module fake_ariane_2636_n_8906 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_730, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_830, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_726, n_603, n_373, n_299, n_836, n_541, n_499, n_789, n_788, n_12, n_771, n_564, n_133, n_610, n_66, n_205, n_752, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_760, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_806, n_367, n_713, n_649, n_598, n_345, n_374, n_318, n_817, n_103, n_244, n_643, n_679, n_226, n_781, n_220, n_261, n_682, n_36, n_663, n_370, n_706, n_189, n_717, n_819, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_776, n_424, n_528, n_584, n_387, n_406, n_826, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_756, n_346, n_214, n_764, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_807, n_138, n_162, n_765, n_264, n_737, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_766, n_372, n_377, n_15, n_396, n_802, n_631, n_23, n_399, n_554, n_520, n_87, n_714, n_279, n_702, n_207, n_790, n_363, n_720, n_354, n_41, n_813, n_140, n_725, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_801, n_202, n_145, n_193, n_733, n_761, n_818, n_500, n_665, n_59, n_336, n_731, n_754, n_779, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_829, n_8, n_668, n_339, n_738, n_758, n_833, n_672, n_487, n_740, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_784, n_269, n_597, n_816, n_75, n_158, n_69, n_259, n_835, n_95, n_808, n_446, n_553, n_143, n_753, n_566, n_814, n_578, n_701, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_822, n_344, n_381, n_795, n_426, n_433, n_481, n_600, n_721, n_840, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_770, n_218, n_821, n_79, n_839, n_3, n_271, n_465, n_486, n_507, n_759, n_247, n_569, n_567, n_825, n_732, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_787, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_703, n_748, n_786, n_510, n_831, n_256, n_326, n_681, n_778, n_227, n_48, n_188, n_323, n_550, n_635, n_707, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_727, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_823, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_777, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_843, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_729, n_661, n_488, n_775, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_846, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_728, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_715, n_579, n_844, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_838, n_237, n_780, n_175, n_711, n_453, n_734, n_74, n_491, n_810, n_19, n_40, n_181, n_723, n_616, n_617, n_658, n_630, n_705, n_570, n_53, n_260, n_362, n_543, n_310, n_709, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_809, n_461, n_209, n_262, n_490, n_743, n_17, n_225, n_235, n_660, n_464, n_735, n_575, n_546, n_297, n_662, n_641, n_503, n_700, n_290, n_527, n_46, n_741, n_747, n_772, n_84, n_847, n_371, n_845, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_708, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_755, n_710, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_842, n_148, n_652, n_451, n_613, n_745, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_716, n_102, n_742, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_798, n_769, n_820, n_43, n_577, n_407, n_774, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_832, n_55, n_535, n_231, n_366, n_744, n_762, n_656, n_555, n_234, n_492, n_574, n_848, n_804, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_794, n_763, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_768, n_514, n_418, n_537, n_223, n_403, n_25, n_750, n_834, n_83, n_389, n_800, n_657, n_513, n_837, n_288, n_179, n_812, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_724, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_722, n_203, n_378, n_436, n_150, n_98, n_757, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_785, n_827, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_746, n_208, n_456, n_156, n_292, n_793, n_174, n_275, n_100, n_704, n_132, n_147, n_204, n_751, n_615, n_521, n_51, n_496, n_739, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_792, n_824, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_719, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_773, n_165, n_144, n_317, n_101, n_243, n_803, n_134, n_329, n_718, n_185, n_340, n_749, n_289, n_9, n_112, n_45, n_542, n_548, n_815, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_782, n_425, n_431, n_811, n_508, n_624, n_118, n_121, n_791, n_618, n_411, n_484, n_712, n_353, n_22, n_736, n_767, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_797, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_828, n_595, n_322, n_251, n_506, n_602, n_799, n_558, n_592, n_116, n_397, n_841, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_796, n_805, n_127, n_531, n_783, n_675, n_8906);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_730;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_830;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_726;
input n_603;
input n_373;
input n_299;
input n_836;
input n_541;
input n_499;
input n_789;
input n_788;
input n_12;
input n_771;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_752;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_760;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_806;
input n_367;
input n_713;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_817;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_781;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_706;
input n_189;
input n_717;
input n_819;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_776;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_826;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_756;
input n_346;
input n_214;
input n_764;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_807;
input n_138;
input n_162;
input n_765;
input n_264;
input n_737;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_766;
input n_372;
input n_377;
input n_15;
input n_396;
input n_802;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_714;
input n_279;
input n_702;
input n_207;
input n_790;
input n_363;
input n_720;
input n_354;
input n_41;
input n_813;
input n_140;
input n_725;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_801;
input n_202;
input n_145;
input n_193;
input n_733;
input n_761;
input n_818;
input n_500;
input n_665;
input n_59;
input n_336;
input n_731;
input n_754;
input n_779;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_829;
input n_8;
input n_668;
input n_339;
input n_738;
input n_758;
input n_833;
input n_672;
input n_487;
input n_740;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_597;
input n_816;
input n_75;
input n_158;
input n_69;
input n_259;
input n_835;
input n_95;
input n_808;
input n_446;
input n_553;
input n_143;
input n_753;
input n_566;
input n_814;
input n_578;
input n_701;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_822;
input n_344;
input n_381;
input n_795;
input n_426;
input n_433;
input n_481;
input n_600;
input n_721;
input n_840;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_770;
input n_218;
input n_821;
input n_79;
input n_839;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_759;
input n_247;
input n_569;
input n_567;
input n_825;
input n_732;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_787;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_703;
input n_748;
input n_786;
input n_510;
input n_831;
input n_256;
input n_326;
input n_681;
input n_778;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_707;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_727;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_823;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_777;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_843;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_729;
input n_661;
input n_488;
input n_775;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_846;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_728;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_715;
input n_579;
input n_844;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_838;
input n_237;
input n_780;
input n_175;
input n_711;
input n_453;
input n_734;
input n_74;
input n_491;
input n_810;
input n_19;
input n_40;
input n_181;
input n_723;
input n_616;
input n_617;
input n_658;
input n_630;
input n_705;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_709;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_809;
input n_461;
input n_209;
input n_262;
input n_490;
input n_743;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_735;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_700;
input n_290;
input n_527;
input n_46;
input n_741;
input n_747;
input n_772;
input n_84;
input n_847;
input n_371;
input n_845;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_708;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_755;
input n_710;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_842;
input n_148;
input n_652;
input n_451;
input n_613;
input n_745;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_716;
input n_102;
input n_742;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_798;
input n_769;
input n_820;
input n_43;
input n_577;
input n_407;
input n_774;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_832;
input n_55;
input n_535;
input n_231;
input n_366;
input n_744;
input n_762;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_848;
input n_804;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_794;
input n_763;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_768;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_750;
input n_834;
input n_83;
input n_389;
input n_800;
input n_657;
input n_513;
input n_837;
input n_288;
input n_179;
input n_812;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_724;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_722;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_757;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_785;
input n_827;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_746;
input n_208;
input n_456;
input n_156;
input n_292;
input n_793;
input n_174;
input n_275;
input n_100;
input n_704;
input n_132;
input n_147;
input n_204;
input n_751;
input n_615;
input n_521;
input n_51;
input n_496;
input n_739;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_792;
input n_824;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_719;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_773;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_803;
input n_134;
input n_329;
input n_718;
input n_185;
input n_340;
input n_749;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_815;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_782;
input n_425;
input n_431;
input n_811;
input n_508;
input n_624;
input n_118;
input n_121;
input n_791;
input n_618;
input n_411;
input n_484;
input n_712;
input n_353;
input n_22;
input n_736;
input n_767;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_797;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_828;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_799;
input n_558;
input n_592;
input n_116;
input n_397;
input n_841;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_796;
input n_805;
input n_127;
input n_531;
input n_783;
input n_675;

output n_8906;

wire n_2752;
wire n_4474;
wire n_3527;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_8165;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_8139;
wire n_4962;
wire n_1430;
wire n_7832;
wire n_8438;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_8321;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_7922;
wire n_7805;
wire n_2790;
wire n_7542;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_8699;
wire n_1131;
wire n_8037;
wire n_5479;
wire n_2646;
wire n_8257;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_8546;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_7001;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_4853;
wire n_8744;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_8449;
wire n_4260;
wire n_903;
wire n_7626;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_7965;
wire n_7368;
wire n_1690;
wire n_8399;
wire n_2807;
wire n_6664;
wire n_8598;
wire n_7562;
wire n_7534;
wire n_1018;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_8460;
wire n_4132;
wire n_1364;
wire n_7373;
wire n_2390;
wire n_8068;
wire n_6891;
wire n_4500;
wire n_2322;
wire n_8734;
wire n_1107;
wire n_8720;
wire n_2663;
wire n_8097;
wire n_5481;
wire n_6539;
wire n_8114;
wire n_4824;
wire n_8422;
wire n_7467;
wire n_8126;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_4741;
wire n_1284;
wire n_1428;
wire n_1241;
wire n_7526;
wire n_8664;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_8326;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_8504;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_7937;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_863;
wire n_6992;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_8035;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_8660;
wire n_3325;
wire n_6681;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_6452;
wire n_1840;
wire n_5247;
wire n_8469;
wire n_8715;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_7507;
wire n_1267;
wire n_8176;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_1213;
wire n_2382;
wire n_7379;
wire n_7441;
wire n_5292;
wire n_1918;
wire n_8327;
wire n_7438;
wire n_8855;
wire n_4443;
wire n_4119;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_7874;
wire n_8539;
wire n_8630;
wire n_8533;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_8435;
wire n_7695;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_8098;
wire n_3754;
wire n_8204;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_7944;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_7850;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_8542;
wire n_8572;
wire n_5046;
wire n_7607;
wire n_7642;
wire n_8373;
wire n_8424;
wire n_8442;
wire n_1386;
wire n_6236;
wire n_7104;
wire n_8147;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_1842;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_8519;
wire n_1692;
wire n_2611;
wire n_8075;
wire n_5468;
wire n_4745;
wire n_3029;
wire n_7638;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_8642;
wire n_8648;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_7259;
wire n_7838;
wire n_8556;
wire n_5984;
wire n_5204;
wire n_6724;
wire n_6705;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_7840;
wire n_8585;
wire n_2745;
wire n_8455;
wire n_2087;
wire n_8444;
wire n_2161;
wire n_6624;
wire n_1357;
wire n_7888;
wire n_8560;
wire n_6710;
wire n_1787;
wire n_6883;
wire n_8108;
wire n_1389;
wire n_8158;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_6659;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_8814;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_7583;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_8130;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_7690;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_7893;
wire n_2954;
wire n_4438;
wire n_6538;
wire n_7966;
wire n_974;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7599;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_7717;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_1447;
wire n_8675;
wire n_1220;
wire n_7900;
wire n_2019;
wire n_5708;
wire n_8123;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_8220;
wire n_2625;
wire n_8355;
wire n_5373;
wire n_7403;
wire n_1578;
wire n_6665;
wire n_8883;
wire n_3147;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_1247;
wire n_6860;
wire n_1568;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_8816;
wire n_4314;
wire n_8418;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_7789;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_8739;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_8243;
wire n_3704;
wire n_8798;
wire n_7963;
wire n_6382;
wire n_8423;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_7938;
wire n_5088;
wire n_6615;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_1743;
wire n_8548;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_8156;
wire n_5138;
wire n_8845;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_8510;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_1665;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_8402;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_8685;
wire n_1828;
wire n_1304;
wire n_7202;
wire n_5960;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_8595;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_7868;
wire n_3370;
wire n_874;
wire n_7654;
wire n_3949;
wire n_2286;
wire n_8779;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_8520;
wire n_4583;
wire n_8555;
wire n_6366;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_7176;
wire n_8565;
wire n_8334;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_7547;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_8030;
wire n_8513;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_8245;
wire n_7942;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_8753;
wire n_1188;
wire n_1498;
wire n_7527;
wire n_4856;
wire n_2618;
wire n_7948;
wire n_7096;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_8485;
wire n_5596;
wire n_6482;
wire n_8106;
wire n_2849;
wire n_1489;
wire n_8325;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_1005;
wire n_8677;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_8626;
wire n_2827;
wire n_7869;
wire n_3214;
wire n_8166;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_6631;
wire n_5889;
wire n_8602;
wire n_7151;
wire n_3944;
wire n_7762;
wire n_5632;
wire n_4729;
wire n_8002;
wire n_6728;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_4800;
wire n_1373;
wire n_7075;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_7611;
wire n_7796;
wire n_6508;
wire n_7989;
wire n_8047;
wire n_2821;
wire n_3696;
wire n_7936;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_8751;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_8800;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_7655;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_951;
wire n_8039;
wire n_8193;
wire n_7546;
wire n_8432;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_8684;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_5463;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_8628;
wire n_3617;
wire n_6012;
wire n_2958;
wire n_7481;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_5435;
wire n_6484;
wire n_5053;
wire n_3340;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_8617;
wire n_7605;
wire n_8591;
wire n_8090;
wire n_1243;
wire n_5511;
wire n_8661;
wire n_3486;
wire n_6639;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_1878;
wire n_7375;
wire n_7076;
wire n_7689;
wire n_6344;
wire n_8189;
wire n_8811;
wire n_7736;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_6600;
wire n_7010;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_8192;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_8573;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_7918;
wire n_1406;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_8339;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_8775;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_8804;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_7295;
wire n_4076;
wire n_7824;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_7600;
wire n_2386;
wire n_5826;
wire n_8697;
wire n_4822;
wire n_6946;
wire n_7947;
wire n_8645;
wire n_5931;
wire n_8820;
wire n_8146;
wire n_1829;
wire n_4635;
wire n_7847;
wire n_8154;
wire n_1450;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_7039;
wire n_8027;
wire n_7807;
wire n_1493;
wire n_2911;
wire n_8063;
wire n_3313;
wire n_8406;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_8480;
wire n_4419;
wire n_8849;
wire n_5405;
wire n_7660;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_5772;
wire n_3345;
wire n_6442;
wire n_8241;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_4906;
wire n_3548;
wire n_6846;
wire n_4630;
wire n_8261;
wire n_6840;
wire n_6645;
wire n_8535;
wire n_8348;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_7831;
wire n_8138;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_8702;
wire n_1995;
wire n_7455;
wire n_8273;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4966;
wire n_2250;
wire n_8235;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_8294;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_8349;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_8429;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_7887;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_8486;
wire n_2070;
wire n_6706;
wire n_7431;
wire n_8140;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_8117;
wire n_3886;
wire n_2619;
wire n_7521;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_8129;
wire n_1291;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_7569;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_7972;
wire n_8672;
wire n_7505;
wire n_3921;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_7524;
wire n_4196;
wire n_1197;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_8847;
wire n_8005;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_6500;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_1398;
wire n_1921;
wire n_8221;
wire n_7573;
wire n_6630;
wire n_5759;
wire n_5629;
wire n_2411;
wire n_4631;
wire n_8191;
wire n_6798;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_7498;
wire n_7895;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_8225;
wire n_3822;
wire n_889;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_7932;
wire n_7890;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6403;
wire n_3497;
wire n_6395;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_8559;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_8689;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_8330;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_8304;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_8163;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_7240;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_1056;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_8777;
wire n_2669;
wire n_8698;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6541;
wire n_6248;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_7927;
wire n_1814;
wire n_7219;
wire n_2441;
wire n_8081;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_7382;
wire n_8384;
wire n_4004;
wire n_5238;
wire n_8650;
wire n_3630;
wire n_1612;
wire n_1910;
wire n_5906;
wire n_7767;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_2931;
wire n_3433;
wire n_8284;
wire n_8374;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_3786;
wire n_875;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_7691;
wire n_3553;
wire n_5323;
wire n_7745;
wire n_6744;
wire n_3645;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_7735;
wire n_8531;
wire n_6116;
wire n_8074;
wire n_3550;
wire n_8780;
wire n_7956;
wire n_5510;
wire n_7651;
wire n_7495;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_8580;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_6757;
wire n_7536;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_8358;
wire n_972;
wire n_7734;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_7671;
wire n_4832;
wire n_8033;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_7926;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_8643;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_7528;
wire n_6209;
wire n_4672;
wire n_8094;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_1127;
wire n_7413;
wire n_7993;
wire n_7821;
wire n_7620;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_8477;
wire n_1775;
wire n_908;
wire n_1036;
wire n_7109;
wire n_8028;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_8530;
wire n_3621;
wire n_5529;
wire n_7561;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_8500;
wire n_6716;
wire n_8713;
wire n_3565;
wire n_7885;
wire n_8297;
wire n_6905;
wire n_8456;
wire n_7722;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_8025;
wire n_5354;
wire n_2453;
wire n_7898;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_4230;
wire n_3040;
wire n_6899;
wire n_7980;
wire n_7817;
wire n_6413;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_8293;
wire n_3211;
wire n_7299;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_8029;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_8880;
wire n_1261;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_857;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_8471;
wire n_1462;
wire n_5701;
wire n_7002;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_8726;
wire n_1813;
wire n_2997;
wire n_7018;
wire n_1573;
wire n_6746;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_8316;
wire n_6174;
wire n_6545;
wire n_7773;
wire n_6763;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_4339;
wire n_7297;
wire n_7730;
wire n_8134;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4169;
wire n_4024;
wire n_3316;
wire n_8610;
wire n_4023;
wire n_4253;
wire n_7637;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_7544;
wire n_2139;
wire n_7613;
wire n_7995;
wire n_8113;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_8724;
wire n_7140;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_8253;
wire n_3303;
wire n_7910;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_7741;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_6668;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_8232;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_8803;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_7679;
wire n_3018;
wire n_8818;
wire n_7698;
wire n_1875;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_1150;
wire n_7800;
wire n_4266;
wire n_6336;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_7835;
wire n_1136;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_8823;
wire n_5399;
wire n_8536;
wire n_8795;
wire n_2846;
wire n_3371;
wire n_8674;
wire n_4918;
wire n_5856;
wire n_8016;
wire n_3872;
wire n_5760;
wire n_7747;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_7552;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_8132;
wire n_7650;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_7535;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_7635;
wire n_4408;
wire n_2115;
wire n_8567;
wire n_8259;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_8578;
wire n_4548;
wire n_7819;
wire n_8495;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_896;
wire n_4574;
wire n_8160;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_8336;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_5548;
wire n_7788;
wire n_6974;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_8600;
wire n_8229;
wire n_4686;
wire n_2384;
wire n_7794;
wire n_1705;
wire n_3895;
wire n_1091;
wire n_3707;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_8761;
wire n_1846;
wire n_7630;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6951;
wire n_6963;
wire n_1581;
wire n_946;
wire n_3058;
wire n_5355;
wire n_2047;
wire n_1655;
wire n_3709;
wire n_3398;
wire n_1146;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_8473;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_8351;
wire n_5915;
wire n_7276;
wire n_6379;
wire n_1368;
wire n_963;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_925;
wire n_7753;
wire n_6834;
wire n_2880;
wire n_4716;
wire n_1001;
wire n_1313;
wire n_3722;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_7541;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_7913;
wire n_8020;
wire n_7946;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_8875;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_7920;
wire n_1931;
wire n_5559;
wire n_8649;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_1820;
wire n_7841;
wire n_7160;
wire n_7324;
wire n_8205;
wire n_6046;
wire n_7054;
wire n_4493;
wire n_1233;
wire n_6055;
wire n_7161;
wire n_1808;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_1635;
wire n_8440;
wire n_1704;
wire n_4896;
wire n_8041;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_886;
wire n_7837;
wire n_6788;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_5528;
wire n_7806;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_8076;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_8757;
wire n_1355;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_8897;
wire n_7676;
wire n_8177;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_1169;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_7644;
wire n_4602;
wire n_1713;
wire n_7816;
wire n_8829;
wire n_2818;
wire n_1436;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_8638;
wire n_1515;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_952;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_7724;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_8101;
wire n_2374;
wire n_5439;
wire n_8687;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_8721;
wire n_1366;
wire n_8749;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_7879;
wire n_8730;
wire n_6607;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_4660;
wire n_8503;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_8315;
wire n_1961;
wire n_1535;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_871;
wire n_6807;
wire n_2844;
wire n_8197;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_4814;
wire n_8019;
wire n_8801;
wire n_6178;
wire n_8707;
wire n_6677;
wire n_2221;
wire n_7875;
wire n_5502;
wire n_8248;
wire n_1283;
wire n_7550;
wire n_8554;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_8501;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_7804;
wire n_5098;
wire n_1084;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_1276;
wire n_8263;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_8040;
wire n_5466;
wire n_1528;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_7826;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_8102;
wire n_3999;
wire n_8196;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_8822;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_7971;
wire n_8885;
wire n_5592;
wire n_5620;
wire n_5491;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_8474;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_4597;
wire n_1636;
wire n_8152;
wire n_8269;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_4576;
wire n_7577;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_8144;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_7812;
wire n_5330;
wire n_6935;
wire n_1560;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_8058;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_2722;
wire n_3728;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_6781;
wire n_7667;
wire n_4593;
wire n_8024;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_1391;
wire n_8107;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_6741;
wire n_1245;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_6593;
wire n_7827;
wire n_3758;
wire n_7631;
wire n_8748;
wire n_8452;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_8742;
wire n_3777;
wire n_8393;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_8122;
wire n_2426;
wire n_6947;
wire n_8403;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_8740;
wire n_5574;
wire n_8310;
wire n_3391;
wire n_5877;
wire n_912;
wire n_6375;
wire n_7781;
wire n_4786;
wire n_6042;
wire n_8238;
wire n_5203;
wire n_7908;
wire n_8296;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_7855;
wire n_8850;
wire n_2855;
wire n_2848;
wire n_7886;
wire n_7675;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_7774;
wire n_8634;
wire n_8831;
wire n_6970;
wire n_1026;
wire n_6948;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_8676;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_8758;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_8544;
wire n_3240;
wire n_7999;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_8652;
wire n_2836;
wire n_7873;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_8646;
wire n_2172;
wire n_2601;
wire n_2365;
wire n_1880;
wire n_5684;
wire n_1399;
wire n_7228;
wire n_5981;
wire n_7784;
wire n_1855;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_7713;
wire n_6623;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_2224;
wire n_1226;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_8031;
wire n_3257;
wire n_5737;
wire n_8015;
wire n_8412;
wire n_3730;
wire n_8439;
wire n_8575;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_976;
wire n_4003;
wire n_1832;
wire n_8499;
wire n_6390;
wire n_7640;
wire n_2302;
wire n_6799;
wire n_8772;
wire n_3014;
wire n_7912;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_8557;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_7641;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_8815;
wire n_7949;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_8679;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_1020;
wire n_7764;
wire n_8446;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_8789;
wire n_8128;
wire n_7520;
wire n_5314;
wire n_7616;
wire n_8359;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_1279;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_8678;
wire n_1689;
wire n_8605;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_8443;
wire n_8525;
wire n_1401;
wire n_3138;
wire n_8312;
wire n_2860;
wire n_8901;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_6387;
wire n_4201;
wire n_6470;
wire n_7206;
wire n_8869;
wire n_5287;
wire n_8272;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_1217;
wire n_6341;
wire n_2662;
wire n_4386;
wire n_6374;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_8870;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_8178;
wire n_5524;
wire n_7854;
wire n_926;
wire n_2296;
wire n_5735;
wire n_7959;
wire n_8234;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_7897;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_8488;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_1570;
wire n_7533;
wire n_3377;
wire n_6722;
wire n_1518;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_7766;
wire n_855;
wire n_8862;
wire n_2059;
wire n_8184;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_1287;
wire n_1611;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_7776;
wire n_4818;
wire n_8001;
wire n_8695;
wire n_7436;
wire n_8767;
wire n_8571;
wire n_7020;
wire n_5935;
wire n_8064;
wire n_6696;
wire n_4916;
wire n_8472;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_7978;
wire n_5488;
wire n_1105;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_8787;
wire n_8131;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_7694;
wire n_8771;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_983;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_8150;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_1092;
wire n_4374;
wire n_3205;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_8230;
wire n_6222;
wire n_2218;
wire n_8352;
wire n_1122;
wire n_7760;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_8821;
wire n_8465;
wire n_6587;
wire n_6688;
wire n_8360;
wire n_6505;
wire n_5362;
wire n_8209;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_7629;
wire n_6987;
wire n_877;
wire n_3995;
wire n_7567;
wire n_8743;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_1055;
wire n_8396;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_8514;
wire n_8550;
wire n_1089;
wire n_7449;
wire n_8151;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3568;
wire n_3216;
wire n_2708;
wire n_6187;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_7479;
wire n_7882;
wire n_1649;
wire n_2470;
wire n_7517;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_8070;
wire n_4525;
wire n_8866;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_7878;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_8797;
wire n_6547;
wire n_7177;
wire n_7902;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_8054;
wire n_982;
wire n_3791;
wire n_915;
wire n_6478;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_8841;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_7590;
wire n_6906;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_1319;
wire n_3669;
wire n_3367;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_7818;
wire n_7645;
wire n_5385;
wire n_7482;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_8618;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_8538;
wire n_3582;
wire n_8590;
wire n_7907;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_8791;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_7862;
wire n_3735;
wire n_8703;
wire n_7565;
wire n_7410;
wire n_6422;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_7721;
wire n_4524;
wire n_8061;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_8754;
wire n_8864;
wire n_5941;
wire n_4891;
wire n_8837;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_8784;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_8768;
wire n_6999;
wire n_8086;
wire n_8072;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_7539;
wire n_6440;
wire n_4977;
wire n_8774;
wire n_2492;
wire n_6976;
wire n_7608;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_2912;
wire n_5936;
wire n_8307;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1757;
wire n_8470;
wire n_1950;
wire n_2264;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_7830;
wire n_8050;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_1281;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_5504;
wire n_878;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_8010;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_6464;
wire n_8802;
wire n_5129;
wire n_1350;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_8603;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_1616;
wire n_7935;
wire n_2416;
wire n_8143;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_7933;
wire n_1557;
wire n_6640;
wire n_7155;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_6850;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_7743;
wire n_4990;
wire n_2986;
wire n_8584;
wire n_949;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_8153;
wire n_6972;
wire n_3591;
wire n_8574;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_7043;
wire n_7986;
wire n_3317;
wire n_8049;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_7996;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_8509;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_4790;
wire n_7035;
wire n_4173;
wire n_8354;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_8277;
wire n_7442;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_8583;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_8681;
wire n_6258;
wire n_1288;
wire n_8644;
wire n_7939;
wire n_7715;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_8609;
wire n_1143;
wire n_3973;
wire n_8052;
wire n_4799;
wire n_8733;
wire n_8082;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_7699;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_7580;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_5911;
wire n_7340;
wire n_8080;
wire n_3600;
wire n_7303;
wire n_1023;
wire n_8819;
wire n_914;
wire n_7870;
wire n_6139;
wire n_7568;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_8487;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_8382;
wire n_1417;
wire n_3096;
wire n_8517;
wire n_7207;
wire n_8827;
wire n_4166;
wire n_5356;
wire n_2777;
wire n_7167;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_8203;
wire n_2935;
wire n_4246;
wire n_7618;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_8340;
wire n_4754;
wire n_1534;
wire n_8268;
wire n_8171;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_8008;
wire n_7633;
wire n_3117;
wire n_4684;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_8553;
wire n_2592;
wire n_8824;
wire n_3490;
wire n_7280;
wire n_8369;
wire n_962;
wire n_5043;
wire n_7339;
wire n_7597;
wire n_8884;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_7768;
wire n_918;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_6455;
wire n_2842;
wire n_7615;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_8271;
wire n_3720;
wire n_6183;
wire n_8392;
wire n_8309;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_4256;
wire n_2560;
wire n_1164;
wire n_8874;
wire n_8228;
wire n_1193;
wire n_5035;
wire n_1345;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_8483;
wire n_6003;
wire n_5443;
wire n_8133;
wire n_7612;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_8172;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_8344;
wire n_7594;
wire n_7711;
wire n_7321;
wire n_4457;
wire n_2150;
wire n_8738;
wire n_6785;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_7574;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_8226;
wire n_6695;
wire n_7529;
wire n_5608;
wire n_3354;
wire n_6501;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_7522;
wire n_7188;
wire n_8088;
wire n_5702;
wire n_8662;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_8783;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_8663;
wire n_5277;
wire n_1262;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_4048;
wire n_3807;
wire n_6213;
wire n_1579;
wire n_8364;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_8490;
wire n_923;
wire n_1124;
wire n_7872;
wire n_1326;
wire n_3969;
wire n_6873;
wire n_7958;
wire n_2282;
wire n_4605;
wire n_8118;
wire n_981;
wire n_4649;
wire n_3873;
wire n_5747;
wire n_8671;
wire n_7101;
wire n_8785;
wire n_1204;
wire n_7843;
wire n_2428;
wire n_994;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_7578;
wire n_3410;
wire n_5415;
wire n_856;
wire n_7261;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_6993;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_8100;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_8522;
wire n_1361;
wire n_8381;
wire n_8835;
wire n_6767;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_7263;
wire n_3782;
wire n_1317;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_7688;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7925;
wire n_7310;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_7585;
wire n_8356;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_7772;
wire n_8736;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_1550;
wire n_1358;
wire n_8616;
wire n_1200;
wire n_6105;
wire n_5512;
wire n_7738;
wire n_2808;
wire n_2344;
wire n_8838;
wire n_3520;
wire n_2392;
wire n_7609;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_8607;
wire n_8213;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_8436;
wire n_7282;
wire n_8551;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_7921;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_6331;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_7863;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_7968;
wire n_6023;
wire n_7820;
wire n_8437;
wire n_7833;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_7750;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_7588;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_7697;
wire n_5887;
wire n_7808;
wire n_3068;
wire n_1629;
wire n_7603;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_8704;
wire n_3002;
wire n_7192;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_8613;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_8012;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_8881;
wire n_5531;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_2351;
wire n_1619;
wire n_7988;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_8763;
wire n_6450;
wire n_1152;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_1236;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_8387;
wire n_8105;
wire n_2704;
wire n_1334;
wire n_6745;
wire n_7943;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_8900;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_8353;
wire n_2048;
wire n_7723;
wire n_3028;
wire n_4691;
wire n_7904;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_8323;
wire n_6164;
wire n_8711;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_8731;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_7759;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_8597;
wire n_2515;
wire n_6330;
wire n_1600;
wire n_1144;
wire n_7178;
wire n_1941;
wire n_7045;
wire n_3637;
wire n_8534;
wire n_1017;
wire n_8655;
wire n_4893;
wire n_2240;
wire n_7777;
wire n_8302;
wire n_4258;
wire n_5756;
wire n_8496;
wire n_7693;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_8078;
wire n_2097;
wire n_3461;
wire n_7682;
wire n_7300;
wire n_939;
wire n_2297;
wire n_1410;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_7558;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_8103;
wire n_8719;
wire n_1983;
wire n_7798;
wire n_8879;
wire n_4767;
wire n_4569;
wire n_948;
wire n_6528;
wire n_8896;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_8335;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_8116;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_1571;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_933;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_8462;
wire n_3228;
wire n_8834;
wire n_8286;
wire n_8417;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_7672;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_3088;
wire n_1724;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_8247;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_8639;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_7712;
wire n_6885;
wire n_7681;
wire n_5039;
wire n_1818;
wire n_6580;
wire n_6613;
wire n_8566;
wire n_8727;
wire n_4265;
wire n_8482;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_7491;
wire n_1583;
wire n_8599;
wire n_4612;
wire n_5997;
wire n_8781;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_7954;
wire n_7974;
wire n_1264;
wire n_6530;
wire n_6602;
wire n_7915;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_8839;
wire n_1752;
wire n_2361;
wire n_3030;
wire n_4538;
wire n_5563;
wire n_3505;
wire n_3075;
wire n_8365;
wire n_1102;
wire n_2239;
wire n_6942;
wire n_7860;
wire n_6892;
wire n_1296;
wire n_4730;
wire n_7357;
wire n_8112;
wire n_8489;
wire n_8859;
wire n_8060;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_8244;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_8096;
wire n_7336;
wire n_5932;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_8346;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_8367;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_2797;
wire n_5823;
wire n_8658;
wire n_8898;
wire n_2423;
wire n_2208;
wire n_1421;
wire n_5422;
wire n_5944;
wire n_8905;
wire n_6989;
wire n_8145;
wire n_8237;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_8562;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_7273;
wire n_7901;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_7149;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_8211;
wire n_3268;
wire n_2559;
wire n_8537;
wire n_5616;
wire n_1383;
wire n_8055;
wire n_4259;
wire n_5870;
wire n_7909;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_6758;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_8332;
wire n_5601;
wire n_4965;
wire n_3742;
wire n_7601;
wire n_1837;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_8157;
wire n_2006;
wire n_4953;
wire n_8484;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_7596;
wire n_5294;
wire n_8161;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5670;
wire n_5411;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_7549;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_8692;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_6918;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_8812;
wire n_8682;
wire n_4796;
wire n_8290;
wire n_1088;
wire n_7138;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_7976;
wire n_2750;
wire n_8890;
wire n_2547;
wire n_8747;
wire n_7617;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_8062;
wire n_3281;
wire n_7137;
wire n_5061;
wire n_3535;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7700;
wire n_8275;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_8667;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_5575;
wire n_6654;
wire n_7661;
wire n_4968;
wire n_7801;
wire n_8807;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_7876;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_7323;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_8048;
wire n_5607;
wire n_1514;
wire n_7929;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_8212;
wire n_4950;
wire n_1650;
wire n_7755;
wire n_6504;
wire n_4176;
wire n_7556;
wire n_4124;
wire n_4431;
wire n_3347;
wire n_1404;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_8043;
wire n_8223;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_8159;
wire n_5845;
wire n_8868;
wire n_4608;
wire n_6691;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_8434;
wire n_3634;
wire n_5436;
wire n_7962;
wire n_2341;
wire n_1654;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_8608;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_8656;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_7905;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_8249;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_5718;
wire n_7208;
wire n_7718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_6567;
wire n_5658;
wire n_1112;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_7756;
wire n_5546;
wire n_6294;
wire n_7795;
wire n_7822;
wire n_8717;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_7623;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_7632;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_8842;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_8073;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_8576;
wire n_916;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_1555;
wire n_8799;
wire n_1468;
wire n_4378;
wire n_1253;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_8181;
wire n_5808;
wire n_1182;
wire n_6527;
wire n_4594;
wire n_8447;
wire n_8045;
wire n_7289;
wire n_7538;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_1376;
wire n_7473;
wire n_7242;
wire n_6533;
wire n_7164;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_8022;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_8227;
wire n_7853;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_7483;
wire n_8756;
wire n_5710;
wire n_1491;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_5333;
wire n_1083;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_8604;
wire n_8809;
wire n_3510;
wire n_7046;
wire n_7834;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_8844;
wire n_6148;
wire n_2100;
wire n_8255;
wire n_5538;
wire n_3666;
wire n_990;
wire n_6357;
wire n_867;
wire n_8216;
wire n_8693;
wire n_3479;
wire n_944;
wire n_5499;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_7811;
wire n_8669;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_7880;
wire n_8769;
wire n_909;
wire n_6713;
wire n_8149;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_7851;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_7810;
wire n_6108;
wire n_7664;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_7477;
wire n_1914;
wire n_8208;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_7714;
wire n_7899;
wire n_8710;
wire n_6415;
wire n_8479;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_8512;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_7845;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_7858;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_6392;
wire n_6513;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_6720;
wire n_5883;
wire n_8401;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_7680;
wire n_5630;
wire n_6666;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_6815;
wire n_1387;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_8450;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_7710;
wire n_8788;
wire n_5394;
wire n_8324;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_8104;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_8014;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_8623;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_8651;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_5132;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_7783;
wire n_7662;
wire n_6057;
wire n_6936;
wire n_4728;
wire n_7171;
wire n_7990;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_7003;
wire n_8137;
wire n_2187;
wire n_1413;
wire n_8413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_8300;
wire n_8069;
wire n_7501;
wire n_6432;
wire n_7984;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_1423;
wire n_8173;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_7589;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_1798;
wire n_8091;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_6699;
wire n_3983;
wire n_8254;
wire n_8400;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_6957;
wire n_5074;
wire n_7917;
wire n_3939;
wire n_3788;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_8368;
wire n_6694;
wire n_3260;
wire n_2496;
wire n_8463;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_1602;
wire n_7422;
wire n_3139;
wire n_8889;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_8322;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_7621;
wire n_8274;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_1205;
wire n_6195;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_7572;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_7500;
wire n_1202;
wire n_4084;
wire n_7985;
wire n_1371;
wire n_4240;
wire n_8657;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_8311;
wire n_5748;
wire n_4393;
wire n_6662;
wire n_7494;
wire n_3984;
wire n_1586;
wire n_8728;
wire n_1431;
wire n_4389;
wire n_6433;
wire n_1763;
wire n_8398;
wire n_6200;
wire n_5641;
wire n_8407;
wire n_8071;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3492;
wire n_3044;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_8528;
wire n_5657;
wire n_8475;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_5244;
wire n_1677;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_6956;
wire n_7587;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_7704;
wire n_5420;
wire n_6497;
wire n_8511;
wire n_7865;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_6701;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_8867;
wire n_3417;
wire n_8246;
wire n_8558;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_7881;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_8641;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_1800;
wire n_7198;
wire n_6884;
wire n_7752;
wire n_5081;
wire n_8201;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_7953;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_8046;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_8414;
wire n_3024;
wire n_5567;
wire n_8292;
wire n_5406;
wire n_8647;
wire n_6362;
wire n_4328;
wire n_8543;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_8331;
wire n_999;
wire n_2280;
wire n_8317;
wire n_7126;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_6678;
wire n_7982;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_8187;
wire n_8174;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_8846;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_8032;
wire n_5417;
wire n_4545;
wire n_8200;
wire n_4758;
wire n_1161;
wire n_8036;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_8586;
wire n_8524;
wire n_1191;
wire n_4535;
wire n_7518;
wire n_8828;
wire n_4385;
wire n_7779;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_7575;
wire n_2337;
wire n_7073;
wire n_8092;
wire n_1786;
wire n_6309;
wire n_8370;
wire n_3732;
wire n_1804;
wire n_8135;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1318;
wire n_8764;
wire n_1632;
wire n_1769;
wire n_7349;
wire n_1929;
wire n_8502;
wire n_4319;
wire n_6585;
wire n_7786;
wire n_8454;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_7579;
wire n_7122;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_6490;
wire n_7867;
wire n_4651;
wire n_943;
wire n_4748;
wire n_3167;
wire n_7624;
wire n_1807;
wire n_1123;
wire n_8776;
wire n_2857;
wire n_8564;
wire n_8343;
wire n_7828;
wire n_1784;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_8718;
wire n_985;
wire n_5506;
wire n_7543;
wire n_5475;
wire n_8042;
wire n_7727;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_8379;
wire n_8034;
wire n_7778;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_7019;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_8441;
wire n_2353;
wire n_1429;
wire n_7702;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_6685;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_8569;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_8592;
wire n_8865;
wire n_3976;
wire n_2813;
wire n_897;
wire n_3381;
wire n_2546;
wire n_7952;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_7791;
wire n_6971;
wire n_8362;
wire n_3336;
wire n_8632;
wire n_7739;
wire n_7945;
wire n_8361;
wire n_7656;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_8561;
wire n_6549;
wire n_8611;
wire n_8410;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_5912;
wire n_5745;
wire n_7923;
wire n_6086;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_8878;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_8492;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_8888;
wire n_6820;
wire n_2497;
wire n_879;
wire n_5446;
wire n_7610;
wire n_7107;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_7456;
wire n_8095;
wire n_7369;
wire n_1472;
wire n_1050;
wire n_7548;
wire n_2578;
wire n_1201;
wire n_8735;
wire n_7598;
wire n_2475;
wire n_1185;
wire n_7250;
wire n_8808;
wire n_8902;
wire n_7823;
wire n_8833;
wire n_4715;
wire n_6157;
wire n_8796;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_8794;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_1090;
wire n_8549;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_7525;
wire n_4418;
wire n_7924;
wire n_3341;
wire n_8690;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_8593;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_6923;
wire n_2036;
wire n_7649;
wire n_8009;
wire n_8195;
wire n_8588;
wire n_3358;
wire n_6704;
wire n_7634;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_7406;
wire n_4682;
wire n_1128;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_8805;
wire n_5078;
wire n_4810;
wire n_7659;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_8596;
wire n_1549;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_7844;
wire n_5207;
wire n_7934;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_7009;
wire n_3376;
wire n_7371;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_7463;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5755;
wire n_5700;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_8627;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_1038;
wire n_3723;
wire n_7941;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_8858;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_1022;
wire n_5465;
wire n_8745;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_8169;
wire n_6184;
wire n_8018;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_4138;
wire n_7083;
wire n_1973;
wire n_1444;
wire n_8260;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_7701;
wire n_8688;
wire n_7969;
wire n_8279;
wire n_4384;
wire n_8793;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_7683;
wire n_2154;
wire n_7669;
wire n_1986;
wire n_8298;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_8023;
wire n_7330;
wire n_6007;
wire n_6734;
wire n_6535;
wire n_8053;
wire n_8059;
wire n_1772;
wire n_6879;
wire n_3106;
wire n_1311;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_7692;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_6457;
wire n_4924;
wire n_4044;
wire n_8372;
wire n_6270;
wire n_2305;
wire n_8737;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_1028;
wire n_8723;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_8419;
wire n_2809;
wire n_5652;
wire n_8893;
wire n_975;
wire n_1645;
wire n_5805;
wire n_7304;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_8077;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_7754;
wire n_8826;
wire n_3178;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_7981;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_8712;
wire n_1011;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_8109;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_7877;
wire n_7787;
wire n_7836;
wire n_8515;
wire n_8725;
wire n_8007;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_5902;
wire n_987;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_8301;
wire n_6764;
wire n_7871;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_8892;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_7571;
wire n_8252;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_6955;
wire n_7563;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_8494;
wire n_6569;
wire n_1630;
wire n_7919;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_8278;
wire n_3431;
wire n_8180;
wire n_3355;
wire n_7031;
wire n_1738;
wire n_5716;
wire n_8891;
wire n_3897;
wire n_7103;
wire n_6605;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_8270;
wire n_8231;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_6832;
wire n_5980;
wire n_8683;
wire n_956;
wire n_4092;
wire n_4875;
wire n_7771;
wire n_8903;
wire n_4255;
wire n_2758;
wire n_6544;
wire n_8810;
wire n_6469;
wire n_5036;
wire n_1271;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_8264;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_8288;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_1285;
wire n_6289;
wire n_3838;
wire n_6651;
wire n_8882;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_8388;
wire n_5445;
wire n_2734;
wire n_8067;
wire n_8385;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_8670;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_7706;
wire n_7813;
wire n_8142;
wire n_2420;
wire n_7992;
wire n_7643;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_7628;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_8224;
wire n_5472;
wire n_6035;
wire n_1754;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_8345;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_8614;
wire n_8242;
wire n_6786;
wire n_4564;
wire n_8299;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_8110;
wire n_5072;
wire n_8529;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_8700;
wire n_6766;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_7802;
wire n_7519;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_2933;
wire n_8468;
wire n_7515;
wire n_3387;
wire n_7639;
wire n_6214;
wire n_3952;
wire n_8636;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_7049;
wire n_7884;
wire n_6945;
wire n_8378;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_7749;
wire n_7592;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_8283;
wire n_977;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_7914;
wire n_1866;
wire n_8860;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_6447;
wire n_5859;
wire n_4390;
wire n_1782;
wire n_7892;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4609;
wire n_4361;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_1393;
wire n_7674;
wire n_8686;
wire n_6175;
wire n_6445;
wire n_8563;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_8493;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_6499;
wire n_1982;
wire n_7983;
wire n_5311;
wire n_8765;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_7361;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2982;
wire n_1273;
wire n_8653;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_8601;
wire n_1043;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_8333;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_7309;
wire n_7119;
wire n_1613;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_7696;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_954;
wire n_2051;
wire n_3196;
wire n_8708;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_8659;
wire n_6732;
wire n_8759;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_7646;
wire n_3779;
wire n_6982;
wire n_1063;
wire n_7291;
wire n_8790;
wire n_991;
wire n_2275;
wire n_7668;
wire n_7435;
wire n_4606;
wire n_8832;
wire n_8305;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_8453;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_7017;
wire n_4072;
wire n_7848;
wire n_2792;
wire n_4465;
wire n_8127;
wire n_2596;
wire n_5217;
wire n_8337;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_7861;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_7889;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_7554;
wire n_3202;
wire n_8508;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_7648;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_7653;
wire n_6400;
wire n_1644;
wire n_7846;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_8347;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_5135;
wire n_7551;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_1434;
wire n_8093;
wire n_8899;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_7737;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_8481;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_7606;
wire n_7420;
wire n_8115;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_8182;
wire n_1981;
wire n_2824;
wire n_7973;
wire n_7545;
wire n_5327;
wire n_4417;
wire n_1374;
wire n_2089;
wire n_7896;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_8629;
wire n_8186;
wire n_7319;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_8233;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_8282;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_1463;
wire n_4626;
wire n_7625;
wire n_8750;
wire n_4997;
wire n_8183;
wire n_5065;
wire n_6806;
wire n_924;
wire n_7991;
wire n_8637;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_8792;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_7857;
wire n_7970;
wire n_1706;
wire n_2461;
wire n_8258;
wire n_3719;
wire n_7154;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_5295;
wire n_1503;
wire n_8416;
wire n_8390;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_8696;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_3905;
wire n_1457;
wire n_7163;
wire n_3797;
wire n_1836;
wire n_7027;
wire n_3416;
wire n_8552;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_7964;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_8619;
wire n_7068;
wire n_2908;
wire n_8594;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_8162;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_7327;
wire n_1277;
wire n_1746;
wire n_6610;
wire n_1062;
wire n_5998;
wire n_8318;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_8425;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_7864;
wire n_3451;
wire n_8051;
wire n_4734;
wire n_6675;
wire n_7955;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_1718;
wire n_7814;
wire n_8389;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_8620;
wire n_5555;
wire n_2078;
wire n_8886;
wire n_1145;
wire n_4809;
wire n_7152;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_8202;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_1314;
wire n_8755;
wire n_1512;
wire n_8668;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_7761;
wire n_8141;
wire n_3793;
wire n_5042;
wire n_859;
wire n_3230;
wire n_8199;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_8004;
wire n_8383;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_1751;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_8895;
wire n_8680;
wire n_1548;
wire n_4987;
wire n_6714;
wire n_8394;
wire n_7849;
wire n_7726;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_8198;
wire n_1354;
wire n_8665;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_7859;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_8017;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_7523;
wire n_5234;
wire n_1416;
wire n_6890;
wire n_7559;
wire n_7576;
wire n_6988;
wire n_8303;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_8000;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7769;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_8852;
wire n_5007;
wire n_8709;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_7729;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_8782;
wire n_7081;
wire n_7742;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_4775;
wire n_1442;
wire n_6256;
wire n_2620;
wire n_1833;
wire n_8716;
wire n_1691;
wire n_8250;
wire n_7264;
wire n_7842;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_6649;
wire n_8714;
wire n_1656;
wire n_8357;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_955;
wire n_8466;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_6431;
wire n_8589;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_8266;
wire n_3839;
wire n_8587;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_8876;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_8498;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_8457;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_8267;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_8124;
wire n_3604;
wire n_8545;
wire n_5430;
wire n_6041;
wire n_8526;
wire n_8319;
wire n_7997;
wire n_5659;
wire n_6859;
wire n_7716;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_7950;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_8581;
wire n_8214;
wire n_7793;
wire n_8516;
wire n_2083;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_7746;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_7570;
wire n_2898;
wire n_1825;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_7829;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_1731;
wire n_7894;
wire n_1147;
wire n_7957;
wire n_8262;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_8289;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_7121;
wire n_7531;
wire n_6410;
wire n_6473;
wire n_8087;
wire n_4056;
wire n_4806;
wire n_7961;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_7687;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_8863;
wire n_4517;
wire n_2896;
wire n_8701;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_8705;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_6975;
wire n_7763;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_7703;
wire n_7928;
wire n_4234;
wire n_1483;
wire n_1363;
wire n_8722;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_3179;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_7677;
wire n_5262;
wire n_7665;
wire n_3262;
wire n_5319;
wire n_927;
wire n_7469;
wire n_3699;
wire n_6118;
wire n_2120;
wire n_7125;
wire n_7856;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_1419;
wire n_8622;
wire n_3816;
wire n_8099;
wire n_8729;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_8085;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_7203;
wire n_7797;
wire n_1826;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_5335;
wire n_1259;
wire n_6365;
wire n_8459;
wire n_7111;
wire n_2801;
wire n_4334;
wire n_1177;
wire n_8478;
wire n_5284;
wire n_8786;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_8887;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_8851;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_8540;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_8276;
wire n_7057;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_8706;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_8532;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_6772;
wire n_7088;
wire n_7799;
wire n_5698;
wire n_5731;
wire n_8871;
wire n_4007;
wire n_1456;
wire n_8433;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_7979;
wire n_6617;
wire n_7725;
wire n_5120;
wire n_3572;
wire n_8371;
wire n_2975;
wire n_2399;
wire n_8547;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_8467;
wire n_2027;
wire n_2932;
wire n_8409;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_6777;
wire n_8640;
wire n_6742;
wire n_1467;
wire n_7447;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_8431;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_8415;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_6479;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_8329;
wire n_2599;
wire n_3988;
wire n_7792;
wire n_5022;
wire n_8089;
wire n_6370;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_1098;
wire n_3009;
wire n_8633;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_8541;
wire n_8762;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_1132;
wire n_8125;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_7530;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_7471;
wire n_6465;
wire n_8188;
wire n_5673;
wire n_861;
wire n_8615;
wire n_5814;
wire n_1666;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_8011;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_3326;
wire n_8624;
wire n_8222;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_8206;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_8065;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_7709;
wire n_4269;
wire n_1927;
wire n_7540;
wire n_7581;
wire n_1222;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_7782;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_4913;
wire n_1460;
wire n_8155;
wire n_2449;
wire n_4428;
wire n_6483;
wire n_1572;
wire n_7770;
wire n_8397;
wire n_8568;
wire n_4463;
wire n_5357;
wire n_8175;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_8026;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_8836;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_8168;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7751;
wire n_7951;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_8873;
wire n_7591;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_7911;
wire n_3795;
wire n_7595;
wire n_4931;
wire n_2306;
wire n_7790;
wire n_2071;
wire n_7426;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_6855;
wire n_8170;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_8120;
wire n_8825;
wire n_852;
wire n_2916;
wire n_7252;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_7532;
wire n_4192;
wire n_8003;
wire n_1748;
wire n_1301;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_8395;
wire n_7065;
wire n_1466;
wire n_8083;
wire n_6177;
wire n_8057;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_7367;
wire n_8164;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1037;
wire n_8877;
wire n_1329;
wire n_6825;
wire n_7614;
wire n_1993;
wire n_1545;
wire n_6460;
wire n_4035;
wire n_6952;
wire n_1480;
wire n_3670;
wire n_8366;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_8476;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_7685;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_7619;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_5577;
wire n_876;
wire n_5872;
wire n_7883;
wire n_6692;
wire n_5017;
wire n_8854;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_7560;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_8256;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_1658;
wire n_1072;
wire n_8621;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_8577;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_7731;
wire n_6626;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_7034;
wire n_8654;
wire n_3694;
wire n_6854;
wire n_7940;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_7537;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_1824;
wire n_7740;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_2945;
wire n_3543;
wire n_1971;
wire n_1324;
wire n_8421;
wire n_7179;
wire n_1776;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_3609;
wire n_2936;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_7658;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_7987;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_5401;
wire n_4595;
wire n_960;
wire n_7272;
wire n_8215;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_7906;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_7765;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_4611;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_7815;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_8121;
wire n_5252;
wire n_5777;
wire n_7785;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_8280;
wire n_7728;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_7181;
wire n_2796;
wire n_858;
wire n_5393;
wire n_8328;
wire n_4817;
wire n_8861;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_8427;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_7825;
wire n_1565;
wire n_4437;
wire n_6419;
wire n_7916;
wire n_3055;
wire n_8194;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_7903;
wire n_7089;
wire n_1045;
wire n_8217;
wire n_1881;
wire n_2635;
wire n_7604;
wire n_7647;
wire n_2999;
wire n_988;
wire n_4769;
wire n_4139;
wire n_6130;
wire n_5868;
wire n_6417;
wire n_8285;
wire n_7145;
wire n_8521;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_7803;
wire n_2713;
wire n_1422;
wire n_8448;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_8732;
wire n_7622;
wire n_7839;
wire n_6792;
wire n_7720;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_8136;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_1049;
wire n_8420;
wire n_4430;
wire n_8386;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_1356;
wire n_6831;
wire n_4544;
wire n_3175;
wire n_1773;
wire n_2666;
wire n_5578;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_7809;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_8746;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_8857;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_7564;
wire n_5863;
wire n_8185;
wire n_8313;
wire n_6633;
wire n_3790;
wire n_7775;
wire n_907;
wire n_7118;
wire n_7960;
wire n_6152;
wire n_5734;
wire n_8281;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_7636;
wire n_4341;
wire n_1694;
wire n_6925;
wire n_7186;
wire n_8766;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_8066;
wire n_7666;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_7967;
wire n_5977;
wire n_8314;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_8239;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_8497;
wire n_1157;
wire n_7262;
wire n_5959;
wire n_8056;
wire n_8210;
wire n_3563;
wire n_5945;
wire n_4423;
wire n_2642;
wire n_3310;
wire n_1739;
wire n_3689;
wire n_7584;
wire n_7748;
wire n_1789;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_7686;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_4350;
wire n_1756;
wire n_1606;
wire n_5600;
wire n_6737;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_8404;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_6459;
wire n_1427;
wire n_7670;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_8505;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_8606;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_6448;
wire n_5186;
wire n_7930;
wire n_7487;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_7077;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_8518;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_5604;
wire n_3470;
wire n_7663;
wire n_8350;
wire n_8741;
wire n_5221;
wire n_7024;
wire n_1407;
wire n_8148;
wire n_8408;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_8236;
wire n_7214;
wire n_8806;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_8295;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_7977;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_8167;
wire n_8377;
wire n_3989;
wire n_7652;
wire n_4644;
wire n_4752;
wire n_8673;
wire n_4746;
wire n_7566;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_8760;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_8207;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_8904;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_7678;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_7975;
wire n_8451;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_7553;
wire n_8527;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_7086;
wire n_5689;
wire n_7732;
wire n_7891;
wire n_4578;
wire n_8840;
wire n_5644;
wire n_3644;
wire n_8038;
wire n_8190;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_8179;
wire n_7038;
wire n_7994;
wire n_4470;
wire n_4187;
wire n_8287;
wire n_1904;
wire n_8111;
wire n_8341;
wire n_8830;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_8308;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_8021;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_7593;
wire n_8265;
wire n_898;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_7757;
wire n_1093;
wire n_8251;
wire n_7866;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_8773;
wire n_5947;
wire n_6242;
wire n_6601;
wire n_8570;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_8579;
wire n_2111;
wire n_3743;
wire n_8079;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_8506;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_8291;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_1003;
wire n_7758;
wire n_8320;
wire n_8635;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_8375;
wire n_2973;
wire n_8612;
wire n_8778;
wire n_5893;
wire n_2710;
wire n_7705;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_8872;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_8006;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_8491;
wire n_8218;
wire n_1212;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_5726;
wire n_3933;
wire n_7439;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_7744;
wire n_3898;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_8240;
wire n_4749;
wire n_7707;
wire n_5924;
wire n_1845;
wire n_7733;
wire n_921;
wire n_5545;
wire n_8458;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_8853;
wire n_5083;
wire n_7684;
wire n_3253;
wire n_8306;
wire n_2088;
wire n_1275;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_904;
wire n_7673;
wire n_2005;
wire n_1696;
wire n_7187;
wire n_8013;
wire n_2108;
wire n_3824;
wire n_8342;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_6264;
wire n_5782;
wire n_8119;
wire n_4168;
wire n_1369;
wire n_8582;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_7931;
wire n_4743;
wire n_8445;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_8044;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_8363;
wire n_8464;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_7480;
wire n_8843;
wire n_5185;
wire n_8405;
wire n_2964;
wire n_8376;
wire n_5032;
wire n_6990;
wire n_865;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_1041;
wire n_2451;
wire n_8694;
wire n_2913;
wire n_8848;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_8752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_8625;
wire n_8894;
wire n_7380;
wire n_2839;
wire n_8813;
wire n_3237;
wire n_7708;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_8430;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_8770;
wire n_6277;
wire n_8426;
wire n_5115;
wire n_7376;
wire n_8411;
wire n_902;
wire n_8817;
wire n_8461;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_6409;
wire n_4095;
wire n_8391;
wire n_8507;
wire n_1310;
wire n_5927;
wire n_8691;
wire n_4485;
wire n_7657;
wire n_6388;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_4356;
wire n_3327;
wire n_1896;
wire n_6864;
wire n_1516;
wire n_4890;
wire n_8084;
wire n_8856;
wire n_2485;
wire n_6679;
wire n_8631;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_8219;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_7586;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_8428;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_8338;
wire n_1631;
wire n_7602;
wire n_6566;
wire n_1794;
wire n_5696;
wire n_7998;
wire n_8666;
wire n_5014;
wire n_1375;
wire n_3053;
wire n_7106;
wire n_6346;
wire n_7557;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_7026;
wire n_4335;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_7394;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_7627;
wire n_6436;
wire n_1464;
wire n_7719;
wire n_2798;
wire n_7450;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_7852;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_7462;
wire n_7780;
wire n_3503;
wire n_8523;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_7582;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_7555;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_8380;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_6612;
wire n_5258;

INVx1_ASAP7_75t_SL g849 ( 
.A(n_442),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_156),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_86),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_494),
.Y(n_852)
);

CKINVDCx11_ASAP7_75t_R g853 ( 
.A(n_35),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_526),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_527),
.Y(n_855)
);

CKINVDCx14_ASAP7_75t_R g856 ( 
.A(n_23),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_144),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_622),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_627),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_370),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_816),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_259),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_250),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_780),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_565),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_241),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_478),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_219),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_219),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_821),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_780),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_425),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_46),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_264),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_278),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_485),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_808),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_297),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_35),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_712),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_427),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_696),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_601),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_223),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_421),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_169),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_819),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_504),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_528),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_229),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_529),
.Y(n_891)
);

BUFx8_ASAP7_75t_SL g892 ( 
.A(n_467),
.Y(n_892)
);

CKINVDCx20_ASAP7_75t_R g893 ( 
.A(n_699),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_9),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_622),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_651),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_428),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_792),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_555),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_684),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_835),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_156),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_792),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_644),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_528),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_659),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_794),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_60),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_559),
.Y(n_909)
);

BUFx10_ASAP7_75t_L g910 ( 
.A(n_381),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_137),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_113),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_72),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_717),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_517),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_669),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_353),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_225),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_481),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_714),
.Y(n_920)
);

INVxp67_ASAP7_75t_SL g921 ( 
.A(n_448),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_831),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_547),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_629),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_487),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_833),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_187),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_237),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_210),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_506),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_547),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_837),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_71),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_33),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_810),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_597),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_166),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_650),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_380),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_804),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_159),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_518),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_55),
.Y(n_943)
);

BUFx10_ASAP7_75t_L g944 ( 
.A(n_398),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_629),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_543),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_769),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_416),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_208),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_338),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_62),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_363),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_236),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_462),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_678),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_405),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_191),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_700),
.Y(n_958)
);

BUFx10_ASAP7_75t_L g959 ( 
.A(n_28),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_803),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_737),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_267),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_16),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_63),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_313),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_345),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_830),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_686),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_138),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_243),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_655),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_254),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_685),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_154),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_427),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_222),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_408),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_461),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_381),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_584),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_105),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_460),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_167),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_325),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_499),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_750),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_236),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_38),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_723),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_725),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_679),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_820),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_473),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_78),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_504),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_457),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_497),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_345),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_272),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_710),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_597),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_731),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_75),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_660),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_197),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_150),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_308),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_582),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_848),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_49),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_230),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_571),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_452),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_404),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_571),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_82),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_400),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_491),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_337),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_362),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_632),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_701),
.Y(n_1022)
);

BUFx10_ASAP7_75t_L g1023 ( 
.A(n_220),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_841),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_592),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_519),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_623),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_678),
.Y(n_1028)
);

INVx1_ASAP7_75t_SL g1029 ( 
.A(n_22),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_446),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_749),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_512),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_575),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_201),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_7),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_84),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_409),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_544),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_830),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_269),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_687),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_823),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_50),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_415),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_160),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_385),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_614),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_250),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_824),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_581),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_595),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_457),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_248),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_383),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_147),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_144),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_506),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_157),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_89),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_478),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_350),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_433),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_166),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_569),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_265),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_383),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_114),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_101),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_407),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_729),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_313),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_242),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_372),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_644),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_561),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_443),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_170),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_80),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_56),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_658),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_367),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_180),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_612),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_2),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_771),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_132),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_602),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_812),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_433),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_603),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_196),
.Y(n_1091)
);

INVx1_ASAP7_75t_SL g1092 ( 
.A(n_303),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_13),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_13),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_163),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_331),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_155),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_560),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_472),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_618),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_197),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_668),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_99),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_783),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_272),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_589),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_543),
.Y(n_1107)
);

BUFx5_ASAP7_75t_L g1108 ( 
.A(n_414),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_823),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_261),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_318),
.Y(n_1111)
);

CKINVDCx20_ASAP7_75t_R g1112 ( 
.A(n_245),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_831),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_350),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_799),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_502),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_580),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_186),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_22),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_773),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_663),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_261),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_704),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_577),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_439),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_611),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_23),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_694),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_568),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_782),
.Y(n_1130)
);

CKINVDCx20_ASAP7_75t_R g1131 ( 
.A(n_690),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_443),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_627),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_630),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_104),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_435),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_610),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_208),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_63),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_210),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_122),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_570),
.Y(n_1142)
);

INVxp67_ASAP7_75t_L g1143 ( 
.A(n_406),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_709),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_727),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_784),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_665),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_367),
.Y(n_1148)
);

BUFx3_ASAP7_75t_L g1149 ( 
.A(n_380),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_656),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_278),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_568),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_199),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_808),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_97),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_333),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_164),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_95),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_411),
.Y(n_1159)
);

BUFx10_ASAP7_75t_L g1160 ( 
.A(n_758),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_114),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_760),
.Y(n_1162)
);

BUFx5_ASAP7_75t_L g1163 ( 
.A(n_558),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_196),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_227),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_208),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_784),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_276),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_106),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_446),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_413),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_654),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_196),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_88),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_261),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_767),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_17),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_451),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_573),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_459),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_716),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_635),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_296),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_179),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_39),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_85),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_625),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_492),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_624),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_769),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_417),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_688),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_307),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_467),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_408),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_369),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_612),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_54),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_63),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_255),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_474),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_38),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_162),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_42),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_189),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_742),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_286),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_482),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_306),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_186),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_44),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_262),
.Y(n_1212)
);

CKINVDCx14_ASAP7_75t_R g1213 ( 
.A(n_412),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_562),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_753),
.Y(n_1215)
);

CKINVDCx16_ASAP7_75t_R g1216 ( 
.A(n_666),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_124),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_795),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_604),
.Y(n_1219)
);

BUFx10_ASAP7_75t_L g1220 ( 
.A(n_786),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_393),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_779),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_296),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_186),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_358),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_252),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_240),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_848),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_368),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_602),
.Y(n_1230)
);

INVx1_ASAP7_75t_SL g1231 ( 
.A(n_797),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_164),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_217),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_228),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_729),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_470),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_664),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_298),
.Y(n_1238)
);

CKINVDCx20_ASAP7_75t_R g1239 ( 
.A(n_588),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_768),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_730),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_89),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_445),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_280),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_673),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_834),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_289),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_45),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_143),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_567),
.Y(n_1250)
);

CKINVDCx16_ASAP7_75t_R g1251 ( 
.A(n_663),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_521),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_704),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_406),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_257),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_456),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_172),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_31),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_139),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_356),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_649),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_601),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_93),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_189),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_532),
.Y(n_1265)
);

CKINVDCx14_ASAP7_75t_R g1266 ( 
.A(n_470),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_36),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_41),
.Y(n_1268)
);

CKINVDCx16_ASAP7_75t_R g1269 ( 
.A(n_586),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_128),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_548),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_137),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_518),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_379),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_356),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_621),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_107),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_529),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_34),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_605),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_331),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_590),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_174),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_343),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_426),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_763),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_272),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_292),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_321),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_68),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_378),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_32),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_316),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_184),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_39),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_565),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_184),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_429),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_65),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_452),
.Y(n_1300)
);

INVx1_ASAP7_75t_SL g1301 ( 
.A(n_458),
.Y(n_1301)
);

INVx2_ASAP7_75t_SL g1302 ( 
.A(n_458),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_134),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_788),
.Y(n_1304)
);

BUFx8_ASAP7_75t_SL g1305 ( 
.A(n_834),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_123),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_212),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_92),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_273),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_39),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_501),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_548),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_556),
.Y(n_1313)
);

BUFx10_ASAP7_75t_L g1314 ( 
.A(n_8),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_696),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_114),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_822),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_723),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_322),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_786),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_605),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_113),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_373),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_349),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_762),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_525),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_697),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_596),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_643),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_579),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_531),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_803),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_268),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_722),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_788),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_728),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_656),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_50),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_74),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_634),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_400),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_546),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_407),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_82),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_416),
.Y(n_1345)
);

CKINVDCx14_ASAP7_75t_R g1346 ( 
.A(n_664),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_778),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_60),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_642),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_239),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_126),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_0),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_717),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_76),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_789),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_782),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_647),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_307),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_171),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_58),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_741),
.Y(n_1361)
);

CKINVDCx14_ASAP7_75t_R g1362 ( 
.A(n_14),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_34),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_14),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_666),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_471),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_57),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_635),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_640),
.Y(n_1369)
);

BUFx8_ASAP7_75t_SL g1370 ( 
.A(n_420),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_166),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_465),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_639),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_224),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_662),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_787),
.Y(n_1376)
);

CKINVDCx16_ASAP7_75t_R g1377 ( 
.A(n_263),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_78),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_209),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_317),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_450),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_184),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_231),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_677),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_357),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_670),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_355),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_159),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_31),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_172),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_352),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_498),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_747),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_549),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_698),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_713),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_370),
.Y(n_1397)
);

BUFx5_ASAP7_75t_L g1398 ( 
.A(n_376),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_5),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_542),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_694),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_532),
.Y(n_1402)
);

CKINVDCx16_ASAP7_75t_R g1403 ( 
.A(n_495),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_336),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_842),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_262),
.Y(n_1406)
);

CKINVDCx20_ASAP7_75t_R g1407 ( 
.A(n_48),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_29),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_394),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_16),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_844),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_56),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_475),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_97),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_33),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_3),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_397),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_153),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_520),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_344),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_70),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_495),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_200),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_735),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_607),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_519),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_21),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_410),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_560),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_447),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_615),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_659),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_749),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_683),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_336),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_132),
.Y(n_1436)
);

BUFx8_ASAP7_75t_SL g1437 ( 
.A(n_464),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_250),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_18),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_730),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_167),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_185),
.Y(n_1442)
);

BUFx6f_ASAP7_75t_L g1443 ( 
.A(n_750),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_402),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_139),
.Y(n_1445)
);

CKINVDCx16_ASAP7_75t_R g1446 ( 
.A(n_480),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_785),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_399),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_6),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_140),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_583),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_812),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_776),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_474),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_684),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_288),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_216),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_94),
.Y(n_1458)
);

CKINVDCx14_ASAP7_75t_R g1459 ( 
.A(n_551),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_5),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_403),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_600),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_731),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_129),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_793),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_459),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_195),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_181),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1213),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_852),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1406),
.B(n_0),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_894),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1213),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1266),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1067),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1067),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_864),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1067),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1266),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1346),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_864),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_894),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1346),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1459),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1097),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1459),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1108),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_892),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1097),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_894),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1097),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1258),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1258),
.Y(n_1493)
);

CKINVDCx16_ASAP7_75t_R g1494 ( 
.A(n_856),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1258),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1173),
.B(n_0),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_892),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1406),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1305),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1305),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_1370),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1370),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1437),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1437),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1406),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_894),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_856),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1406),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_894),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1362),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1362),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_929),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_853),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_853),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_863),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1216),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_929),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1216),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1376),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1376),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1251),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1376),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_894),
.Y(n_1523)
);

CKINVDCx20_ASAP7_75t_R g1524 ( 
.A(n_888),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1376),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_1251),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1269),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_855),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1108),
.Y(n_1529)
);

BUFx10_ASAP7_75t_L g1530 ( 
.A(n_894),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_855),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_855),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1269),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1403),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_885),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_885),
.Y(n_1536)
);

NOR2xp67_ASAP7_75t_L g1537 ( 
.A(n_1091),
.B(n_1),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_1403),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1446),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1446),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_852),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1108),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_1377),
.Y(n_1543)
);

NOR2xp67_ASAP7_75t_L g1544 ( 
.A(n_1091),
.B(n_1),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1466),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_854),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_860),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_861),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_885),
.Y(n_1549)
);

NOR2xp67_ASAP7_75t_L g1550 ( 
.A(n_1091),
.B(n_1),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_896),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_896),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1377),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_896),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_981),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1463),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1465),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_930),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_865),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_863),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_867),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_930),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1173),
.B(n_2),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_930),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_934),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_876),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_877),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_981),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1144),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1144),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_888),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_864),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_881),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_887),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1144),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1176),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1149),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_981),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1451),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1452),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_981),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_864),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_934),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1149),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1149),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_959),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1176),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_889),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_893),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1029),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1181),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1181),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1181),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1155),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_981),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_895),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_898),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1155),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1342),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1155),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1287),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_893),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_901),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1287),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_904),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1287),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_873),
.Y(n_1607)
);

BUFx10_ASAP7_75t_L g1608 ( 
.A(n_981),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_873),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_873),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_962),
.Y(n_1611)
);

BUFx10_ASAP7_75t_L g1612 ( 
.A(n_981),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_906),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_962),
.Y(n_1614)
);

BUFx2_ASAP7_75t_SL g1615 ( 
.A(n_959),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_907),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_909),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_962),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1019),
.Y(n_1619)
);

XOR2xp5_ASAP7_75t_L g1620 ( 
.A(n_1468),
.B(n_943),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_914),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_900),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1019),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1135),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1019),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1141),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1141),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1141),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_917),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1158),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1029),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1158),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1158),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1279),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1279),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_864),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1279),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1135),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1108),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1135),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_919),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1316),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1316),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_920),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1135),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_900),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1108),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1316),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1367),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1342),
.Y(n_1650)
);

BUFx10_ASAP7_75t_L g1651 ( 
.A(n_1135),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1367),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1367),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1382),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1382),
.Y(n_1655)
);

CKINVDCx20_ASAP7_75t_R g1656 ( 
.A(n_925),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1382),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1289),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_922),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1289),
.Y(n_1660)
);

INVxp67_ASAP7_75t_L g1661 ( 
.A(n_1356),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1012),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1108),
.B(n_2),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_923),
.Y(n_1664)
);

INVxp67_ASAP7_75t_SL g1665 ( 
.A(n_1135),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_924),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_926),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_935),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_936),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1012),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_925),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_939),
.Y(n_1672)
);

INVx1_ASAP7_75t_SL g1673 ( 
.A(n_1092),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1098),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1108),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1012),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_864),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_864),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1042),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_931),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_940),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1135),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1199),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1042),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1042),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1047),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1047),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1047),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_931),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1199),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1182),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1182),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1182),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1098),
.B(n_3),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1302),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1302),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1302),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_942),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1199),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_938),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1199),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_945),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_959),
.Y(n_1703)
);

CKINVDCx14_ASAP7_75t_R g1704 ( 
.A(n_959),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_948),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_938),
.Y(n_1706)
);

INVxp33_ASAP7_75t_SL g1707 ( 
.A(n_1356),
.Y(n_1707)
);

BUFx2_ASAP7_75t_L g1708 ( 
.A(n_1188),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_956),
.Y(n_1709)
);

INVx4_ASAP7_75t_R g1710 ( 
.A(n_1092),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1199),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_958),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_955),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1199),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1365),
.B(n_3),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_960),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1199),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1264),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_961),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1108),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1264),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_966),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1264),
.Y(n_1723)
);

BUFx10_ASAP7_75t_L g1724 ( 
.A(n_1264),
.Y(n_1724)
);

INVxp33_ASAP7_75t_L g1725 ( 
.A(n_1365),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_955),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1264),
.Y(n_1727)
);

CKINVDCx20_ASAP7_75t_R g1728 ( 
.A(n_989),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1264),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1264),
.Y(n_1730)
);

CKINVDCx16_ASAP7_75t_R g1731 ( 
.A(n_1023),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1259),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1023),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1295),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_967),
.Y(n_1735)
);

BUFx5_ASAP7_75t_L g1736 ( 
.A(n_851),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1295),
.Y(n_1737)
);

BUFx2_ASAP7_75t_SL g1738 ( 
.A(n_1023),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1295),
.Y(n_1739)
);

CKINVDCx16_ASAP7_75t_R g1740 ( 
.A(n_1023),
.Y(n_1740)
);

BUFx5_ASAP7_75t_L g1741 ( 
.A(n_851),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_968),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_971),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1108),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1295),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_973),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1188),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1295),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_989),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1295),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_903),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1295),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1360),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_975),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1360),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1360),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_977),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_982),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1360),
.Y(n_1759)
);

BUFx3_ASAP7_75t_L g1760 ( 
.A(n_1108),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_985),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1360),
.Y(n_1762)
);

BUFx3_ASAP7_75t_L g1763 ( 
.A(n_1163),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1360),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_986),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_903),
.Y(n_1766)
);

CKINVDCx16_ASAP7_75t_R g1767 ( 
.A(n_1314),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_993),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1360),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1412),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_995),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1412),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1412),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1412),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1412),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1412),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_998),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1412),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_857),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_857),
.Y(n_1780)
);

BUFx6f_ASAP7_75t_L g1781 ( 
.A(n_903),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1163),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_879),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_879),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_884),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1163),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_884),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_886),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1001),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1008),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_886),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_890),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_890),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_912),
.Y(n_1794)
);

CKINVDCx5p33_ASAP7_75t_R g1795 ( 
.A(n_1013),
.Y(n_1795)
);

BUFx3_ASAP7_75t_L g1796 ( 
.A(n_1163),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1422),
.Y(n_1797)
);

CKINVDCx5p33_ASAP7_75t_R g1798 ( 
.A(n_1014),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1422),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_997),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_912),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_913),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_913),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1015),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1017),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_933),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_933),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1163),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1163),
.Y(n_1809)
);

CKINVDCx20_ASAP7_75t_R g1810 ( 
.A(n_997),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1018),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1424),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1424),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_937),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1163),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_937),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_969),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_969),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1024),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1163),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_972),
.Y(n_1821)
);

BUFx3_ASAP7_75t_L g1822 ( 
.A(n_1163),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1163),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1025),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_L g1825 ( 
.A(n_903),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_972),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_976),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1026),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1398),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_976),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_988),
.Y(n_1831)
);

CKINVDCx20_ASAP7_75t_R g1832 ( 
.A(n_1064),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_988),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1005),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1005),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_943),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1028),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1035),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1035),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_850),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1036),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_1030),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1036),
.Y(n_1843)
);

BUFx3_ASAP7_75t_L g1844 ( 
.A(n_1398),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1064),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_1031),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1039),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1043),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1398),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1044),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_862),
.Y(n_1851)
);

BUFx5_ASAP7_75t_L g1852 ( 
.A(n_1043),
.Y(n_1852)
);

INVx2_ASAP7_75t_SL g1853 ( 
.A(n_1314),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1046),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1050),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1045),
.Y(n_1856)
);

BUFx3_ASAP7_75t_L g1857 ( 
.A(n_1398),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1052),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1045),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1057),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1055),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1062),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1055),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1056),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1069),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1398),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1070),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1073),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1074),
.Y(n_1869)
);

CKINVDCx20_ASAP7_75t_R g1870 ( 
.A(n_1126),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1398),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1126),
.Y(n_1872)
);

CKINVDCx20_ASAP7_75t_R g1873 ( 
.A(n_1131),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1011),
.Y(n_1874)
);

CKINVDCx20_ASAP7_75t_R g1875 ( 
.A(n_1131),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1056),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1076),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_903),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1398),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1080),
.Y(n_1880)
);

CKINVDCx16_ASAP7_75t_R g1881 ( 
.A(n_1314),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1081),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1063),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1063),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1083),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1087),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1398),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1088),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1089),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1398),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1100),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1147),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1102),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1072),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1147),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1072),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1398),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1104),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1078),
.Y(n_1899)
);

CKINVDCx20_ASAP7_75t_R g1900 ( 
.A(n_1148),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1078),
.Y(n_1901)
);

CKINVDCx16_ASAP7_75t_R g1902 ( 
.A(n_1314),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1084),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1106),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1084),
.Y(n_1905)
);

CKINVDCx5p33_ASAP7_75t_R g1906 ( 
.A(n_1109),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1096),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1114),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1116),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1148),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_903),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1117),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1123),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1124),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1096),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1105),
.Y(n_1916)
);

CKINVDCx5p33_ASAP7_75t_R g1917 ( 
.A(n_1129),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1105),
.Y(n_1918)
);

CKINVDCx16_ASAP7_75t_R g1919 ( 
.A(n_910),
.Y(n_1919)
);

CKINVDCx16_ASAP7_75t_R g1920 ( 
.A(n_910),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1130),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1118),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1118),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1119),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1119),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1139),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1139),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1156),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1156),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_1133),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_903),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1174),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1134),
.Y(n_1933)
);

CKINVDCx16_ASAP7_75t_R g1934 ( 
.A(n_910),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1136),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1174),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_866),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1203),
.B(n_4),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1150),
.Y(n_1939)
);

CKINVDCx5p33_ASAP7_75t_R g1940 ( 
.A(n_1152),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1203),
.Y(n_1941)
);

NOR2xp67_ASAP7_75t_L g1942 ( 
.A(n_1040),
.B(n_4),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1204),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1204),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1205),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1154),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1205),
.Y(n_1947)
);

CKINVDCx16_ASAP7_75t_R g1948 ( 
.A(n_910),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_991),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1207),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1162),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1167),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1171),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1172),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1179),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1207),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1211),
.Y(n_1957)
);

INVxp67_ASAP7_75t_L g1958 ( 
.A(n_921),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1211),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1217),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1217),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_868),
.Y(n_1962)
);

CKINVDCx5p33_ASAP7_75t_R g1963 ( 
.A(n_1180),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1223),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1159),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1223),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1187),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1189),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_944),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1159),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1190),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1249),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1249),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1255),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_991),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1255),
.Y(n_1976)
);

BUFx6f_ASAP7_75t_L g1977 ( 
.A(n_991),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1192),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1194),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1257),
.Y(n_1980)
);

CKINVDCx20_ASAP7_75t_R g1981 ( 
.A(n_1240),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1257),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_991),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1011),
.Y(n_1984)
);

INVxp33_ASAP7_75t_L g1985 ( 
.A(n_870),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1263),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1263),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1267),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1267),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1240),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_991),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_944),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1270),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1270),
.Y(n_1994)
);

CKINVDCx16_ASAP7_75t_R g1995 ( 
.A(n_944),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1195),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1196),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1277),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_1197),
.Y(n_1999)
);

NOR2xp67_ASAP7_75t_L g2000 ( 
.A(n_1040),
.B(n_4),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_1488),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1498),
.Y(n_2002)
);

INVxp33_ASAP7_75t_SL g2003 ( 
.A(n_1513),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1505),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1508),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1519),
.Y(n_2006)
);

CKINVDCx20_ASAP7_75t_R g2007 ( 
.A(n_1524),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1520),
.Y(n_2008)
);

CKINVDCx16_ASAP7_75t_R g2009 ( 
.A(n_1494),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1522),
.Y(n_2010)
);

INVxp67_ASAP7_75t_SL g2011 ( 
.A(n_1665),
.Y(n_2011)
);

INVxp67_ASAP7_75t_SL g2012 ( 
.A(n_1729),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1525),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1488),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1594),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1598),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1600),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1601),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1604),
.Y(n_2019)
);

INVxp67_ASAP7_75t_SL g2020 ( 
.A(n_1778),
.Y(n_2020)
);

INVxp67_ASAP7_75t_SL g2021 ( 
.A(n_1487),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1606),
.Y(n_2022)
);

INVxp67_ASAP7_75t_SL g2023 ( 
.A(n_1487),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1662),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1499),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1670),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1499),
.Y(n_2027)
);

CKINVDCx16_ASAP7_75t_R g2028 ( 
.A(n_1586),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1676),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1501),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1571),
.Y(n_2031)
);

INVxp33_ASAP7_75t_L g2032 ( 
.A(n_1512),
.Y(n_2032)
);

INVx1_ASAP7_75t_SL g2033 ( 
.A(n_1515),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1472),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1472),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1679),
.Y(n_2036)
);

CKINVDCx5p33_ASAP7_75t_R g2037 ( 
.A(n_1501),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1684),
.Y(n_2038)
);

CKINVDCx16_ASAP7_75t_R g2039 ( 
.A(n_1731),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1685),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1502),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1482),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1686),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_1589),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1502),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1687),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1688),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_1602),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_1560),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_1516),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1691),
.Y(n_2051)
);

CKINVDCx20_ASAP7_75t_R g2052 ( 
.A(n_1622),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1692),
.Y(n_2053)
);

INVxp67_ASAP7_75t_L g2054 ( 
.A(n_1565),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1503),
.Y(n_2055)
);

INVxp67_ASAP7_75t_SL g2056 ( 
.A(n_1529),
.Y(n_2056)
);

INVxp67_ASAP7_75t_SL g2057 ( 
.A(n_1529),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1503),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1693),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1695),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1704),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1482),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1696),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_1646),
.Y(n_2064)
);

INVxp33_ASAP7_75t_L g2065 ( 
.A(n_1517),
.Y(n_2065)
);

CKINVDCx20_ASAP7_75t_R g2066 ( 
.A(n_1656),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1697),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1490),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1497),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1500),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1528),
.Y(n_2071)
);

INVxp67_ASAP7_75t_SL g2072 ( 
.A(n_1542),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1531),
.Y(n_2073)
);

INVxp67_ASAP7_75t_SL g2074 ( 
.A(n_1542),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1532),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1535),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1536),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1549),
.Y(n_2078)
);

INVxp67_ASAP7_75t_SL g2079 ( 
.A(n_1639),
.Y(n_2079)
);

INVxp33_ASAP7_75t_L g2080 ( 
.A(n_1553),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1551),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_1583),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1552),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1554),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1558),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1562),
.Y(n_2086)
);

INVxp67_ASAP7_75t_SL g2087 ( 
.A(n_1639),
.Y(n_2087)
);

BUFx2_ASAP7_75t_L g2088 ( 
.A(n_1516),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1564),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1569),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1490),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1570),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_1504),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1575),
.Y(n_2094)
);

INVxp33_ASAP7_75t_SL g2095 ( 
.A(n_1513),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_1647),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1577),
.Y(n_2097)
);

HB1xp67_ASAP7_75t_L g2098 ( 
.A(n_1590),
.Y(n_2098)
);

CKINVDCx20_ASAP7_75t_R g2099 ( 
.A(n_1671),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1584),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1585),
.Y(n_2101)
);

INVxp33_ASAP7_75t_SL g2102 ( 
.A(n_1514),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1591),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1592),
.Y(n_2104)
);

CKINVDCx20_ASAP7_75t_R g2105 ( 
.A(n_1680),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1545),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_1631),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1593),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1663),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1545),
.Y(n_2110)
);

CKINVDCx16_ASAP7_75t_R g2111 ( 
.A(n_1733),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1787),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1859),
.Y(n_2113)
);

INVxp67_ASAP7_75t_SL g2114 ( 
.A(n_1647),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1546),
.Y(n_2115)
);

CKINVDCx20_ASAP7_75t_R g2116 ( 
.A(n_1689),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1475),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1673),
.Y(n_2118)
);

CKINVDCx20_ASAP7_75t_R g2119 ( 
.A(n_1700),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1546),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1476),
.Y(n_2121)
);

CKINVDCx20_ASAP7_75t_R g2122 ( 
.A(n_1706),
.Y(n_2122)
);

CKINVDCx16_ASAP7_75t_R g2123 ( 
.A(n_1740),
.Y(n_2123)
);

BUFx2_ASAP7_75t_SL g2124 ( 
.A(n_1484),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1547),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1547),
.Y(n_2126)
);

INVxp33_ASAP7_75t_L g2127 ( 
.A(n_1840),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1478),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_1548),
.Y(n_2129)
);

INVxp67_ASAP7_75t_SL g2130 ( 
.A(n_1675),
.Y(n_2130)
);

INVxp67_ASAP7_75t_SL g2131 ( 
.A(n_1675),
.Y(n_2131)
);

INVxp67_ASAP7_75t_SL g2132 ( 
.A(n_1720),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_1732),
.Y(n_2133)
);

INVxp67_ASAP7_75t_SL g2134 ( 
.A(n_1720),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_1548),
.Y(n_2135)
);

INVxp33_ASAP7_75t_SL g2136 ( 
.A(n_1514),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_1556),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1485),
.Y(n_2138)
);

INVxp67_ASAP7_75t_SL g2139 ( 
.A(n_1744),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1506),
.Y(n_2140)
);

CKINVDCx20_ASAP7_75t_R g2141 ( 
.A(n_1713),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1489),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1491),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1492),
.Y(n_2144)
);

CKINVDCx16_ASAP7_75t_R g2145 ( 
.A(n_1767),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1477),
.Y(n_2146)
);

INVxp67_ASAP7_75t_L g2147 ( 
.A(n_1615),
.Y(n_2147)
);

CKINVDCx20_ASAP7_75t_R g2148 ( 
.A(n_1726),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1493),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1506),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1495),
.Y(n_2151)
);

CKINVDCx20_ASAP7_75t_R g2152 ( 
.A(n_1728),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1779),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1780),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1556),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1783),
.Y(n_2156)
);

CKINVDCx16_ASAP7_75t_R g2157 ( 
.A(n_1881),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1557),
.Y(n_2158)
);

INVx3_ASAP7_75t_L g2159 ( 
.A(n_1530),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1784),
.Y(n_2160)
);

CKINVDCx20_ASAP7_75t_R g2161 ( 
.A(n_1749),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1785),
.Y(n_2162)
);

CKINVDCx20_ASAP7_75t_R g2163 ( 
.A(n_1800),
.Y(n_2163)
);

CKINVDCx5p33_ASAP7_75t_R g2164 ( 
.A(n_1557),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1559),
.Y(n_2165)
);

CKINVDCx16_ASAP7_75t_R g2166 ( 
.A(n_1902),
.Y(n_2166)
);

CKINVDCx20_ASAP7_75t_R g2167 ( 
.A(n_1810),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1788),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1791),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1792),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1793),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1794),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1801),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1802),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1559),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1803),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_1543),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_1744),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1806),
.Y(n_2179)
);

CKINVDCx20_ASAP7_75t_R g2180 ( 
.A(n_1832),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1807),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1760),
.Y(n_2182)
);

INVxp67_ASAP7_75t_SL g2183 ( 
.A(n_1760),
.Y(n_2183)
);

INVxp33_ASAP7_75t_L g2184 ( 
.A(n_1851),
.Y(n_2184)
);

CKINVDCx20_ASAP7_75t_R g2185 ( 
.A(n_1845),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1814),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1816),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1817),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1818),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1821),
.Y(n_2190)
);

CKINVDCx20_ASAP7_75t_R g2191 ( 
.A(n_1870),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1826),
.Y(n_2192)
);

CKINVDCx5p33_ASAP7_75t_R g2193 ( 
.A(n_1561),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1827),
.Y(n_2194)
);

CKINVDCx20_ASAP7_75t_R g2195 ( 
.A(n_1872),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1830),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1831),
.Y(n_2197)
);

CKINVDCx20_ASAP7_75t_R g2198 ( 
.A(n_1873),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1833),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1834),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1835),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1838),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1839),
.Y(n_2203)
);

INVxp67_ASAP7_75t_SL g2204 ( 
.A(n_1763),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1841),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1561),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1843),
.Y(n_2207)
);

CKINVDCx5p33_ASAP7_75t_R g2208 ( 
.A(n_1566),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1848),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1856),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1861),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1863),
.Y(n_2212)
);

INVxp67_ASAP7_75t_L g2213 ( 
.A(n_1738),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1864),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1876),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1883),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1884),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1894),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1896),
.Y(n_2219)
);

INVxp67_ASAP7_75t_SL g2220 ( 
.A(n_1763),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1899),
.Y(n_2221)
);

BUFx2_ASAP7_75t_SL g2222 ( 
.A(n_1507),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1566),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1901),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1509),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1903),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1905),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1907),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1915),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1916),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1918),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1922),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1923),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1924),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1509),
.Y(n_2235)
);

CKINVDCx20_ASAP7_75t_R g2236 ( 
.A(n_1875),
.Y(n_2236)
);

INVx1_ASAP7_75t_SL g2237 ( 
.A(n_1510),
.Y(n_2237)
);

CKINVDCx20_ASAP7_75t_R g2238 ( 
.A(n_1892),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_1469),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1925),
.Y(n_2240)
);

INVxp67_ASAP7_75t_L g2241 ( 
.A(n_1937),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_1567),
.Y(n_2242)
);

INVxp33_ASAP7_75t_SL g2243 ( 
.A(n_1469),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_1926),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1927),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1928),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_1567),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1523),
.Y(n_2248)
);

CKINVDCx5p33_ASAP7_75t_R g2249 ( 
.A(n_1573),
.Y(n_2249)
);

CKINVDCx5p33_ASAP7_75t_R g2250 ( 
.A(n_1573),
.Y(n_2250)
);

CKINVDCx20_ASAP7_75t_R g2251 ( 
.A(n_1895),
.Y(n_2251)
);

CKINVDCx20_ASAP7_75t_R g2252 ( 
.A(n_1900),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1929),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1932),
.Y(n_2254)
);

INVx1_ASAP7_75t_SL g2255 ( 
.A(n_1518),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1936),
.Y(n_2256)
);

CKINVDCx5p33_ASAP7_75t_R g2257 ( 
.A(n_1574),
.Y(n_2257)
);

CKINVDCx20_ASAP7_75t_R g2258 ( 
.A(n_1910),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1941),
.Y(n_2259)
);

CKINVDCx20_ASAP7_75t_R g2260 ( 
.A(n_1965),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1943),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_1518),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1944),
.Y(n_2263)
);

CKINVDCx16_ASAP7_75t_R g2264 ( 
.A(n_1919),
.Y(n_2264)
);

CKINVDCx20_ASAP7_75t_R g2265 ( 
.A(n_1970),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1945),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_1477),
.Y(n_2267)
);

CKINVDCx20_ASAP7_75t_R g2268 ( 
.A(n_1981),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_1962),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1947),
.Y(n_2270)
);

CKINVDCx20_ASAP7_75t_R g2271 ( 
.A(n_1990),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1950),
.Y(n_2272)
);

INVxp67_ASAP7_75t_SL g2273 ( 
.A(n_1796),
.Y(n_2273)
);

INVxp67_ASAP7_75t_L g2274 ( 
.A(n_1674),
.Y(n_2274)
);

INVxp33_ASAP7_75t_SL g2275 ( 
.A(n_1473),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1956),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1957),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1959),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_1574),
.Y(n_2279)
);

CKINVDCx16_ASAP7_75t_R g2280 ( 
.A(n_1920),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_1521),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1960),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1961),
.Y(n_2283)
);

CKINVDCx5p33_ASAP7_75t_R g2284 ( 
.A(n_1579),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1964),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1966),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1972),
.Y(n_2287)
);

INVxp67_ASAP7_75t_SL g2288 ( 
.A(n_1796),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1973),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1974),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1976),
.Y(n_2291)
);

INVxp67_ASAP7_75t_SL g2292 ( 
.A(n_1822),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1980),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1982),
.Y(n_2294)
);

INVxp67_ASAP7_75t_SL g2295 ( 
.A(n_1822),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1986),
.Y(n_2296)
);

CKINVDCx20_ASAP7_75t_R g2297 ( 
.A(n_1620),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1523),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1987),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1988),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_1579),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1989),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1993),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1994),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1998),
.Y(n_2305)
);

CKINVDCx20_ASAP7_75t_R g2306 ( 
.A(n_1934),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1471),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_1580),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1736),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1736),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1736),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1736),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1736),
.Y(n_2313)
);

INVxp67_ASAP7_75t_SL g2314 ( 
.A(n_1844),
.Y(n_2314)
);

CKINVDCx20_ASAP7_75t_R g2315 ( 
.A(n_1948),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1736),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_1844),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1555),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1736),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_1473),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1736),
.Y(n_2321)
);

INVxp67_ASAP7_75t_L g2322 ( 
.A(n_1708),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_1474),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1555),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1741),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_1474),
.Y(n_2326)
);

INVxp67_ASAP7_75t_SL g2327 ( 
.A(n_1857),
.Y(n_2327)
);

CKINVDCx20_ASAP7_75t_R g2328 ( 
.A(n_1995),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_1479),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1741),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1741),
.Y(n_2331)
);

CKINVDCx20_ASAP7_75t_R g2332 ( 
.A(n_1836),
.Y(n_2332)
);

CKINVDCx16_ASAP7_75t_R g2333 ( 
.A(n_1703),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1741),
.Y(n_2334)
);

INVxp67_ASAP7_75t_L g2335 ( 
.A(n_1797),
.Y(n_2335)
);

CKINVDCx16_ASAP7_75t_R g2336 ( 
.A(n_1703),
.Y(n_2336)
);

CKINVDCx20_ASAP7_75t_R g2337 ( 
.A(n_1874),
.Y(n_2337)
);

CKINVDCx16_ASAP7_75t_R g2338 ( 
.A(n_1853),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1741),
.Y(n_2339)
);

CKINVDCx5p33_ASAP7_75t_R g2340 ( 
.A(n_1479),
.Y(n_2340)
);

BUFx2_ASAP7_75t_L g2341 ( 
.A(n_1521),
.Y(n_2341)
);

CKINVDCx20_ASAP7_75t_R g2342 ( 
.A(n_1984),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_1480),
.Y(n_2343)
);

CKINVDCx20_ASAP7_75t_R g2344 ( 
.A(n_1984),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_1480),
.Y(n_2345)
);

CKINVDCx16_ASAP7_75t_R g2346 ( 
.A(n_1853),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_1483),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1741),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_1568),
.Y(n_2349)
);

INVxp67_ASAP7_75t_SL g2350 ( 
.A(n_1857),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1568),
.Y(n_2351)
);

INVxp67_ASAP7_75t_L g2352 ( 
.A(n_1812),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_1483),
.Y(n_2353)
);

CKINVDCx16_ASAP7_75t_R g2354 ( 
.A(n_1812),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1741),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1741),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_1852),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1852),
.Y(n_2358)
);

CKINVDCx20_ASAP7_75t_R g2359 ( 
.A(n_1526),
.Y(n_2359)
);

CKINVDCx20_ASAP7_75t_R g2360 ( 
.A(n_1526),
.Y(n_2360)
);

CKINVDCx20_ASAP7_75t_R g2361 ( 
.A(n_1527),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1852),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1852),
.Y(n_2363)
);

CKINVDCx20_ASAP7_75t_R g2364 ( 
.A(n_1527),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_1852),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_1533),
.Y(n_2366)
);

CKINVDCx16_ASAP7_75t_R g2367 ( 
.A(n_1969),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1578),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1852),
.Y(n_2369)
);

INVxp67_ASAP7_75t_L g2370 ( 
.A(n_1969),
.Y(n_2370)
);

INVxp33_ASAP7_75t_L g2371 ( 
.A(n_1725),
.Y(n_2371)
);

INVxp67_ASAP7_75t_L g2372 ( 
.A(n_1992),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_1852),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1852),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_1607),
.Y(n_2375)
);

HB1xp67_ASAP7_75t_L g2376 ( 
.A(n_1533),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1578),
.Y(n_2377)
);

INVxp67_ASAP7_75t_L g2378 ( 
.A(n_1992),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1609),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_1486),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1610),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_1534),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1611),
.Y(n_2383)
);

CKINVDCx5p33_ASAP7_75t_R g2384 ( 
.A(n_1486),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1614),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1618),
.Y(n_2386)
);

INVxp67_ASAP7_75t_SL g2387 ( 
.A(n_1983),
.Y(n_2387)
);

BUFx2_ASAP7_75t_L g2388 ( 
.A(n_1534),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1619),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1623),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_1625),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1626),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_1580),
.Y(n_2393)
);

AND2x6_ASAP7_75t_L g2394 ( 
.A(n_1581),
.B(n_858),
.Y(n_2394)
);

CKINVDCx20_ASAP7_75t_R g2395 ( 
.A(n_1538),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1627),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1628),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1630),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_1538),
.Y(n_2399)
);

INVxp67_ASAP7_75t_SL g2400 ( 
.A(n_1983),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1632),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1633),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_1581),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_1588),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1634),
.Y(n_2405)
);

CKINVDCx16_ASAP7_75t_R g2406 ( 
.A(n_1587),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_1635),
.Y(n_2407)
);

CKINVDCx20_ASAP7_75t_R g2408 ( 
.A(n_1539),
.Y(n_2408)
);

BUFx3_ASAP7_75t_L g2409 ( 
.A(n_1530),
.Y(n_2409)
);

INVxp67_ASAP7_75t_SL g2410 ( 
.A(n_1958),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1637),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_1588),
.Y(n_2412)
);

CKINVDCx20_ASAP7_75t_R g2413 ( 
.A(n_1539),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1595),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_1596),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2034),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2011),
.Y(n_2417)
);

OA21x2_ASAP7_75t_L g2418 ( 
.A1(n_2109),
.A2(n_1786),
.B(n_1782),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2033),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2034),
.Y(n_2420)
);

BUFx6f_ASAP7_75t_L g2421 ( 
.A(n_2182),
.Y(n_2421)
);

INVx6_ASAP7_75t_L g2422 ( 
.A(n_2182),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2112),
.B(n_1496),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_2317),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2012),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2035),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_2317),
.Y(n_2427)
);

BUFx6f_ASAP7_75t_L g2428 ( 
.A(n_2146),
.Y(n_2428)
);

INVxp33_ASAP7_75t_SL g2429 ( 
.A(n_2393),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2020),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2307),
.B(n_1511),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2015),
.Y(n_2432)
);

INVx6_ASAP7_75t_L g2433 ( 
.A(n_2409),
.Y(n_2433)
);

BUFx8_ASAP7_75t_L g2434 ( 
.A(n_2050),
.Y(n_2434)
);

BUFx2_ASAP7_75t_L g2435 ( 
.A(n_2049),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2035),
.Y(n_2436)
);

AND2x4_ASAP7_75t_L g2437 ( 
.A(n_2113),
.B(n_2410),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2016),
.Y(n_2438)
);

BUFx6f_ASAP7_75t_L g2439 ( 
.A(n_2146),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2042),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2159),
.B(n_1511),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2017),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2042),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2018),
.Y(n_2444)
);

OA21x2_ASAP7_75t_L g2445 ( 
.A1(n_2309),
.A2(n_1786),
.B(n_1782),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_2370),
.B(n_1496),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2062),
.Y(n_2447)
);

BUFx6f_ASAP7_75t_L g2448 ( 
.A(n_2146),
.Y(n_2448)
);

OAI21x1_ASAP7_75t_L g2449 ( 
.A1(n_2310),
.A2(n_1809),
.B(n_1808),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2019),
.Y(n_2450)
);

OAI22xp5_ASAP7_75t_SL g2451 ( 
.A1(n_2342),
.A2(n_1312),
.B1(n_1361),
.B2(n_1296),
.Y(n_2451)
);

BUFx6f_ASAP7_75t_L g2452 ( 
.A(n_2146),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2267),
.Y(n_2453)
);

OAI22xp5_ASAP7_75t_SL g2454 ( 
.A1(n_2342),
.A2(n_1312),
.B1(n_1361),
.B2(n_1296),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2371),
.B(n_1985),
.Y(n_2455)
);

BUFx2_ASAP7_75t_L g2456 ( 
.A(n_2054),
.Y(n_2456)
);

OAI22xp5_ASAP7_75t_L g2457 ( 
.A1(n_2333),
.A2(n_1707),
.B1(n_1715),
.B2(n_1563),
.Y(n_2457)
);

AOI22xp5_ASAP7_75t_L g2458 ( 
.A1(n_2147),
.A2(n_1707),
.B1(n_1694),
.B2(n_1540),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2062),
.Y(n_2459)
);

AND2x4_ASAP7_75t_L g2460 ( 
.A(n_2372),
.B(n_1563),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2068),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2068),
.Y(n_2462)
);

INVx4_ASAP7_75t_L g2463 ( 
.A(n_2159),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2022),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2091),
.Y(n_2465)
);

HB1xp67_ASAP7_75t_L g2466 ( 
.A(n_2082),
.Y(n_2466)
);

INVx3_ASAP7_75t_L g2467 ( 
.A(n_2267),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2024),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2091),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2061),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2140),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2140),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2159),
.B(n_1537),
.Y(n_2473)
);

BUFx3_ASAP7_75t_L g2474 ( 
.A(n_2409),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2026),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2378),
.B(n_1715),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2021),
.B(n_2023),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2336),
.A2(n_1540),
.B1(n_1799),
.B2(n_1747),
.Y(n_2478)
);

INVx2_ASAP7_75t_L g2479 ( 
.A(n_2150),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_2267),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_SL g2481 ( 
.A1(n_2344),
.A2(n_1420),
.B1(n_1430),
.B2(n_1411),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2371),
.B(n_1596),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2150),
.Y(n_2483)
);

AND2x6_ASAP7_75t_L g2484 ( 
.A(n_2002),
.B(n_1277),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2225),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2225),
.Y(n_2486)
);

INVxp67_ASAP7_75t_L g2487 ( 
.A(n_2098),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2235),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2029),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2036),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2038),
.Y(n_2491)
);

INVx4_ASAP7_75t_L g2492 ( 
.A(n_2394),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2040),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2056),
.B(n_1544),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2043),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2057),
.B(n_1550),
.Y(n_2496)
);

BUFx3_ASAP7_75t_L g2497 ( 
.A(n_2117),
.Y(n_2497)
);

AND2x6_ASAP7_75t_L g2498 ( 
.A(n_2004),
.B(n_1299),
.Y(n_2498)
);

INVx3_ASAP7_75t_L g2499 ( 
.A(n_2394),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_2118),
.Y(n_2500)
);

CKINVDCx20_ASAP7_75t_R g2501 ( 
.A(n_2007),
.Y(n_2501)
);

OAI22xp5_ASAP7_75t_SL g2502 ( 
.A1(n_2344),
.A2(n_1420),
.B1(n_1430),
.B2(n_1411),
.Y(n_2502)
);

BUFx2_ASAP7_75t_L g2503 ( 
.A(n_2107),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2046),
.Y(n_2504)
);

INVx3_ASAP7_75t_L g2505 ( 
.A(n_2394),
.Y(n_2505)
);

HB1xp67_ASAP7_75t_L g2506 ( 
.A(n_2133),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2394),
.Y(n_2507)
);

INVxp33_ASAP7_75t_SL g2508 ( 
.A(n_2393),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2375),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2072),
.B(n_1597),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2047),
.Y(n_2511)
);

OAI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2338),
.A2(n_1813),
.B1(n_1470),
.B2(n_1576),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2235),
.Y(n_2513)
);

AND2x4_ASAP7_75t_L g2514 ( 
.A(n_2071),
.B(n_1938),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_2248),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2006),
.B(n_1597),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2354),
.Y(n_2517)
);

INVx4_ASAP7_75t_L g2518 ( 
.A(n_2394),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2061),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2248),
.Y(n_2520)
);

AOI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_2213),
.A2(n_2346),
.B1(n_2367),
.B2(n_2269),
.Y(n_2521)
);

BUFx3_ASAP7_75t_L g2522 ( 
.A(n_2121),
.Y(n_2522)
);

CKINVDCx16_ASAP7_75t_R g2523 ( 
.A(n_2028),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2243),
.B(n_2275),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2298),
.Y(n_2525)
);

AND2x4_ASAP7_75t_L g2526 ( 
.A(n_2073),
.B(n_1938),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2298),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2318),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2093),
.Y(n_2529)
);

AOI22xp5_ASAP7_75t_L g2530 ( 
.A1(n_2241),
.A2(n_1605),
.B1(n_1613),
.B2(n_1603),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2051),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_SL g2532 ( 
.A(n_2106),
.B(n_1967),
.Y(n_2532)
);

INVx2_ASAP7_75t_SL g2533 ( 
.A(n_2177),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2394),
.Y(n_2534)
);

BUFx2_ASAP7_75t_L g2535 ( 
.A(n_2274),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2053),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2059),
.Y(n_2537)
);

OAI22xp5_ASAP7_75t_SL g2538 ( 
.A1(n_2332),
.A2(n_1453),
.B1(n_1065),
.B2(n_1101),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2074),
.B(n_1603),
.Y(n_2539)
);

HB1xp67_ASAP7_75t_L g2540 ( 
.A(n_2406),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2008),
.B(n_1605),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2318),
.Y(n_2542)
);

BUFx3_ASAP7_75t_L g2543 ( 
.A(n_2128),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2324),
.Y(n_2544)
);

BUFx6f_ASAP7_75t_L g2545 ( 
.A(n_2324),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2079),
.B(n_2087),
.Y(n_2546)
);

HB1xp67_ASAP7_75t_L g2547 ( 
.A(n_2322),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2060),
.Y(n_2548)
);

BUFx2_ASAP7_75t_L g2549 ( 
.A(n_2335),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2349),
.Y(n_2550)
);

BUFx3_ASAP7_75t_L g2551 ( 
.A(n_2138),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2349),
.Y(n_2552)
);

HB1xp67_ASAP7_75t_L g2553 ( 
.A(n_2352),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2063),
.Y(n_2554)
);

BUFx6f_ASAP7_75t_L g2555 ( 
.A(n_2351),
.Y(n_2555)
);

AOI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2243),
.A2(n_1616),
.B1(n_1617),
.B2(n_1613),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2067),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2096),
.B(n_2114),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2005),
.Y(n_2559)
);

BUFx3_ASAP7_75t_L g2560 ( 
.A(n_2142),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2110),
.B(n_1978),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2130),
.B(n_1616),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2143),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2144),
.Y(n_2564)
);

INVx2_ASAP7_75t_L g2565 ( 
.A(n_2351),
.Y(n_2565)
);

CKINVDCx8_ASAP7_75t_R g2566 ( 
.A(n_2124),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2149),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2010),
.B(n_1617),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2151),
.Y(n_2569)
);

BUFx6f_ASAP7_75t_L g2570 ( 
.A(n_2379),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2381),
.Y(n_2571)
);

BUFx6f_ASAP7_75t_L g2572 ( 
.A(n_2383),
.Y(n_2572)
);

AND2x6_ASAP7_75t_L g2573 ( 
.A(n_2013),
.B(n_1299),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2368),
.Y(n_2574)
);

BUFx6f_ASAP7_75t_L g2575 ( 
.A(n_2385),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2368),
.Y(n_2576)
);

AND2x2_ASAP7_75t_SL g2577 ( 
.A(n_2009),
.B(n_858),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2153),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2377),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2377),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2154),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2156),
.Y(n_2582)
);

BUFx6f_ASAP7_75t_L g2583 ( 
.A(n_2386),
.Y(n_2583)
);

INVx6_ASAP7_75t_L g2584 ( 
.A(n_2131),
.Y(n_2584)
);

INVx3_ASAP7_75t_L g2585 ( 
.A(n_2403),
.Y(n_2585)
);

NOR2x1_ASAP7_75t_L g2586 ( 
.A(n_2160),
.B(n_1658),
.Y(n_2586)
);

INVxp67_ASAP7_75t_L g2587 ( 
.A(n_2088),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2403),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2414),
.Y(n_2589)
);

INVx6_ASAP7_75t_L g2590 ( 
.A(n_2132),
.Y(n_2590)
);

OAI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2239),
.A2(n_1541),
.B1(n_1661),
.B2(n_1143),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2414),
.Y(n_2592)
);

AND2x2_ASAP7_75t_SL g2593 ( 
.A(n_2039),
.B(n_858),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2162),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2311),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2312),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2134),
.B(n_1621),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2168),
.B(n_2169),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2139),
.B(n_1621),
.Y(n_2599)
);

INVx3_ASAP7_75t_L g2600 ( 
.A(n_2313),
.Y(n_2600)
);

BUFx6f_ASAP7_75t_L g2601 ( 
.A(n_2389),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_SL g2602 ( 
.A1(n_2359),
.A2(n_1065),
.B1(n_1101),
.B2(n_1059),
.Y(n_2602)
);

NAND3xp33_ASAP7_75t_L g2603 ( 
.A(n_2115),
.B(n_1641),
.C(n_1629),
.Y(n_2603)
);

AND2x6_ASAP7_75t_L g2604 ( 
.A(n_2075),
.B(n_1303),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2170),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2178),
.B(n_1629),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2171),
.Y(n_2607)
);

OAI22xp5_ASAP7_75t_SL g2608 ( 
.A1(n_2332),
.A2(n_1453),
.B1(n_1112),
.B2(n_1161),
.Y(n_2608)
);

BUFx3_ASAP7_75t_L g2609 ( 
.A(n_2076),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2316),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2183),
.B(n_1641),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2077),
.B(n_1660),
.Y(n_2612)
);

INVx2_ASAP7_75t_SL g2613 ( 
.A(n_2120),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2319),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2172),
.Y(n_2615)
);

INVx3_ASAP7_75t_L g2616 ( 
.A(n_2321),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2173),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2174),
.Y(n_2618)
);

AOI22x1_ASAP7_75t_SL g2619 ( 
.A1(n_2297),
.A2(n_1112),
.B1(n_1161),
.B2(n_1059),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_2204),
.B(n_1644),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2325),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2176),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2330),
.Y(n_2623)
);

AND2x6_ASAP7_75t_L g2624 ( 
.A(n_2078),
.B(n_1303),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2331),
.Y(n_2625)
);

AND2x4_ASAP7_75t_L g2626 ( 
.A(n_2081),
.B(n_1942),
.Y(n_2626)
);

AND2x4_ASAP7_75t_L g2627 ( 
.A(n_2083),
.B(n_2000),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2390),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2334),
.Y(n_2629)
);

AND2x6_ASAP7_75t_L g2630 ( 
.A(n_2084),
.B(n_1308),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2339),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2348),
.Y(n_2632)
);

XNOR2x2_ASAP7_75t_R g2633 ( 
.A(n_2007),
.B(n_1710),
.Y(n_2633)
);

BUFx6f_ASAP7_75t_L g2634 ( 
.A(n_2391),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2179),
.B(n_1644),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_2355),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2220),
.B(n_1659),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2356),
.Y(n_2638)
);

BUFx6f_ASAP7_75t_L g2639 ( 
.A(n_2357),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2085),
.B(n_921),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2086),
.B(n_1308),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2181),
.B(n_1659),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2186),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_SL g2644 ( 
.A1(n_2337),
.A2(n_1351),
.B1(n_1407),
.B2(n_1306),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2187),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2358),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2362),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_2404),
.Y(n_2648)
);

AND2x4_ASAP7_75t_L g2649 ( 
.A(n_2089),
.B(n_1310),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2188),
.Y(n_2650)
);

INVx3_ASAP7_75t_L g2651 ( 
.A(n_2363),
.Y(n_2651)
);

OA21x2_ASAP7_75t_L g2652 ( 
.A1(n_2365),
.A2(n_1809),
.B(n_1808),
.Y(n_2652)
);

INVx3_ASAP7_75t_L g2653 ( 
.A(n_2369),
.Y(n_2653)
);

OAI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2239),
.A2(n_1143),
.B1(n_869),
.B2(n_875),
.Y(n_2654)
);

CKINVDCx20_ASAP7_75t_R g2655 ( 
.A(n_2031),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2373),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2275),
.B(n_1664),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2404),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2374),
.Y(n_2659)
);

BUFx6f_ASAP7_75t_L g2660 ( 
.A(n_2392),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2189),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2396),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2190),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2397),
.Y(n_2664)
);

BUFx6f_ASAP7_75t_L g2665 ( 
.A(n_2398),
.Y(n_2665)
);

INVx5_ASAP7_75t_L g2666 ( 
.A(n_2273),
.Y(n_2666)
);

BUFx6f_ASAP7_75t_L g2667 ( 
.A(n_2401),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_2402),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2192),
.B(n_1664),
.Y(n_2669)
);

XOR2xp5_ASAP7_75t_L g2670 ( 
.A(n_2297),
.B(n_1306),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2194),
.B(n_1666),
.Y(n_2671)
);

INVx3_ASAP7_75t_L g2672 ( 
.A(n_2405),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_2407),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2288),
.B(n_2292),
.Y(n_2674)
);

INVx3_ASAP7_75t_L g2675 ( 
.A(n_2411),
.Y(n_2675)
);

AOI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2127),
.A2(n_1667),
.B1(n_1668),
.B2(n_1666),
.Y(n_2676)
);

OAI22x1_ASAP7_75t_L g2677 ( 
.A1(n_2412),
.A2(n_1650),
.B1(n_1599),
.B2(n_1272),
.Y(n_2677)
);

INVx6_ASAP7_75t_L g2678 ( 
.A(n_2295),
.Y(n_2678)
);

BUFx12f_ASAP7_75t_L g2679 ( 
.A(n_2025),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2196),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2314),
.B(n_1667),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2197),
.Y(n_2682)
);

BUFx12f_ASAP7_75t_L g2683 ( 
.A(n_2027),
.Y(n_2683)
);

BUFx3_ASAP7_75t_L g2684 ( 
.A(n_2090),
.Y(n_2684)
);

OA21x2_ASAP7_75t_L g2685 ( 
.A1(n_2387),
.A2(n_1820),
.B(n_1815),
.Y(n_2685)
);

AND2x4_ASAP7_75t_L g2686 ( 
.A(n_2092),
.B(n_1310),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2094),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2097),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2199),
.Y(n_2689)
);

BUFx6f_ASAP7_75t_L g2690 ( 
.A(n_2100),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2101),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2327),
.B(n_1668),
.Y(n_2692)
);

CKINVDCx8_ASAP7_75t_R g2693 ( 
.A(n_2222),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2103),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2200),
.Y(n_2695)
);

AOI22xp5_ASAP7_75t_L g2696 ( 
.A1(n_2127),
.A2(n_1672),
.B1(n_1681),
.B2(n_1669),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2125),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2104),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2108),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2201),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2350),
.B(n_1669),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2412),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_SL g2703 ( 
.A(n_2255),
.B(n_1672),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2202),
.Y(n_2704)
);

INVx6_ASAP7_75t_L g2705 ( 
.A(n_2400),
.Y(n_2705)
);

OAI21x1_ASAP7_75t_L g2706 ( 
.A1(n_2203),
.A2(n_1820),
.B(n_1815),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2205),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2207),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2184),
.B(n_1681),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2184),
.B(n_1698),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2209),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2210),
.B(n_2211),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2212),
.B(n_1698),
.Y(n_2713)
);

CKINVDCx20_ASAP7_75t_R g2714 ( 
.A(n_2031),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2214),
.B(n_1702),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_SL g2716 ( 
.A(n_2126),
.B(n_1955),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2215),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2216),
.Y(n_2718)
);

BUFx8_ASAP7_75t_L g2719 ( 
.A(n_2341),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2217),
.B(n_1702),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2218),
.Y(n_2721)
);

BUFx6f_ASAP7_75t_L g2722 ( 
.A(n_2219),
.Y(n_2722)
);

OA21x2_ASAP7_75t_L g2723 ( 
.A1(n_2221),
.A2(n_1829),
.B(n_1823),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2224),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2226),
.B(n_1705),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_2227),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2228),
.B(n_1705),
.Y(n_2727)
);

OAI22xp5_ASAP7_75t_SL g2728 ( 
.A1(n_2337),
.A2(n_1407),
.B1(n_1418),
.B2(n_1351),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_2229),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2032),
.B(n_1709),
.Y(n_2730)
);

NAND2xp5_ASAP7_75t_L g2731 ( 
.A(n_2230),
.B(n_2231),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2232),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2233),
.B(n_1709),
.Y(n_2733)
);

INVx4_ASAP7_75t_L g2734 ( 
.A(n_2234),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2240),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2244),
.B(n_1712),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2245),
.Y(n_2737)
);

OAI22xp5_ASAP7_75t_SL g2738 ( 
.A1(n_2044),
.A2(n_1427),
.B1(n_1468),
.B2(n_1418),
.Y(n_2738)
);

CKINVDCx6p67_ASAP7_75t_R g2739 ( 
.A(n_2111),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2246),
.B(n_1712),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2253),
.B(n_1319),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2254),
.Y(n_2742)
);

BUFx6f_ASAP7_75t_L g2743 ( 
.A(n_2256),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2259),
.B(n_1716),
.Y(n_2744)
);

INVx4_ASAP7_75t_L g2745 ( 
.A(n_2261),
.Y(n_2745)
);

AOI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2320),
.A2(n_1719),
.B1(n_1722),
.B2(n_1716),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2263),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2266),
.Y(n_2748)
);

BUFx3_ASAP7_75t_L g2749 ( 
.A(n_2270),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2272),
.Y(n_2750)
);

HB1xp67_ASAP7_75t_L g2751 ( 
.A(n_2388),
.Y(n_2751)
);

AOI22xp5_ASAP7_75t_L g2752 ( 
.A1(n_2320),
.A2(n_1722),
.B1(n_1735),
.B2(n_1719),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2276),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2415),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2277),
.B(n_1735),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2278),
.B(n_2282),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2283),
.Y(n_2757)
);

BUFx12f_ASAP7_75t_L g2758 ( 
.A(n_2030),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2285),
.Y(n_2759)
);

HB1xp67_ASAP7_75t_L g2760 ( 
.A(n_2399),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2286),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2287),
.B(n_2289),
.Y(n_2762)
);

BUFx3_ASAP7_75t_L g2763 ( 
.A(n_2290),
.Y(n_2763)
);

BUFx8_ASAP7_75t_L g2764 ( 
.A(n_2123),
.Y(n_2764)
);

INVx5_ASAP7_75t_L g2765 ( 
.A(n_2145),
.Y(n_2765)
);

OAI21x1_ASAP7_75t_L g2766 ( 
.A1(n_2291),
.A2(n_1829),
.B(n_1823),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2293),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2294),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2296),
.Y(n_2769)
);

BUFx2_ASAP7_75t_L g2770 ( 
.A(n_2359),
.Y(n_2770)
);

AND2x2_ASAP7_75t_SL g2771 ( 
.A(n_2157),
.B(n_859),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2299),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2300),
.Y(n_2773)
);

BUFx6f_ASAP7_75t_L g2774 ( 
.A(n_2302),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2303),
.Y(n_2775)
);

OAI22xp5_ASAP7_75t_SL g2776 ( 
.A1(n_2044),
.A2(n_1427),
.B1(n_1209),
.B2(n_1068),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_2304),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2305),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2032),
.B(n_1742),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2129),
.Y(n_2780)
);

CKINVDCx5p33_ASAP7_75t_R g2781 ( 
.A(n_2135),
.Y(n_2781)
);

BUFx8_ASAP7_75t_L g2782 ( 
.A(n_2166),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2137),
.Y(n_2783)
);

BUFx6f_ASAP7_75t_L g2784 ( 
.A(n_2323),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2155),
.Y(n_2785)
);

NOR2xp33_ASAP7_75t_L g2786 ( 
.A(n_2065),
.B(n_1742),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2262),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2281),
.Y(n_2788)
);

INVx3_ASAP7_75t_L g2789 ( 
.A(n_2323),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2326),
.A2(n_874),
.B1(n_902),
.B2(n_878),
.Y(n_2790)
);

BUFx2_ASAP7_75t_L g2791 ( 
.A(n_2360),
.Y(n_2791)
);

OA21x2_ASAP7_75t_L g2792 ( 
.A1(n_2326),
.A2(n_1866),
.B(n_1849),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2158),
.Y(n_2793)
);

BUFx8_ASAP7_75t_L g2794 ( 
.A(n_2264),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2366),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2164),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2376),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2382),
.Y(n_2798)
);

INVx3_ASAP7_75t_L g2799 ( 
.A(n_2329),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2165),
.Y(n_2800)
);

BUFx6f_ASAP7_75t_L g2801 ( 
.A(n_2175),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2329),
.B(n_1319),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2193),
.B(n_1743),
.Y(n_2803)
);

OAI22xp5_ASAP7_75t_SL g2804 ( 
.A1(n_2048),
.A2(n_1021),
.B1(n_1038),
.B2(n_1020),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2206),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_2208),
.Y(n_2806)
);

BUFx12f_ASAP7_75t_L g2807 ( 
.A(n_2037),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2223),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2242),
.Y(n_2809)
);

BUFx6f_ASAP7_75t_L g2810 ( 
.A(n_2247),
.Y(n_2810)
);

OAI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2340),
.A2(n_908),
.B1(n_918),
.B2(n_911),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2249),
.Y(n_2812)
);

NOR2xp33_ASAP7_75t_L g2813 ( 
.A(n_2065),
.B(n_1743),
.Y(n_2813)
);

AND2x6_ASAP7_75t_L g2814 ( 
.A(n_2237),
.B(n_1352),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_L g2815 ( 
.A(n_2080),
.B(n_1746),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2250),
.Y(n_2816)
);

BUFx12f_ASAP7_75t_L g2817 ( 
.A(n_2041),
.Y(n_2817)
);

INVx3_ASAP7_75t_L g2818 ( 
.A(n_2340),
.Y(n_2818)
);

AND2x4_ASAP7_75t_L g2819 ( 
.A(n_2343),
.B(n_1352),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2080),
.B(n_1746),
.Y(n_2820)
);

AND2x2_ASAP7_75t_SL g2821 ( 
.A(n_2280),
.B(n_859),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2343),
.B(n_1754),
.Y(n_2822)
);

OA21x2_ASAP7_75t_L g2823 ( 
.A1(n_2345),
.A2(n_1866),
.B(n_1849),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2257),
.Y(n_2824)
);

BUFx8_ASAP7_75t_L g2825 ( 
.A(n_2003),
.Y(n_2825)
);

INVxp67_ASAP7_75t_L g2826 ( 
.A(n_2279),
.Y(n_2826)
);

HB1xp67_ASAP7_75t_L g2827 ( 
.A(n_2284),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2301),
.Y(n_2828)
);

INVx3_ASAP7_75t_L g2829 ( 
.A(n_2345),
.Y(n_2829)
);

BUFx3_ASAP7_75t_L g2830 ( 
.A(n_2308),
.Y(n_2830)
);

BUFx6f_ASAP7_75t_L g2831 ( 
.A(n_2347),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2347),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2353),
.B(n_1754),
.Y(n_2833)
);

AND2x6_ASAP7_75t_L g2834 ( 
.A(n_2353),
.B(n_1358),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2380),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2380),
.Y(n_2836)
);

CKINVDCx6p67_ASAP7_75t_R g2837 ( 
.A(n_2306),
.Y(n_2837)
);

INVx5_ASAP7_75t_L g2838 ( 
.A(n_2384),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2384),
.B(n_1757),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_2045),
.Y(n_2840)
);

BUFx6f_ASAP7_75t_L g2841 ( 
.A(n_2055),
.Y(n_2841)
);

OAI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2003),
.A2(n_927),
.B1(n_941),
.B2(n_928),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2001),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2001),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2095),
.B(n_1757),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2095),
.A2(n_1761),
.B1(n_1765),
.B2(n_1758),
.Y(n_2846)
);

INVx6_ASAP7_75t_L g2847 ( 
.A(n_2102),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2014),
.Y(n_2848)
);

BUFx3_ASAP7_75t_L g2849 ( 
.A(n_2014),
.Y(n_2849)
);

BUFx6f_ASAP7_75t_L g2850 ( 
.A(n_2058),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2058),
.Y(n_2851)
);

CKINVDCx16_ASAP7_75t_R g2852 ( 
.A(n_2306),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2102),
.B(n_1758),
.Y(n_2853)
);

CKINVDCx5p33_ASAP7_75t_R g2854 ( 
.A(n_2069),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_L g2855 ( 
.A(n_2069),
.Y(n_2855)
);

BUFx2_ASAP7_75t_L g2856 ( 
.A(n_2360),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2361),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2136),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2136),
.Y(n_2859)
);

CKINVDCx6p67_ASAP7_75t_R g2860 ( 
.A(n_2315),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2361),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2364),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2364),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2315),
.B(n_1761),
.Y(n_2864)
);

OAI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2395),
.A2(n_949),
.B1(n_951),
.B2(n_950),
.Y(n_2865)
);

CKINVDCx20_ASAP7_75t_R g2866 ( 
.A(n_2048),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2395),
.Y(n_2867)
);

INVx3_ASAP7_75t_L g2868 ( 
.A(n_2070),
.Y(n_2868)
);

BUFx3_ASAP7_75t_L g2869 ( 
.A(n_2328),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2408),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2408),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2413),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2413),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2328),
.B(n_1765),
.Y(n_2874)
);

AND2x6_ASAP7_75t_L g2875 ( 
.A(n_2070),
.B(n_1358),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2052),
.Y(n_2876)
);

INVx5_ASAP7_75t_L g2877 ( 
.A(n_2052),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2064),
.Y(n_2878)
);

CKINVDCx5p33_ASAP7_75t_R g2879 ( 
.A(n_2064),
.Y(n_2879)
);

BUFx3_ASAP7_75t_L g2880 ( 
.A(n_2066),
.Y(n_2880)
);

AND2x4_ASAP7_75t_L g2881 ( 
.A(n_2066),
.B(n_1371),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2271),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_2421),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2416),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2416),
.Y(n_2885)
);

HB1xp67_ASAP7_75t_L g2886 ( 
.A(n_2455),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2455),
.B(n_1804),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2420),
.Y(n_2888)
);

INVx2_ASAP7_75t_L g2889 ( 
.A(n_2420),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2426),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2426),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2436),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2436),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2437),
.B(n_1768),
.Y(n_2894)
);

AND2x6_ASAP7_75t_L g2895 ( 
.A(n_2499),
.B(n_859),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2440),
.Y(n_2896)
);

CKINVDCx8_ASAP7_75t_R g2897 ( 
.A(n_2523),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2598),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2598),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2756),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2440),
.Y(n_2901)
);

OA21x2_ASAP7_75t_L g2902 ( 
.A1(n_2706),
.A2(n_1879),
.B(n_1871),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_2754),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_SL g2904 ( 
.A(n_2838),
.B(n_1768),
.Y(n_2904)
);

NOR2xp33_ASAP7_75t_L g2905 ( 
.A(n_2435),
.B(n_1771),
.Y(n_2905)
);

BUFx6f_ASAP7_75t_L g2906 ( 
.A(n_2421),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2756),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2443),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2437),
.B(n_2417),
.Y(n_2909)
);

AND2x2_ASAP7_75t_L g2910 ( 
.A(n_2435),
.B(n_2456),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2443),
.Y(n_2911)
);

AND2x4_ASAP7_75t_L g2912 ( 
.A(n_2765),
.B(n_870),
.Y(n_2912)
);

BUFx6f_ASAP7_75t_L g2913 ( 
.A(n_2421),
.Y(n_2913)
);

BUFx6f_ASAP7_75t_L g2914 ( 
.A(n_2421),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2762),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2762),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2447),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2447),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2687),
.Y(n_2919)
);

CKINVDCx5p33_ASAP7_75t_R g2920 ( 
.A(n_2754),
.Y(n_2920)
);

HB1xp67_ASAP7_75t_L g2921 ( 
.A(n_2503),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2459),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2459),
.Y(n_2923)
);

BUFx6f_ASAP7_75t_L g2924 ( 
.A(n_2424),
.Y(n_2924)
);

HB1xp67_ASAP7_75t_L g2925 ( 
.A(n_2503),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2461),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2838),
.B(n_1819),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2461),
.Y(n_2928)
);

INVx2_ASAP7_75t_L g2929 ( 
.A(n_2462),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2462),
.Y(n_2930)
);

CKINVDCx5p33_ASAP7_75t_R g2931 ( 
.A(n_2781),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_SL g2932 ( 
.A(n_2838),
.B(n_1819),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2465),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2465),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2437),
.B(n_1771),
.Y(n_2935)
);

CKINVDCx5p33_ASAP7_75t_R g2936 ( 
.A(n_2781),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2469),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2425),
.B(n_1777),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2687),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2688),
.Y(n_2940)
);

INVx3_ASAP7_75t_L g2941 ( 
.A(n_2499),
.Y(n_2941)
);

BUFx2_ASAP7_75t_L g2942 ( 
.A(n_2517),
.Y(n_2942)
);

BUFx6f_ASAP7_75t_L g2943 ( 
.A(n_2424),
.Y(n_2943)
);

INVx4_ASAP7_75t_L g2944 ( 
.A(n_2584),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2430),
.B(n_1777),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2688),
.Y(n_2946)
);

HB1xp67_ASAP7_75t_L g2947 ( 
.A(n_2456),
.Y(n_2947)
);

OA21x2_ASAP7_75t_L g2948 ( 
.A1(n_2706),
.A2(n_1879),
.B(n_1871),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2469),
.Y(n_2949)
);

BUFx8_ASAP7_75t_L g2950 ( 
.A(n_2517),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2471),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2471),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2472),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2717),
.B(n_1789),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2472),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2691),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2765),
.B(n_872),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2691),
.Y(n_2958)
);

AND2x6_ASAP7_75t_L g2959 ( 
.A(n_2499),
.B(n_871),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2479),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2479),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2694),
.Y(n_2962)
);

INVx3_ASAP7_75t_L g2963 ( 
.A(n_2505),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2424),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2483),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2717),
.B(n_1789),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2483),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2485),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2485),
.Y(n_2969)
);

BUFx6f_ASAP7_75t_L g2970 ( 
.A(n_2424),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_SL g2971 ( 
.A(n_2838),
.B(n_1795),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2486),
.Y(n_2972)
);

BUFx6f_ASAP7_75t_L g2973 ( 
.A(n_2639),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2486),
.Y(n_2974)
);

INVx2_ASAP7_75t_L g2975 ( 
.A(n_2488),
.Y(n_2975)
);

NOR2xp33_ASAP7_75t_L g2976 ( 
.A(n_2500),
.B(n_1790),
.Y(n_2976)
);

BUFx6f_ASAP7_75t_L g2977 ( 
.A(n_2639),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2488),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2513),
.Y(n_2979)
);

NAND3xp33_ASAP7_75t_L g2980 ( 
.A(n_2709),
.B(n_1795),
.C(n_1790),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2513),
.Y(n_2981)
);

AND2x4_ASAP7_75t_L g2982 ( 
.A(n_2765),
.B(n_872),
.Y(n_2982)
);

BUFx8_ASAP7_75t_L g2983 ( 
.A(n_2770),
.Y(n_2983)
);

AND2x2_ASAP7_75t_SL g2984 ( 
.A(n_2577),
.B(n_871),
.Y(n_2984)
);

AND2x6_ASAP7_75t_L g2985 ( 
.A(n_2505),
.B(n_871),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2525),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2525),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2717),
.B(n_1798),
.Y(n_2988)
);

INVx3_ASAP7_75t_L g2989 ( 
.A(n_2505),
.Y(n_2989)
);

INVxp67_ASAP7_75t_L g2990 ( 
.A(n_2500),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2527),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2527),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2542),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2542),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2552),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2552),
.Y(n_2996)
);

NAND2xp33_ASAP7_75t_SL g2997 ( 
.A(n_2831),
.B(n_1142),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_2565),
.Y(n_2998)
);

AND2x4_ASAP7_75t_L g2999 ( 
.A(n_2765),
.B(n_880),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2565),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2574),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_SL g3002 ( 
.A(n_2838),
.B(n_1824),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2574),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_SL g3004 ( 
.A(n_2831),
.B(n_1824),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2576),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2576),
.Y(n_3006)
);

INVx2_ASAP7_75t_L g3007 ( 
.A(n_2579),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2579),
.Y(n_3008)
);

BUFx2_ASAP7_75t_L g3009 ( 
.A(n_2540),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2446),
.B(n_1798),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2580),
.Y(n_3011)
);

OA21x2_ASAP7_75t_L g3012 ( 
.A1(n_2766),
.A2(n_1890),
.B(n_1887),
.Y(n_3012)
);

INVxp67_ASAP7_75t_L g3013 ( 
.A(n_2466),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2580),
.Y(n_3014)
);

BUFx12f_ASAP7_75t_L g3015 ( 
.A(n_2764),
.Y(n_3015)
);

BUFx6f_ASAP7_75t_L g3016 ( 
.A(n_2639),
.Y(n_3016)
);

BUFx6f_ASAP7_75t_L g3017 ( 
.A(n_2639),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2588),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2446),
.B(n_1804),
.Y(n_3019)
);

INVx3_ASAP7_75t_L g3020 ( 
.A(n_2507),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2588),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2589),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2589),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2446),
.B(n_1805),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2592),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2460),
.B(n_1805),
.Y(n_3026)
);

HB1xp67_ASAP7_75t_L g3027 ( 
.A(n_2535),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2592),
.Y(n_3028)
);

AND2x6_ASAP7_75t_L g3029 ( 
.A(n_2507),
.B(n_915),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_SL g3030 ( 
.A(n_2419),
.B(n_1206),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2449),
.Y(n_3031)
);

NOR2xp33_ASAP7_75t_L g3032 ( 
.A(n_2710),
.B(n_1811),
.Y(n_3032)
);

NOR2xp33_ASAP7_75t_L g3033 ( 
.A(n_2487),
.B(n_1811),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_2449),
.Y(n_3034)
);

BUFx6f_ASAP7_75t_L g3035 ( 
.A(n_2639),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2766),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2550),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2460),
.B(n_1828),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2550),
.Y(n_3039)
);

AND2x4_ASAP7_75t_L g3040 ( 
.A(n_2765),
.B(n_880),
.Y(n_3040)
);

AOI22xp5_ASAP7_75t_L g3041 ( 
.A1(n_2834),
.A2(n_1837),
.B1(n_1842),
.B2(n_1828),
.Y(n_3041)
);

AND2x4_ASAP7_75t_L g3042 ( 
.A(n_2831),
.B(n_882),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2723),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2723),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2550),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2448),
.Y(n_3046)
);

AND2x4_ASAP7_75t_L g3047 ( 
.A(n_2831),
.B(n_882),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2723),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2445),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2423),
.B(n_2460),
.Y(n_3050)
);

INVx3_ASAP7_75t_L g3051 ( 
.A(n_2507),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2585),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2585),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2445),
.Y(n_3054)
);

BUFx6f_ASAP7_75t_L g3055 ( 
.A(n_2448),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2476),
.B(n_1837),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2445),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2694),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2652),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_L g3060 ( 
.A(n_2448),
.Y(n_3060)
);

AOI22xp5_ASAP7_75t_L g3061 ( 
.A1(n_2834),
.A2(n_1846),
.B1(n_1847),
.B2(n_1842),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2476),
.B(n_1846),
.Y(n_3062)
);

AND2x4_ASAP7_75t_L g3063 ( 
.A(n_2831),
.B(n_883),
.Y(n_3063)
);

AND2x2_ASAP7_75t_SL g3064 ( 
.A(n_2577),
.B(n_915),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2652),
.Y(n_3065)
);

HB1xp67_ASAP7_75t_L g3066 ( 
.A(n_2535),
.Y(n_3066)
);

HB1xp67_ASAP7_75t_L g3067 ( 
.A(n_2549),
.Y(n_3067)
);

INVx1_ASAP7_75t_L g3068 ( 
.A(n_2698),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2476),
.B(n_1847),
.Y(n_3069)
);

BUFx6f_ASAP7_75t_L g3070 ( 
.A(n_2448),
.Y(n_3070)
);

INVx3_ASAP7_75t_L g3071 ( 
.A(n_2534),
.Y(n_3071)
);

BUFx6f_ASAP7_75t_L g3072 ( 
.A(n_2448),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2652),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2783),
.B(n_1865),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2783),
.B(n_1865),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2698),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2699),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2699),
.Y(n_3078)
);

BUFx2_ASAP7_75t_SL g3079 ( 
.A(n_2492),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2700),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2834),
.B(n_1850),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2700),
.Y(n_3082)
);

INVx2_ASAP7_75t_L g3083 ( 
.A(n_2585),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2418),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_SL g3085 ( 
.A(n_2783),
.B(n_1867),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_L g3086 ( 
.A(n_2549),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2418),
.Y(n_3087)
);

AND2x2_ASAP7_75t_L g3088 ( 
.A(n_2423),
.B(n_1867),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2423),
.B(n_1868),
.Y(n_3089)
);

OA21x2_ASAP7_75t_L g3090 ( 
.A1(n_2596),
.A2(n_1890),
.B(n_1887),
.Y(n_3090)
);

AND2x4_ASAP7_75t_L g3091 ( 
.A(n_2812),
.B(n_883),
.Y(n_3091)
);

INVx5_ASAP7_75t_L g3092 ( 
.A(n_2492),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2704),
.Y(n_3093)
);

INVx2_ASAP7_75t_L g3094 ( 
.A(n_2418),
.Y(n_3094)
);

INVx1_ASAP7_75t_SL g3095 ( 
.A(n_2419),
.Y(n_3095)
);

INVx2_ASAP7_75t_L g3096 ( 
.A(n_2685),
.Y(n_3096)
);

HB1xp67_ASAP7_75t_L g3097 ( 
.A(n_2880),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2704),
.Y(n_3098)
);

AND2x4_ASAP7_75t_L g3099 ( 
.A(n_2812),
.B(n_891),
.Y(n_3099)
);

INVx3_ASAP7_75t_L g3100 ( 
.A(n_2534),
.Y(n_3100)
);

BUFx6f_ASAP7_75t_L g3101 ( 
.A(n_2452),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2707),
.Y(n_3102)
);

AND2x2_ASAP7_75t_L g3103 ( 
.A(n_2514),
.B(n_1869),
.Y(n_3103)
);

INVx2_ASAP7_75t_L g3104 ( 
.A(n_2685),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2685),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2707),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_SL g3107 ( 
.A(n_2783),
.B(n_1869),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2735),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2735),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2742),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2830),
.B(n_2783),
.Y(n_3111)
);

HB1xp67_ASAP7_75t_L g3112 ( 
.A(n_2880),
.Y(n_3112)
);

BUFx6f_ASAP7_75t_L g3113 ( 
.A(n_2452),
.Y(n_3113)
);

BUFx2_ASAP7_75t_L g3114 ( 
.A(n_2506),
.Y(n_3114)
);

BUFx6f_ASAP7_75t_L g3115 ( 
.A(n_2452),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2742),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2515),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2750),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2801),
.B(n_1877),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2515),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2515),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2515),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2750),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_2515),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_SL g3125 ( 
.A(n_2801),
.B(n_1877),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2753),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2596),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2514),
.B(n_1893),
.Y(n_3128)
);

BUFx6f_ASAP7_75t_L g3129 ( 
.A(n_2452),
.Y(n_3129)
);

OA21x2_ASAP7_75t_L g3130 ( 
.A1(n_2610),
.A2(n_2621),
.B(n_2614),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2801),
.B(n_1893),
.Y(n_3131)
);

OA21x2_ASAP7_75t_L g3132 ( 
.A1(n_2610),
.A2(n_1897),
.B(n_1711),
.Y(n_3132)
);

INVxp67_ASAP7_75t_L g3133 ( 
.A(n_2482),
.Y(n_3133)
);

AND2x2_ASAP7_75t_L g3134 ( 
.A(n_2514),
.B(n_1850),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2520),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2614),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_2621),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2623),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_2801),
.B(n_1854),
.Y(n_3139)
);

BUFx6f_ASAP7_75t_L g3140 ( 
.A(n_2452),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2623),
.Y(n_3141)
);

NOR2xp33_ASAP7_75t_SL g3142 ( 
.A(n_2470),
.B(n_1208),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2625),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2453),
.Y(n_3144)
);

AND2x4_ASAP7_75t_L g3145 ( 
.A(n_2830),
.B(n_891),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2526),
.B(n_1858),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2526),
.B(n_1858),
.Y(n_3147)
);

INVxp67_ASAP7_75t_L g3148 ( 
.A(n_2482),
.Y(n_3148)
);

INVx3_ASAP7_75t_L g3149 ( 
.A(n_2534),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2520),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2625),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2834),
.B(n_1854),
.Y(n_3152)
);

AND2x4_ASAP7_75t_L g3153 ( 
.A(n_2801),
.B(n_897),
.Y(n_3153)
);

CKINVDCx8_ASAP7_75t_R g3154 ( 
.A(n_2852),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2629),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2453),
.Y(n_3156)
);

XNOR2xp5_ASAP7_75t_SL g3157 ( 
.A(n_2670),
.B(n_2099),
.Y(n_3157)
);

BUFx2_ASAP7_75t_L g3158 ( 
.A(n_2882),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2520),
.Y(n_3159)
);

AND2x4_ASAP7_75t_L g3160 ( 
.A(n_2808),
.B(n_897),
.Y(n_3160)
);

INVx3_ASAP7_75t_L g3161 ( 
.A(n_2492),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2753),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2761),
.Y(n_3163)
);

HB1xp67_ASAP7_75t_L g3164 ( 
.A(n_2879),
.Y(n_3164)
);

OAI22xp5_ASAP7_75t_SL g3165 ( 
.A1(n_2602),
.A2(n_2105),
.B1(n_2116),
.B2(n_2099),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2520),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2520),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2761),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2432),
.Y(n_3169)
);

HB1xp67_ASAP7_75t_L g3170 ( 
.A(n_2879),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2438),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2528),
.Y(n_3172)
);

INVx2_ASAP7_75t_L g3173 ( 
.A(n_2528),
.Y(n_3173)
);

OR2x6_ASAP7_75t_L g3174 ( 
.A(n_2679),
.B(n_1371),
.Y(n_3174)
);

INVxp67_ASAP7_75t_L g3175 ( 
.A(n_2547),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2834),
.B(n_1855),
.Y(n_3176)
);

INVx3_ASAP7_75t_L g3177 ( 
.A(n_2518),
.Y(n_3177)
);

AND2x4_ASAP7_75t_L g3178 ( 
.A(n_2808),
.B(n_899),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2528),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2803),
.B(n_1855),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2442),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2444),
.Y(n_3182)
);

BUFx8_ASAP7_75t_L g3183 ( 
.A(n_2770),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2450),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2464),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2468),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2475),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2528),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2489),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_2526),
.B(n_1880),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2528),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2490),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2544),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2544),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2544),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2544),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2544),
.Y(n_3197)
);

BUFx6f_ASAP7_75t_L g3198 ( 
.A(n_2453),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2491),
.Y(n_3199)
);

CKINVDCx5p33_ASAP7_75t_R g3200 ( 
.A(n_2806),
.Y(n_3200)
);

INVx3_ASAP7_75t_L g3201 ( 
.A(n_2518),
.Y(n_3201)
);

AND2x2_ASAP7_75t_L g3202 ( 
.A(n_2820),
.B(n_1880),
.Y(n_3202)
);

BUFx6f_ASAP7_75t_L g3203 ( 
.A(n_2453),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2493),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_2545),
.Y(n_3205)
);

AND2x4_ASAP7_75t_L g3206 ( 
.A(n_2808),
.B(n_899),
.Y(n_3206)
);

INVx2_ASAP7_75t_L g3207 ( 
.A(n_2545),
.Y(n_3207)
);

INVx3_ASAP7_75t_L g3208 ( 
.A(n_2518),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2495),
.Y(n_3209)
);

OA21x2_ASAP7_75t_L g3210 ( 
.A1(n_2629),
.A2(n_1897),
.B(n_1714),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2545),
.Y(n_3211)
);

AND2x2_ASAP7_75t_L g3212 ( 
.A(n_2820),
.B(n_1886),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2504),
.Y(n_3213)
);

OA21x2_ASAP7_75t_L g3214 ( 
.A1(n_2631),
.A2(n_1718),
.B(n_1699),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2545),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2511),
.Y(n_3216)
);

AND2x6_ASAP7_75t_L g3217 ( 
.A(n_2635),
.B(n_915),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2531),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_2545),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_2808),
.B(n_1862),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2555),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2536),
.Y(n_3222)
);

INVx2_ASAP7_75t_L g3223 ( 
.A(n_2555),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_2834),
.B(n_1860),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2537),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2555),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_2808),
.B(n_905),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_2533),
.Y(n_3228)
);

AND2x2_ASAP7_75t_L g3229 ( 
.A(n_2635),
.B(n_1862),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2555),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2555),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2672),
.B(n_1860),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2631),
.Y(n_3233)
);

OR2x6_ASAP7_75t_L g3234 ( 
.A(n_2679),
.B(n_1378),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2548),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2632),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2554),
.Y(n_3237)
);

INVxp67_ASAP7_75t_L g3238 ( 
.A(n_2751),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2557),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2563),
.Y(n_3240)
);

CKINVDCx20_ASAP7_75t_R g3241 ( 
.A(n_2501),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_2642),
.B(n_1904),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2564),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_SL g3244 ( 
.A(n_2809),
.B(n_1904),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_2567),
.Y(n_3245)
);

OAI22xp5_ASAP7_75t_SL g3246 ( 
.A1(n_2451),
.A2(n_2116),
.B1(n_2119),
.B2(n_2105),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2632),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2569),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2636),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2636),
.Y(n_3250)
);

XNOR2xp5_ASAP7_75t_L g3251 ( 
.A(n_2670),
.B(n_2119),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_2638),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2642),
.B(n_1906),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_2669),
.B(n_1906),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2672),
.B(n_1868),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2657),
.B(n_1882),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2578),
.Y(n_3257)
);

INVxp67_ASAP7_75t_L g3258 ( 
.A(n_2760),
.Y(n_3258)
);

AND2x6_ASAP7_75t_L g3259 ( 
.A(n_2669),
.B(n_946),
.Y(n_3259)
);

INVx2_ASAP7_75t_L g3260 ( 
.A(n_2638),
.Y(n_3260)
);

AND2x2_ASAP7_75t_L g3261 ( 
.A(n_2671),
.B(n_1882),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2646),
.Y(n_3262)
);

BUFx2_ASAP7_75t_L g3263 ( 
.A(n_2882),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2646),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2647),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2647),
.Y(n_3266)
);

BUFx2_ASAP7_75t_L g3267 ( 
.A(n_2533),
.Y(n_3267)
);

OR2x2_ASAP7_75t_L g3268 ( 
.A(n_2881),
.B(n_1885),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2656),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2656),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2659),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2659),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2672),
.Y(n_3273)
);

OAI21x1_ASAP7_75t_L g3274 ( 
.A1(n_2595),
.A2(n_1624),
.B(n_1595),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_2673),
.Y(n_3275)
);

INVx2_ASAP7_75t_L g3276 ( 
.A(n_2673),
.Y(n_3276)
);

BUFx2_ASAP7_75t_L g3277 ( 
.A(n_2501),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2673),
.Y(n_3278)
);

BUFx2_ASAP7_75t_L g3279 ( 
.A(n_2655),
.Y(n_3279)
);

NAND2xp33_ASAP7_75t_SL g3280 ( 
.A(n_2809),
.B(n_1219),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_2675),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_2675),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2675),
.Y(n_3283)
);

HB1xp67_ASAP7_75t_L g3284 ( 
.A(n_2877),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2664),
.Y(n_3285)
);

HB1xp67_ASAP7_75t_L g3286 ( 
.A(n_2877),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2664),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2730),
.B(n_1885),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2595),
.Y(n_3289)
);

INVx3_ASAP7_75t_L g3290 ( 
.A(n_2427),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2595),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_2428),
.Y(n_3292)
);

INVx3_ASAP7_75t_L g3293 ( 
.A(n_2427),
.Y(n_3293)
);

INVx2_ASAP7_75t_L g3294 ( 
.A(n_2600),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_2600),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2600),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2616),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2616),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2616),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2651),
.Y(n_3300)
);

HB1xp67_ASAP7_75t_L g3301 ( 
.A(n_2877),
.Y(n_3301)
);

INVx3_ASAP7_75t_L g3302 ( 
.A(n_2427),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2651),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2651),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2653),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2734),
.B(n_1886),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_2809),
.B(n_2810),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2653),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2734),
.B(n_1888),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2653),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_2660),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_2660),
.Y(n_3312)
);

AND2x2_ASAP7_75t_L g3313 ( 
.A(n_2671),
.B(n_1891),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2660),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_2660),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2660),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_2662),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2662),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_2806),
.Y(n_3319)
);

INVx3_ASAP7_75t_L g3320 ( 
.A(n_2662),
.Y(n_3320)
);

BUFx3_ASAP7_75t_L g3321 ( 
.A(n_2422),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2662),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_2662),
.Y(n_3323)
);

INVx3_ASAP7_75t_L g3324 ( 
.A(n_2665),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_SL g3325 ( 
.A(n_2809),
.B(n_1891),
.Y(n_3325)
);

INVx3_ASAP7_75t_L g3326 ( 
.A(n_2665),
.Y(n_3326)
);

INVx1_ASAP7_75t_L g3327 ( 
.A(n_2665),
.Y(n_3327)
);

OAI21x1_ASAP7_75t_L g3328 ( 
.A1(n_2467),
.A2(n_1638),
.B(n_1624),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_2665),
.Y(n_3329)
);

OA21x2_ASAP7_75t_L g3330 ( 
.A1(n_2473),
.A2(n_1723),
.B(n_1721),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2665),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_2734),
.B(n_1888),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_2667),
.Y(n_3333)
);

INVx1_ASAP7_75t_SL g3334 ( 
.A(n_2655),
.Y(n_3334)
);

BUFx6f_ASAP7_75t_L g3335 ( 
.A(n_2428),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_2667),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_L g3337 ( 
.A(n_2745),
.B(n_1889),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_2667),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_2745),
.B(n_1889),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2667),
.Y(n_3340)
);

INVx2_ASAP7_75t_L g3341 ( 
.A(n_2667),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_2713),
.B(n_1913),
.Y(n_3342)
);

CKINVDCx20_ASAP7_75t_R g3343 ( 
.A(n_2714),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_2668),
.Y(n_3344)
);

BUFx6f_ASAP7_75t_L g3345 ( 
.A(n_2428),
.Y(n_3345)
);

AND2x4_ASAP7_75t_L g3346 ( 
.A(n_2809),
.B(n_905),
.Y(n_3346)
);

AND2x6_ASAP7_75t_L g3347 ( 
.A(n_2713),
.B(n_946),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2668),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_SL g3349 ( 
.A(n_2810),
.B(n_1914),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_2725),
.B(n_1914),
.Y(n_3350)
);

NAND2xp33_ASAP7_75t_SL g3351 ( 
.A(n_2810),
.B(n_1239),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_2668),
.Y(n_3352)
);

BUFx2_ASAP7_75t_L g3353 ( 
.A(n_2714),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2668),
.Y(n_3354)
);

AND2x2_ASAP7_75t_L g3355 ( 
.A(n_2725),
.B(n_1921),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2810),
.B(n_1921),
.Y(n_3356)
);

BUFx2_ASAP7_75t_L g3357 ( 
.A(n_2866),
.Y(n_3357)
);

BUFx6f_ASAP7_75t_L g3358 ( 
.A(n_2428),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2668),
.Y(n_3359)
);

BUFx3_ASAP7_75t_L g3360 ( 
.A(n_2422),
.Y(n_3360)
);

AND2x4_ASAP7_75t_L g3361 ( 
.A(n_2810),
.B(n_916),
.Y(n_3361)
);

BUFx8_ASAP7_75t_L g3362 ( 
.A(n_2791),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_2509),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_2509),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_2784),
.B(n_1930),
.Y(n_3365)
);

HB1xp67_ASAP7_75t_L g3366 ( 
.A(n_2877),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2581),
.Y(n_3367)
);

BUFx3_ASAP7_75t_L g3368 ( 
.A(n_2422),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_2582),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_2745),
.B(n_2431),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_2494),
.B(n_1898),
.Y(n_3371)
);

AND2x4_ASAP7_75t_L g3372 ( 
.A(n_2784),
.B(n_916),
.Y(n_3372)
);

INVx6_ASAP7_75t_L g3373 ( 
.A(n_2422),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_2984),
.A2(n_2771),
.B1(n_2821),
.B2(n_2593),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_2973),
.Y(n_3375)
);

BUFx10_ASAP7_75t_L g3376 ( 
.A(n_2905),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_2884),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3050),
.B(n_2593),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3233),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_2984),
.A2(n_2821),
.B1(n_2771),
.B2(n_2814),
.Y(n_3380)
);

BUFx6f_ASAP7_75t_L g3381 ( 
.A(n_2973),
.Y(n_3381)
);

OR2x6_ASAP7_75t_L g3382 ( 
.A(n_3079),
.B(n_2784),
.Y(n_3382)
);

INVx3_ASAP7_75t_L g3383 ( 
.A(n_2973),
.Y(n_3383)
);

INVx2_ASAP7_75t_L g3384 ( 
.A(n_3233),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3127),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_3236),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3127),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_2944),
.Y(n_3388)
);

INVx4_ASAP7_75t_L g3389 ( 
.A(n_3092),
.Y(n_3389)
);

AOI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3064),
.A2(n_2814),
.B1(n_2875),
.B2(n_2819),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3236),
.Y(n_3391)
);

CKINVDCx20_ASAP7_75t_R g3392 ( 
.A(n_3157),
.Y(n_3392)
);

INVx3_ASAP7_75t_L g3393 ( 
.A(n_2973),
.Y(n_3393)
);

BUFx4f_ASAP7_75t_L g3394 ( 
.A(n_3307),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_3256),
.B(n_2789),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3136),
.Y(n_3396)
);

OAI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_3291),
.A2(n_2823),
.B(n_2792),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3136),
.Y(n_3398)
);

OR2x6_ASAP7_75t_L g3399 ( 
.A(n_3079),
.B(n_2784),
.Y(n_3399)
);

BUFx6f_ASAP7_75t_SL g3400 ( 
.A(n_3111),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_3137),
.Y(n_3401)
);

INVxp33_ASAP7_75t_L g3402 ( 
.A(n_3251),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3032),
.B(n_2789),
.Y(n_3403)
);

CKINVDCx5p33_ASAP7_75t_R g3404 ( 
.A(n_2903),
.Y(n_3404)
);

INVx3_ASAP7_75t_L g3405 ( 
.A(n_2973),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_SL g3406 ( 
.A(n_3307),
.B(n_2850),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_3247),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3247),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_SL g3409 ( 
.A1(n_3064),
.A2(n_2728),
.B1(n_2644),
.B2(n_2608),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_SL g3410 ( 
.A(n_3307),
.B(n_2850),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_3092),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3137),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3288),
.B(n_2789),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_3249),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3180),
.B(n_2799),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3095),
.B(n_2429),
.Y(n_3416)
);

INVx1_ASAP7_75t_SL g3417 ( 
.A(n_2942),
.Y(n_3417)
);

INVx2_ASAP7_75t_L g3418 ( 
.A(n_3249),
.Y(n_3418)
);

NAND2xp33_ASAP7_75t_SL g3419 ( 
.A(n_2903),
.B(n_2850),
.Y(n_3419)
);

INVxp67_ASAP7_75t_SL g3420 ( 
.A(n_2944),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3250),
.Y(n_3421)
);

NOR2xp33_ASAP7_75t_L g3422 ( 
.A(n_2976),
.B(n_2429),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3138),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_2977),
.Y(n_3424)
);

INVx4_ASAP7_75t_L g3425 ( 
.A(n_3092),
.Y(n_3425)
);

AND3x2_ASAP7_75t_L g3426 ( 
.A(n_3142),
.B(n_2856),
.C(n_2791),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_2997),
.A2(n_2814),
.B1(n_2875),
.B2(n_2819),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3250),
.Y(n_3428)
);

INVxp67_ASAP7_75t_L g3429 ( 
.A(n_2947),
.Y(n_3429)
);

NOR2xp33_ASAP7_75t_L g3430 ( 
.A(n_2990),
.B(n_2508),
.Y(n_3430)
);

INVx2_ASAP7_75t_L g3431 ( 
.A(n_3252),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3138),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3141),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3252),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3260),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_2909),
.B(n_2799),
.Y(n_3436)
);

INVx2_ASAP7_75t_SL g3437 ( 
.A(n_2944),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3042),
.B(n_2799),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_3238),
.B(n_2508),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3042),
.B(n_2818),
.Y(n_3440)
);

INVx2_ASAP7_75t_SL g3441 ( 
.A(n_3373),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_L g3442 ( 
.A(n_3042),
.B(n_2818),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3260),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3141),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3143),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3264),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3143),
.Y(n_3447)
);

INVx2_ASAP7_75t_SL g3448 ( 
.A(n_3373),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_SL g3449 ( 
.A(n_3267),
.B(n_2850),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3047),
.B(n_2818),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_3264),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3151),
.Y(n_3452)
);

INVx1_ASAP7_75t_L g3453 ( 
.A(n_3151),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_SL g3454 ( 
.A(n_3267),
.B(n_2829),
.Y(n_3454)
);

AND3x2_ASAP7_75t_L g3455 ( 
.A(n_3030),
.B(n_2856),
.C(n_2703),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3155),
.Y(n_3456)
);

AO21x2_ASAP7_75t_L g3457 ( 
.A1(n_3096),
.A2(n_2496),
.B(n_2715),
.Y(n_3457)
);

OR2x6_ASAP7_75t_L g3458 ( 
.A(n_3111),
.B(n_2855),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3272),
.Y(n_3459)
);

BUFx10_ASAP7_75t_L g3460 ( 
.A(n_2920),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_SL g3461 ( 
.A(n_3111),
.B(n_2829),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_2910),
.B(n_2829),
.Y(n_3462)
);

AND2x2_ASAP7_75t_L g3463 ( 
.A(n_3050),
.B(n_2839),
.Y(n_3463)
);

INVx2_ASAP7_75t_L g3464 ( 
.A(n_3272),
.Y(n_3464)
);

AOI22xp33_ASAP7_75t_L g3465 ( 
.A1(n_2997),
.A2(n_2814),
.B1(n_2875),
.B2(n_2819),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_SL g3466 ( 
.A(n_2910),
.B(n_2841),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_SL g3467 ( 
.A(n_3306),
.B(n_2841),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3155),
.Y(n_3468)
);

BUFx2_ASAP7_75t_L g3469 ( 
.A(n_2942),
.Y(n_3469)
);

AND2x4_ASAP7_75t_L g3470 ( 
.A(n_3092),
.B(n_2877),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3262),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3047),
.B(n_2524),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_2884),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_SL g3474 ( 
.A(n_3309),
.B(n_2841),
.Y(n_3474)
);

AND2x2_ASAP7_75t_L g3475 ( 
.A(n_2898),
.B(n_2899),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3262),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_2885),
.Y(n_3477)
);

INVx2_ASAP7_75t_L g3478 ( 
.A(n_2885),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_3332),
.B(n_2841),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3265),
.Y(n_3480)
);

BUFx6f_ASAP7_75t_L g3481 ( 
.A(n_2977),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_2889),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_2889),
.Y(n_3483)
);

INVx3_ASAP7_75t_L g3484 ( 
.A(n_2977),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3047),
.B(n_3063),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3063),
.B(n_2510),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3265),
.Y(n_3487)
);

INVx4_ASAP7_75t_L g3488 ( 
.A(n_3092),
.Y(n_3488)
);

INVx3_ASAP7_75t_L g3489 ( 
.A(n_2977),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_2891),
.Y(n_3490)
);

INVx2_ASAP7_75t_L g3491 ( 
.A(n_2891),
.Y(n_3491)
);

BUFx3_ASAP7_75t_L g3492 ( 
.A(n_3321),
.Y(n_3492)
);

CKINVDCx5p33_ASAP7_75t_R g3493 ( 
.A(n_2920),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_SL g3494 ( 
.A(n_2931),
.B(n_2529),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3266),
.Y(n_3495)
);

INVx2_ASAP7_75t_L g3496 ( 
.A(n_2892),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3063),
.B(n_2539),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3370),
.B(n_2562),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3266),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_L g3500 ( 
.A1(n_3217),
.A2(n_2814),
.B1(n_2875),
.B2(n_2802),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_2892),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_2900),
.B(n_2822),
.Y(n_3502)
);

XNOR2xp5_ASAP7_75t_L g3503 ( 
.A(n_3251),
.B(n_2454),
.Y(n_3503)
);

NOR2xp33_ASAP7_75t_L g3504 ( 
.A(n_3258),
.B(n_2648),
.Y(n_3504)
);

INVx2_ASAP7_75t_L g3505 ( 
.A(n_2901),
.Y(n_3505)
);

NOR2xp33_ASAP7_75t_L g3506 ( 
.A(n_3033),
.B(n_2648),
.Y(n_3506)
);

BUFx6f_ASAP7_75t_L g3507 ( 
.A(n_2977),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_2901),
.Y(n_3508)
);

BUFx3_ASAP7_75t_L g3509 ( 
.A(n_3321),
.Y(n_3509)
);

OAI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3273),
.A2(n_2463),
.B1(n_2836),
.B2(n_2832),
.Y(n_3510)
);

BUFx3_ASAP7_75t_L g3511 ( 
.A(n_3360),
.Y(n_3511)
);

BUFx2_ASAP7_75t_L g3512 ( 
.A(n_3009),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_2922),
.Y(n_3513)
);

BUFx10_ASAP7_75t_L g3514 ( 
.A(n_2931),
.Y(n_3514)
);

AOI22xp33_ASAP7_75t_L g3515 ( 
.A1(n_3217),
.A2(n_2814),
.B1(n_2875),
.B2(n_2802),
.Y(n_3515)
);

INVx2_ASAP7_75t_L g3516 ( 
.A(n_2922),
.Y(n_3516)
);

BUFx2_ASAP7_75t_L g3517 ( 
.A(n_3009),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3269),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_SL g3519 ( 
.A(n_3337),
.B(n_2613),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3269),
.Y(n_3520)
);

INVx3_ASAP7_75t_L g3521 ( 
.A(n_3016),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3270),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_2929),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_2929),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3270),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_3271),
.Y(n_3526)
);

INVx2_ASAP7_75t_SL g3527 ( 
.A(n_3373),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_2937),
.Y(n_3528)
);

INVx3_ASAP7_75t_L g3529 ( 
.A(n_3016),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3271),
.Y(n_3530)
);

INVx3_ASAP7_75t_L g3531 ( 
.A(n_3016),
.Y(n_3531)
);

INVx2_ASAP7_75t_L g3532 ( 
.A(n_2937),
.Y(n_3532)
);

INVx4_ASAP7_75t_L g3533 ( 
.A(n_3161),
.Y(n_3533)
);

INVx2_ASAP7_75t_SL g3534 ( 
.A(n_3373),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_2949),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_L g3536 ( 
.A(n_3133),
.B(n_2658),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_2888),
.Y(n_3537)
);

INVx1_ASAP7_75t_SL g3538 ( 
.A(n_3114),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_2949),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_2953),
.Y(n_3540)
);

AND2x2_ASAP7_75t_L g3541 ( 
.A(n_2907),
.B(n_2839),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_2888),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3339),
.B(n_2613),
.Y(n_3543)
);

OAI22xp33_ASAP7_75t_L g3544 ( 
.A1(n_3041),
.A2(n_2658),
.B1(n_2702),
.B2(n_2697),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_2890),
.Y(n_3545)
);

INVx2_ASAP7_75t_SL g3546 ( 
.A(n_3360),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_2890),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_2953),
.Y(n_3548)
);

INVx4_ASAP7_75t_L g3549 ( 
.A(n_3161),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2915),
.B(n_2597),
.Y(n_3550)
);

NOR2xp33_ASAP7_75t_L g3551 ( 
.A(n_3148),
.B(n_2702),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_2916),
.B(n_2599),
.Y(n_3552)
);

NOR2xp33_ASAP7_75t_L g3553 ( 
.A(n_3175),
.B(n_2826),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_3061),
.B(n_2697),
.Y(n_3554)
);

BUFx3_ASAP7_75t_L g3555 ( 
.A(n_3368),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_2893),
.Y(n_3556)
);

BUFx3_ASAP7_75t_L g3557 ( 
.A(n_3368),
.Y(n_3557)
);

INVx3_ASAP7_75t_L g3558 ( 
.A(n_3016),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_2955),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_2954),
.B(n_2606),
.Y(n_3560)
);

INVx5_ASAP7_75t_L g3561 ( 
.A(n_3161),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_SL g3562 ( 
.A(n_3229),
.B(n_2780),
.Y(n_3562)
);

INVx2_ASAP7_75t_L g3563 ( 
.A(n_2955),
.Y(n_3563)
);

NAND3xp33_ASAP7_75t_SL g3564 ( 
.A(n_2936),
.B(n_2840),
.C(n_2854),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3229),
.B(n_2822),
.Y(n_3565)
);

INVx2_ASAP7_75t_SL g3566 ( 
.A(n_3228),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_L g3567 ( 
.A(n_3013),
.B(n_2847),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_2966),
.B(n_2988),
.Y(n_3568)
);

INVx3_ASAP7_75t_L g3569 ( 
.A(n_3016),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3242),
.B(n_2780),
.Y(n_3570)
);

INVx2_ASAP7_75t_L g3571 ( 
.A(n_2960),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2893),
.Y(n_3572)
);

INVx2_ASAP7_75t_L g3573 ( 
.A(n_2960),
.Y(n_3573)
);

BUFx6f_ASAP7_75t_L g3574 ( 
.A(n_3017),
.Y(n_3574)
);

INVx2_ASAP7_75t_L g3575 ( 
.A(n_2961),
.Y(n_3575)
);

BUFx3_ASAP7_75t_L g3576 ( 
.A(n_3017),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_2896),
.Y(n_3577)
);

NOR2xp33_ASAP7_75t_R g3578 ( 
.A(n_2936),
.B(n_2840),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_2896),
.Y(n_3579)
);

CKINVDCx6p67_ASAP7_75t_R g3580 ( 
.A(n_3015),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2908),
.Y(n_3581)
);

INVx2_ASAP7_75t_SL g3582 ( 
.A(n_3017),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_2908),
.Y(n_3583)
);

INVx3_ASAP7_75t_L g3584 ( 
.A(n_3017),
.Y(n_3584)
);

INVx4_ASAP7_75t_L g3585 ( 
.A(n_3177),
.Y(n_3585)
);

INVx4_ASAP7_75t_L g3586 ( 
.A(n_3177),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3232),
.B(n_2611),
.Y(n_3587)
);

CKINVDCx5p33_ASAP7_75t_R g3588 ( 
.A(n_3200),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_2961),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_2974),
.Y(n_3590)
);

NOR2xp33_ASAP7_75t_L g3591 ( 
.A(n_3027),
.B(n_2847),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_2911),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_3242),
.B(n_2785),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_2911),
.Y(n_3594)
);

INVx8_ASAP7_75t_L g3595 ( 
.A(n_3217),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3066),
.B(n_2847),
.Y(n_3596)
);

BUFx4f_ASAP7_75t_L g3597 ( 
.A(n_3217),
.Y(n_3597)
);

INVx5_ASAP7_75t_L g3598 ( 
.A(n_3177),
.Y(n_3598)
);

BUFx3_ASAP7_75t_L g3599 ( 
.A(n_3017),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_2974),
.Y(n_3600)
);

OAI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_2894),
.A2(n_2849),
.B1(n_2836),
.B2(n_2832),
.Y(n_3601)
);

NOR2xp33_ASAP7_75t_L g3602 ( 
.A(n_3067),
.B(n_2847),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_2917),
.Y(n_3603)
);

INVx2_ASAP7_75t_SL g3604 ( 
.A(n_3035),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_2975),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_2917),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_2975),
.Y(n_3607)
);

OR2x6_ASAP7_75t_L g3608 ( 
.A(n_3015),
.B(n_2855),
.Y(n_3608)
);

INVx2_ASAP7_75t_SL g3609 ( 
.A(n_3035),
.Y(n_3609)
);

INVxp33_ASAP7_75t_L g3610 ( 
.A(n_2921),
.Y(n_3610)
);

AOI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3217),
.A2(n_2498),
.B1(n_2573),
.B2(n_2484),
.Y(n_3611)
);

OR2x2_ASAP7_75t_L g3612 ( 
.A(n_3334),
.B(n_2925),
.Y(n_3612)
);

NOR2xp33_ASAP7_75t_L g3613 ( 
.A(n_3086),
.B(n_2587),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2918),
.Y(n_3614)
);

INVx2_ASAP7_75t_L g3615 ( 
.A(n_2978),
.Y(n_3615)
);

INVx2_ASAP7_75t_L g3616 ( 
.A(n_2978),
.Y(n_3616)
);

INVxp33_ASAP7_75t_L g3617 ( 
.A(n_3165),
.Y(n_3617)
);

INVx3_ASAP7_75t_L g3618 ( 
.A(n_3035),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_2918),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3371),
.B(n_2779),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_3253),
.B(n_2786),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_2979),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3255),
.B(n_2620),
.Y(n_3623)
);

NAND2xp5_ASAP7_75t_L g3624 ( 
.A(n_3153),
.B(n_2637),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3253),
.B(n_2785),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_2923),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_2979),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_2923),
.Y(n_3628)
);

INVx4_ASAP7_75t_L g3629 ( 
.A(n_3201),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_SL g3630 ( 
.A(n_3254),
.B(n_2793),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_3153),
.B(n_2681),
.Y(n_3631)
);

BUFx3_ASAP7_75t_L g3632 ( 
.A(n_3035),
.Y(n_3632)
);

INVx3_ASAP7_75t_L g3633 ( 
.A(n_3035),
.Y(n_3633)
);

INVx2_ASAP7_75t_L g3634 ( 
.A(n_2993),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_2926),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_2993),
.Y(n_3636)
);

BUFx2_ASAP7_75t_L g3637 ( 
.A(n_3114),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3153),
.B(n_2701),
.Y(n_3638)
);

OR2x6_ASAP7_75t_L g3639 ( 
.A(n_3174),
.B(n_2855),
.Y(n_3639)
);

AND2x2_ASAP7_75t_L g3640 ( 
.A(n_3254),
.B(n_3261),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_3200),
.Y(n_3641)
);

INVx5_ASAP7_75t_L g3642 ( 
.A(n_3201),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_2994),
.Y(n_3643)
);

OR2x2_ASAP7_75t_L g3644 ( 
.A(n_3277),
.B(n_2876),
.Y(n_3644)
);

INVx2_ASAP7_75t_SL g3645 ( 
.A(n_2883),
.Y(n_3645)
);

INVx3_ASAP7_75t_L g3646 ( 
.A(n_3201),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_2926),
.Y(n_3647)
);

INVx3_ASAP7_75t_L g3648 ( 
.A(n_3208),
.Y(n_3648)
);

CKINVDCx5p33_ASAP7_75t_R g3649 ( 
.A(n_3319),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_2928),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3160),
.B(n_2692),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_2928),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_2930),
.Y(n_3653)
);

AOI22xp33_ASAP7_75t_L g3654 ( 
.A1(n_3217),
.A2(n_2875),
.B1(n_2802),
.B2(n_2881),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_2930),
.Y(n_3655)
);

AOI22xp33_ASAP7_75t_L g3656 ( 
.A1(n_3259),
.A2(n_3347),
.B1(n_3351),
.B2(n_3280),
.Y(n_3656)
);

INVx3_ASAP7_75t_L g3657 ( 
.A(n_3208),
.Y(n_3657)
);

INVx2_ASAP7_75t_SL g3658 ( 
.A(n_2883),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_2994),
.Y(n_3659)
);

BUFx4f_ASAP7_75t_L g3660 ( 
.A(n_3259),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_2933),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3160),
.B(n_2733),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3160),
.B(n_2733),
.Y(n_3663)
);

BUFx6f_ASAP7_75t_SL g3664 ( 
.A(n_3174),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_2996),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_2996),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_2933),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_2934),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_2934),
.Y(n_3669)
);

INVx5_ASAP7_75t_L g3670 ( 
.A(n_3208),
.Y(n_3670)
);

INVx3_ASAP7_75t_L g3671 ( 
.A(n_3046),
.Y(n_3671)
);

INVx1_ASAP7_75t_L g3672 ( 
.A(n_2951),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_2883),
.Y(n_3673)
);

NOR2xp33_ASAP7_75t_L g3674 ( 
.A(n_3261),
.B(n_2813),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_2951),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3313),
.B(n_2815),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_2998),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_2998),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3001),
.Y(n_3679)
);

INVx3_ASAP7_75t_L g3680 ( 
.A(n_3046),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_3313),
.B(n_2874),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_SL g3682 ( 
.A(n_3342),
.B(n_2793),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_2952),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3178),
.B(n_2736),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3001),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3006),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_2952),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_2883),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_2965),
.Y(n_3689)
);

HB1xp67_ASAP7_75t_L g3690 ( 
.A(n_3277),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_L g3691 ( 
.A(n_3289),
.B(n_2796),
.Y(n_3691)
);

OAI22xp5_ASAP7_75t_L g3692 ( 
.A1(n_3273),
.A2(n_2463),
.B1(n_2805),
.B2(n_2796),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3006),
.Y(n_3693)
);

INVxp33_ASAP7_75t_L g3694 ( 
.A(n_3202),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3342),
.B(n_2844),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_2965),
.Y(n_3696)
);

AOI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3036),
.A2(n_2823),
.B(n_2792),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_2967),
.Y(n_3698)
);

INVxp33_ASAP7_75t_L g3699 ( 
.A(n_3202),
.Y(n_3699)
);

INVx4_ASAP7_75t_L g3700 ( 
.A(n_3046),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_2967),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_SL g3702 ( 
.A(n_3350),
.B(n_2805),
.Y(n_3702)
);

NAND3x1_ASAP7_75t_L g3703 ( 
.A(n_3350),
.B(n_2868),
.C(n_2844),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3007),
.Y(n_3704)
);

AOI22xp5_ASAP7_75t_L g3705 ( 
.A1(n_3259),
.A2(n_2498),
.B1(n_2573),
.B2(n_2484),
.Y(n_3705)
);

NAND2xp33_ASAP7_75t_L g3706 ( 
.A(n_3289),
.B(n_2816),
.Y(n_3706)
);

INVx3_ASAP7_75t_L g3707 ( 
.A(n_3046),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_SL g3708 ( 
.A(n_3355),
.B(n_2816),
.Y(n_3708)
);

AND2x2_ASAP7_75t_L g3709 ( 
.A(n_3355),
.B(n_2736),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3007),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_2968),
.Y(n_3711)
);

NAND3xp33_ASAP7_75t_L g3712 ( 
.A(n_2980),
.B(n_2727),
.C(n_2720),
.Y(n_3712)
);

BUFx8_ASAP7_75t_SL g3713 ( 
.A(n_3319),
.Y(n_3713)
);

INVx3_ASAP7_75t_L g3714 ( 
.A(n_3046),
.Y(n_3714)
);

INVx8_ASAP7_75t_L g3715 ( 
.A(n_3259),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3008),
.Y(n_3716)
);

OAI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_3281),
.A2(n_2463),
.B1(n_2824),
.B2(n_2844),
.Y(n_3717)
);

AOI22xp33_ASAP7_75t_SL g3718 ( 
.A1(n_3246),
.A2(n_2538),
.B1(n_2502),
.B2(n_2481),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_2968),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_2969),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_2969),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3008),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_3212),
.B(n_2845),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3011),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_SL g3725 ( 
.A(n_2935),
.B(n_2824),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_2972),
.Y(n_3726)
);

AND2x6_ASAP7_75t_L g3727 ( 
.A(n_3096),
.B(n_2849),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3011),
.Y(n_3728)
);

AOI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_3259),
.A2(n_3347),
.B1(n_2498),
.B2(n_2573),
.Y(n_3729)
);

AND2x2_ASAP7_75t_L g3730 ( 
.A(n_3103),
.B(n_2640),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3259),
.A2(n_2881),
.B1(n_2624),
.B2(n_2630),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3022),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_2972),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_2981),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_2981),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3022),
.Y(n_3736)
);

INVx2_ASAP7_75t_L g3737 ( 
.A(n_3130),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3130),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_2897),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3178),
.B(n_2712),
.Y(n_3740)
);

AOI22xp5_ASAP7_75t_L g3741 ( 
.A1(n_3347),
.A2(n_2498),
.B1(n_2573),
.B2(n_2484),
.Y(n_3741)
);

INVx3_ASAP7_75t_L g3742 ( 
.A(n_3055),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3130),
.Y(n_3743)
);

BUFx10_ASAP7_75t_L g3744 ( 
.A(n_3091),
.Y(n_3744)
);

NOR2xp33_ASAP7_75t_L g3745 ( 
.A(n_3212),
.B(n_2853),
.Y(n_3745)
);

INVx2_ASAP7_75t_L g3746 ( 
.A(n_2986),
.Y(n_3746)
);

AND3x2_ASAP7_75t_L g3747 ( 
.A(n_3279),
.B(n_3357),
.C(n_3353),
.Y(n_3747)
);

BUFx2_ASAP7_75t_L g3748 ( 
.A(n_3241),
.Y(n_3748)
);

CKINVDCx6p67_ASAP7_75t_R g3749 ( 
.A(n_3241),
.Y(n_3749)
);

BUFx2_ASAP7_75t_L g3750 ( 
.A(n_3343),
.Y(n_3750)
);

OAI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3010),
.A2(n_3024),
.B1(n_3026),
.B2(n_3019),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_2986),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_2987),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_L g3754 ( 
.A(n_3178),
.B(n_2712),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_SL g3755 ( 
.A(n_3103),
.B(n_2848),
.Y(n_3755)
);

OAI21xp33_ASAP7_75t_SL g3756 ( 
.A1(n_3281),
.A2(n_2605),
.B(n_2594),
.Y(n_3756)
);

CKINVDCx6p67_ASAP7_75t_R g3757 ( 
.A(n_3343),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_2987),
.Y(n_3758)
);

INVx2_ASAP7_75t_SL g3759 ( 
.A(n_2883),
.Y(n_3759)
);

INVx4_ASAP7_75t_L g3760 ( 
.A(n_3055),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_2991),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_2991),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_2992),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3038),
.B(n_2858),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_2992),
.Y(n_3765)
);

AO21x2_ASAP7_75t_L g3766 ( 
.A1(n_3104),
.A2(n_2744),
.B(n_2740),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_2995),
.Y(n_3767)
);

INVx4_ASAP7_75t_L g3768 ( 
.A(n_3055),
.Y(n_3768)
);

BUFx6f_ASAP7_75t_L g3769 ( 
.A(n_3055),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_2995),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3000),
.Y(n_3771)
);

OAI21xp33_ASAP7_75t_SL g3772 ( 
.A1(n_3282),
.A2(n_2615),
.B(n_2607),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3000),
.Y(n_3773)
);

NOR2xp33_ASAP7_75t_L g3774 ( 
.A(n_3056),
.B(n_2859),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3003),
.Y(n_3775)
);

AND2x2_ASAP7_75t_L g3776 ( 
.A(n_3128),
.B(n_2640),
.Y(n_3776)
);

INVx3_ASAP7_75t_L g3777 ( 
.A(n_3055),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3003),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3005),
.Y(n_3779)
);

AOI22xp5_ASAP7_75t_L g3780 ( 
.A1(n_3347),
.A2(n_2498),
.B1(n_2573),
.B2(n_2484),
.Y(n_3780)
);

AND2x2_ASAP7_75t_L g3781 ( 
.A(n_3128),
.B(n_2640),
.Y(n_3781)
);

NAND2xp33_ASAP7_75t_L g3782 ( 
.A(n_3294),
.B(n_2827),
.Y(n_3782)
);

BUFx3_ASAP7_75t_L g3783 ( 
.A(n_2906),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3005),
.Y(n_3784)
);

OAI22xp33_ASAP7_75t_SL g3785 ( 
.A1(n_3206),
.A2(n_2457),
.B1(n_1272),
.B2(n_1259),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_SL g3786 ( 
.A(n_3134),
.B(n_2848),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3206),
.B(n_2712),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3014),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3014),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_SL g3790 ( 
.A(n_3134),
.B(n_2851),
.Y(n_3790)
);

INVx2_ASAP7_75t_L g3791 ( 
.A(n_3018),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3206),
.B(n_2516),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3018),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3021),
.Y(n_3794)
);

AO22x2_ASAP7_75t_L g3795 ( 
.A1(n_3372),
.A2(n_3346),
.B1(n_3361),
.B2(n_3227),
.Y(n_3795)
);

AND2x2_ASAP7_75t_L g3796 ( 
.A(n_3146),
.B(n_2516),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3021),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_SL g3798 ( 
.A(n_3146),
.B(n_2851),
.Y(n_3798)
);

CKINVDCx20_ASAP7_75t_R g3799 ( 
.A(n_3157),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3023),
.Y(n_3800)
);

INVx2_ASAP7_75t_SL g3801 ( 
.A(n_2906),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3049),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3062),
.B(n_2833),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3049),
.Y(n_3804)
);

CKINVDCx5p33_ASAP7_75t_R g3805 ( 
.A(n_2897),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_3227),
.B(n_2541),
.Y(n_3806)
);

BUFx3_ASAP7_75t_L g3807 ( 
.A(n_2906),
.Y(n_3807)
);

NOR2xp33_ASAP7_75t_R g3808 ( 
.A(n_3154),
.B(n_2529),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3023),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3054),
.Y(n_3810)
);

CKINVDCx5p33_ASAP7_75t_R g3811 ( 
.A(n_2950),
.Y(n_3811)
);

NOR2x1p5_ASAP7_75t_L g3812 ( 
.A(n_3268),
.B(n_2683),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3025),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3054),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3057),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_SL g3816 ( 
.A(n_3147),
.B(n_2800),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3025),
.Y(n_3817)
);

INVx5_ASAP7_75t_L g3818 ( 
.A(n_2895),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3057),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3147),
.B(n_2828),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_SL g3821 ( 
.A(n_3190),
.B(n_2835),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3028),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_SL g3823 ( 
.A(n_3190),
.B(n_2521),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3059),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3227),
.B(n_2541),
.Y(n_3825)
);

OAI22xp33_ASAP7_75t_L g3826 ( 
.A1(n_3069),
.A2(n_2746),
.B1(n_2752),
.B2(n_2556),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3059),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3028),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3285),
.Y(n_3829)
);

CKINVDCx5p33_ASAP7_75t_R g3830 ( 
.A(n_2950),
.Y(n_3830)
);

BUFx6f_ASAP7_75t_SL g3831 ( 
.A(n_3174),
.Y(n_3831)
);

AOI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3036),
.A2(n_2823),
.B(n_2792),
.Y(n_3832)
);

BUFx6f_ASAP7_75t_L g3833 ( 
.A(n_3060),
.Y(n_3833)
);

AO22x2_ASAP7_75t_L g3834 ( 
.A1(n_3372),
.A2(n_2619),
.B1(n_2863),
.B2(n_2857),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3285),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_SL g3836 ( 
.A(n_3088),
.B(n_2843),
.Y(n_3836)
);

AND2x6_ASAP7_75t_L g3837 ( 
.A(n_3104),
.B(n_2741),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3214),
.Y(n_3838)
);

INVx4_ASAP7_75t_L g3839 ( 
.A(n_3060),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_SL g3840 ( 
.A(n_3088),
.B(n_2855),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3287),
.Y(n_3841)
);

INVx2_ASAP7_75t_L g3842 ( 
.A(n_3214),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3214),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3287),
.Y(n_3844)
);

BUFx6f_ASAP7_75t_SL g3845 ( 
.A(n_3174),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3065),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3089),
.B(n_2568),
.Y(n_3847)
);

AO22x1_ASAP7_75t_L g3848 ( 
.A1(n_3347),
.A2(n_2484),
.B1(n_2573),
.B2(n_2498),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3291),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3065),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3073),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3295),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_L g3853 ( 
.A(n_3346),
.B(n_2568),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3089),
.B(n_2855),
.Y(n_3854)
);

CKINVDCx6p67_ASAP7_75t_R g3855 ( 
.A(n_3234),
.Y(n_3855)
);

AOI22xp5_ASAP7_75t_L g3856 ( 
.A1(n_3347),
.A2(n_2484),
.B1(n_2624),
.B2(n_2604),
.Y(n_3856)
);

BUFx6f_ASAP7_75t_L g3857 ( 
.A(n_3060),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3295),
.Y(n_3858)
);

INVx2_ASAP7_75t_SL g3859 ( 
.A(n_2906),
.Y(n_3859)
);

INVx2_ASAP7_75t_L g3860 ( 
.A(n_3073),
.Y(n_3860)
);

AO21x2_ASAP7_75t_L g3861 ( 
.A1(n_3105),
.A2(n_3087),
.B(n_3084),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3132),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3346),
.B(n_3361),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3296),
.Y(n_3864)
);

INVx3_ASAP7_75t_L g3865 ( 
.A(n_3060),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3132),
.Y(n_3866)
);

NOR2x1p5_ASAP7_75t_L g3867 ( 
.A(n_3268),
.B(n_2683),
.Y(n_3867)
);

CKINVDCx5p33_ASAP7_75t_R g3868 ( 
.A(n_2950),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3361),
.B(n_2749),
.Y(n_3869)
);

OR2x2_ASAP7_75t_L g3870 ( 
.A(n_3279),
.B(n_2878),
.Y(n_3870)
);

INVx4_ASAP7_75t_L g3871 ( 
.A(n_3060),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3132),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3210),
.Y(n_3873)
);

INVx2_ASAP7_75t_SL g3874 ( 
.A(n_2906),
.Y(n_3874)
);

NOR2xp33_ASAP7_75t_L g3875 ( 
.A(n_2886),
.B(n_2532),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3210),
.Y(n_3876)
);

INVx3_ASAP7_75t_L g3877 ( 
.A(n_3070),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_2887),
.B(n_2532),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3210),
.Y(n_3879)
);

AND3x2_ASAP7_75t_L g3880 ( 
.A(n_3353),
.B(n_2863),
.C(n_2857),
.Y(n_3880)
);

CKINVDCx5p33_ASAP7_75t_R g3881 ( 
.A(n_3154),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3296),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3297),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_3275),
.Y(n_3884)
);

BUFx3_ASAP7_75t_L g3885 ( 
.A(n_2913),
.Y(n_3885)
);

INVx4_ASAP7_75t_L g3886 ( 
.A(n_3070),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_3070),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3297),
.Y(n_3888)
);

INVx4_ASAP7_75t_L g3889 ( 
.A(n_3070),
.Y(n_3889)
);

INVxp67_ASAP7_75t_L g3890 ( 
.A(n_3357),
.Y(n_3890)
);

BUFx10_ASAP7_75t_L g3891 ( 
.A(n_3091),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3275),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3298),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_2887),
.B(n_2741),
.Y(n_3894)
);

NOR2xp33_ASAP7_75t_L g3895 ( 
.A(n_2938),
.B(n_2561),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3298),
.Y(n_3896)
);

AO21x2_ASAP7_75t_L g3897 ( 
.A1(n_3105),
.A2(n_2755),
.B(n_2731),
.Y(n_3897)
);

BUFx3_ASAP7_75t_L g3898 ( 
.A(n_2913),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_SL g3899 ( 
.A(n_2945),
.B(n_2474),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3299),
.Y(n_3900)
);

AND2x2_ASAP7_75t_SL g3901 ( 
.A(n_3372),
.B(n_946),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3299),
.Y(n_3902)
);

NAND3xp33_ASAP7_75t_L g3903 ( 
.A(n_3081),
.B(n_2603),
.C(n_2441),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3152),
.B(n_2474),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3303),
.Y(n_3905)
);

INVx1_ASAP7_75t_L g3906 ( 
.A(n_3303),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3304),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3276),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3169),
.B(n_2749),
.Y(n_3909)
);

INVxp67_ASAP7_75t_L g3910 ( 
.A(n_3164),
.Y(n_3910)
);

NOR2x1p5_ASAP7_75t_L g3911 ( 
.A(n_3091),
.B(n_2758),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3304),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3276),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_SL g3914 ( 
.A1(n_3234),
.A2(n_2738),
.B1(n_2776),
.B2(n_2804),
.Y(n_3914)
);

INVx5_ASAP7_75t_L g3915 ( 
.A(n_2895),
.Y(n_3915)
);

BUFx6f_ASAP7_75t_L g3916 ( 
.A(n_3070),
.Y(n_3916)
);

AND2x4_ASAP7_75t_L g3917 ( 
.A(n_2912),
.B(n_2763),
.Y(n_3917)
);

AND2x4_ASAP7_75t_L g3918 ( 
.A(n_2912),
.B(n_2957),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3278),
.Y(n_3919)
);

NOR2xp33_ASAP7_75t_L g3920 ( 
.A(n_3170),
.B(n_2561),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3305),
.Y(n_3921)
);

INVx4_ASAP7_75t_L g3922 ( 
.A(n_3072),
.Y(n_3922)
);

INVx3_ASAP7_75t_L g3923 ( 
.A(n_3072),
.Y(n_3923)
);

AOI21x1_ASAP7_75t_L g3924 ( 
.A1(n_3031),
.A2(n_1734),
.B(n_1730),
.Y(n_3924)
);

INVx2_ASAP7_75t_SL g3925 ( 
.A(n_2913),
.Y(n_3925)
);

BUFx3_ASAP7_75t_L g3926 ( 
.A(n_2913),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3305),
.Y(n_3927)
);

INVx3_ASAP7_75t_L g3928 ( 
.A(n_3072),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3171),
.B(n_2763),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3308),
.Y(n_3930)
);

NOR2xp33_ASAP7_75t_L g3931 ( 
.A(n_3158),
.B(n_2716),
.Y(n_3931)
);

INVx2_ASAP7_75t_L g3932 ( 
.A(n_3278),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3283),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3308),
.Y(n_3934)
);

NAND2xp5_ASAP7_75t_SL g3935 ( 
.A(n_3176),
.B(n_2676),
.Y(n_3935)
);

INVx1_ASAP7_75t_SL g3936 ( 
.A(n_3097),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_2983),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3283),
.Y(n_3938)
);

CKINVDCx20_ASAP7_75t_R g3939 ( 
.A(n_2983),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3294),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3300),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3181),
.B(n_2726),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3300),
.Y(n_3943)
);

NAND2xp5_ASAP7_75t_L g3944 ( 
.A(n_3182),
.B(n_2726),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3917),
.B(n_3158),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3475),
.Y(n_3946)
);

OR2x2_ASAP7_75t_L g3947 ( 
.A(n_3538),
.B(n_2871),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3746),
.Y(n_3948)
);

NAND2x1p5_ASAP7_75t_L g3949 ( 
.A(n_3394),
.B(n_3320),
.Y(n_3949)
);

INVx1_ASAP7_75t_L g3950 ( 
.A(n_3475),
.Y(n_3950)
);

NOR2xp33_ASAP7_75t_L g3951 ( 
.A(n_3621),
.B(n_2716),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3385),
.Y(n_3952)
);

AND2x2_ASAP7_75t_L g3953 ( 
.A(n_3709),
.B(n_2553),
.Y(n_3953)
);

XNOR2x2_ASAP7_75t_L g3954 ( 
.A(n_3503),
.B(n_2677),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3385),
.Y(n_3955)
);

XOR2xp5_ASAP7_75t_L g3956 ( 
.A(n_3503),
.B(n_2866),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3387),
.Y(n_3957)
);

XOR2x2_ASAP7_75t_L g3958 ( 
.A(n_3455),
.B(n_2869),
.Y(n_3958)
);

CKINVDCx20_ASAP7_75t_R g3959 ( 
.A(n_3713),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3387),
.Y(n_3960)
);

AND2x2_ASAP7_75t_L g3961 ( 
.A(n_3709),
.B(n_3640),
.Y(n_3961)
);

AND2x4_ASAP7_75t_L g3962 ( 
.A(n_3917),
.B(n_3263),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3396),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3640),
.B(n_3263),
.Y(n_3964)
);

AND2x4_ASAP7_75t_L g3965 ( 
.A(n_3917),
.B(n_3184),
.Y(n_3965)
);

NOR2xp33_ASAP7_75t_L g3966 ( 
.A(n_3674),
.B(n_3676),
.Y(n_3966)
);

INVx8_ASAP7_75t_L g3967 ( 
.A(n_3400),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3681),
.B(n_2871),
.Y(n_3968)
);

XNOR2x2_ASAP7_75t_L g3969 ( 
.A(n_3834),
.B(n_2677),
.Y(n_3969)
);

INVx2_ASAP7_75t_L g3970 ( 
.A(n_3746),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3396),
.Y(n_3971)
);

XOR2xp5_ASAP7_75t_L g3972 ( 
.A(n_3404),
.B(n_2122),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3565),
.B(n_3099),
.Y(n_3973)
);

XOR2xp5_ASAP7_75t_L g3974 ( 
.A(n_3493),
.B(n_2122),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3398),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3398),
.Y(n_3976)
);

INVx4_ASAP7_75t_L g3977 ( 
.A(n_3394),
.Y(n_3977)
);

INVx2_ASAP7_75t_SL g3978 ( 
.A(n_3578),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3401),
.Y(n_3979)
);

NOR2xp33_ASAP7_75t_L g3980 ( 
.A(n_3422),
.B(n_2787),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3401),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3412),
.Y(n_3982)
);

CKINVDCx5p33_ASAP7_75t_R g3983 ( 
.A(n_3808),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3412),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3423),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3620),
.B(n_3282),
.Y(n_3986)
);

CKINVDCx5p33_ASAP7_75t_R g3987 ( 
.A(n_3588),
.Y(n_3987)
);

NOR2xp33_ASAP7_75t_L g3988 ( 
.A(n_3723),
.B(n_2788),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3803),
.B(n_2919),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3637),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3423),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3432),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3565),
.B(n_3099),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3432),
.Y(n_3994)
);

NOR2xp33_ASAP7_75t_L g3995 ( 
.A(n_3745),
.B(n_2795),
.Y(n_3995)
);

NOR2xp67_ASAP7_75t_L g3996 ( 
.A(n_3564),
.B(n_2758),
.Y(n_3996)
);

NAND2x1p5_ASAP7_75t_L g3997 ( 
.A(n_3394),
.B(n_3320),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3433),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_3796),
.B(n_3099),
.Y(n_3999)
);

XOR2xp5_ASAP7_75t_L g4000 ( 
.A(n_3641),
.B(n_2141),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3758),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3433),
.Y(n_4002)
);

OR2x6_ASAP7_75t_L g4003 ( 
.A(n_3595),
.B(n_2807),
.Y(n_4003)
);

INVx1_ASAP7_75t_L g4004 ( 
.A(n_3444),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3444),
.Y(n_4005)
);

INVxp33_ASAP7_75t_L g4006 ( 
.A(n_3504),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3445),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3445),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3447),
.Y(n_4009)
);

XOR2xp5_ASAP7_75t_L g4010 ( 
.A(n_3649),
.B(n_2141),
.Y(n_4010)
);

INVxp67_ASAP7_75t_SL g4011 ( 
.A(n_3795),
.Y(n_4011)
);

INVxp67_ASAP7_75t_SL g4012 ( 
.A(n_3795),
.Y(n_4012)
);

BUFx6f_ASAP7_75t_L g4013 ( 
.A(n_3769),
.Y(n_4013)
);

XNOR2xp5_ASAP7_75t_L g4014 ( 
.A(n_3392),
.B(n_2148),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3769),
.Y(n_4015)
);

NOR2xp33_ASAP7_75t_L g4016 ( 
.A(n_3694),
.B(n_2797),
.Y(n_4016)
);

AND2x6_ASAP7_75t_L g4017 ( 
.A(n_3729),
.B(n_2941),
.Y(n_4017)
);

INVxp67_ASAP7_75t_L g4018 ( 
.A(n_3637),
.Y(n_4018)
);

AND2x6_ASAP7_75t_L g4019 ( 
.A(n_3729),
.B(n_2941),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3447),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3452),
.Y(n_4021)
);

BUFx6f_ASAP7_75t_L g4022 ( 
.A(n_3769),
.Y(n_4022)
);

AOI21xp5_ASAP7_75t_L g4023 ( 
.A1(n_3403),
.A2(n_3034),
.B(n_3031),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3452),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3453),
.Y(n_4025)
);

XOR2xp5_ASAP7_75t_L g4026 ( 
.A(n_3939),
.B(n_2148),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3796),
.B(n_3145),
.Y(n_4027)
);

CKINVDCx16_ASAP7_75t_R g4028 ( 
.A(n_3494),
.Y(n_4028)
);

CKINVDCx20_ASAP7_75t_R g4029 ( 
.A(n_3580),
.Y(n_4029)
);

XNOR2x1_ASAP7_75t_L g4030 ( 
.A(n_3834),
.B(n_2854),
.Y(n_4030)
);

NAND2xp33_ASAP7_75t_R g4031 ( 
.A(n_3881),
.B(n_2868),
.Y(n_4031)
);

NOR2xp33_ASAP7_75t_L g4032 ( 
.A(n_3699),
.B(n_2798),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_3847),
.B(n_3145),
.Y(n_4033)
);

NOR2xp33_ASAP7_75t_SL g4034 ( 
.A(n_3416),
.B(n_2807),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3453),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_SL g4036 ( 
.A(n_3561),
.B(n_3320),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3456),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3456),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3847),
.B(n_3145),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_L g4040 ( 
.A(n_3472),
.B(n_2458),
.Y(n_4040)
);

CKINVDCx5p33_ASAP7_75t_R g4041 ( 
.A(n_3739),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3468),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3758),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3468),
.Y(n_4044)
);

INVx2_ASAP7_75t_SL g4045 ( 
.A(n_3512),
.Y(n_4045)
);

NOR2xp33_ASAP7_75t_L g4046 ( 
.A(n_3506),
.B(n_2864),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3471),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3471),
.Y(n_4048)
);

NOR2xp33_ASAP7_75t_L g4049 ( 
.A(n_3764),
.B(n_2846),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3476),
.Y(n_4050)
);

NAND2xp33_ASAP7_75t_R g4051 ( 
.A(n_3805),
.B(n_2868),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3476),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3480),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3480),
.Y(n_4054)
);

INVx1_ASAP7_75t_L g4055 ( 
.A(n_3487),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3774),
.B(n_2696),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3730),
.B(n_2530),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3487),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3495),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3495),
.Y(n_4060)
);

XOR2x2_ASAP7_75t_L g4061 ( 
.A(n_3426),
.B(n_2869),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3499),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3499),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3518),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3518),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3520),
.Y(n_4066)
);

AND2x2_ASAP7_75t_L g4067 ( 
.A(n_3730),
.B(n_3234),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3520),
.Y(n_4068)
);

AO21x1_ASAP7_75t_L g4069 ( 
.A1(n_3413),
.A2(n_3224),
.B(n_3311),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3522),
.Y(n_4070)
);

CKINVDCx5p33_ASAP7_75t_R g4071 ( 
.A(n_3580),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3522),
.Y(n_4072)
);

INVx1_ASAP7_75t_L g4073 ( 
.A(n_3525),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3525),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3526),
.Y(n_4075)
);

XNOR2x2_ASAP7_75t_L g4076 ( 
.A(n_3834),
.B(n_2865),
.Y(n_4076)
);

INVxp67_ASAP7_75t_SL g4077 ( 
.A(n_3795),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3761),
.Y(n_4078)
);

INVx2_ASAP7_75t_SL g4079 ( 
.A(n_3512),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_3761),
.Y(n_4080)
);

NOR2xp33_ASAP7_75t_L g4081 ( 
.A(n_3895),
.B(n_2478),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3526),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3776),
.B(n_3781),
.Y(n_4083)
);

BUFx6f_ASAP7_75t_L g4084 ( 
.A(n_3769),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_3530),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3530),
.Y(n_4086)
);

NOR2xp33_ASAP7_75t_L g4087 ( 
.A(n_3878),
.B(n_3112),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3829),
.Y(n_4088)
);

INVxp33_ASAP7_75t_L g4089 ( 
.A(n_3613),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3829),
.Y(n_4090)
);

NOR2xp33_ASAP7_75t_L g4091 ( 
.A(n_3463),
.B(n_3004),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_L g4092 ( 
.A(n_3901),
.B(n_2939),
.Y(n_4092)
);

XOR2xp5_ASAP7_75t_L g4093 ( 
.A(n_3799),
.B(n_2152),
.Y(n_4093)
);

XOR2xp5_ASAP7_75t_L g4094 ( 
.A(n_3811),
.B(n_2152),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3835),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3835),
.Y(n_4096)
);

AOI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_3395),
.A2(n_3034),
.B(n_3310),
.Y(n_4097)
);

XOR2xp5_ASAP7_75t_L g4098 ( 
.A(n_3830),
.B(n_2161),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_3776),
.B(n_3234),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3841),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3841),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3844),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3781),
.B(n_2739),
.Y(n_4103)
);

XNOR2x2_ASAP7_75t_L g4104 ( 
.A(n_3834),
.B(n_2654),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3844),
.Y(n_4105)
);

INVx1_ASAP7_75t_L g4106 ( 
.A(n_3537),
.Y(n_4106)
);

XOR2xp5_ASAP7_75t_L g4107 ( 
.A(n_3868),
.B(n_2161),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3901),
.B(n_2940),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3537),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3542),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3542),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3545),
.Y(n_4112)
);

XOR2xp5_ASAP7_75t_L g4113 ( 
.A(n_3937),
.B(n_2163),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3545),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_3378),
.B(n_2739),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3547),
.Y(n_4116)
);

XOR2xp5_ASAP7_75t_L g4117 ( 
.A(n_3402),
.B(n_2163),
.Y(n_4117)
);

INVxp67_ASAP7_75t_SL g4118 ( 
.A(n_3795),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3547),
.Y(n_4119)
);

OR2x6_ASAP7_75t_L g4120 ( 
.A(n_3595),
.B(n_2817),
.Y(n_4120)
);

CKINVDCx5p33_ASAP7_75t_R g4121 ( 
.A(n_3749),
.Y(n_4121)
);

NAND2x1p5_ASAP7_75t_L g4122 ( 
.A(n_3470),
.B(n_3324),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_3378),
.B(n_2512),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3556),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3556),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3572),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3894),
.B(n_2837),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3572),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_3894),
.B(n_2837),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3577),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3577),
.Y(n_4131)
);

INVx1_ASAP7_75t_L g4132 ( 
.A(n_3579),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3579),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3581),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3463),
.B(n_2860),
.Y(n_4135)
);

INVx2_ASAP7_75t_SL g4136 ( 
.A(n_3517),
.Y(n_4136)
);

OAI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_3756),
.A2(n_3274),
.B(n_3310),
.Y(n_4137)
);

XOR2xp5_ASAP7_75t_L g4138 ( 
.A(n_3718),
.B(n_2167),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3581),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3583),
.Y(n_4140)
);

NOR2xp33_ASAP7_75t_L g4141 ( 
.A(n_3469),
.B(n_3365),
.Y(n_4141)
);

NOR2xp33_ASAP7_75t_L g4142 ( 
.A(n_3469),
.B(n_2861),
.Y(n_4142)
);

INVx2_ASAP7_75t_SL g4143 ( 
.A(n_3517),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3583),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3592),
.Y(n_4145)
);

BUFx3_ASAP7_75t_L g4146 ( 
.A(n_3749),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_3762),
.Y(n_4147)
);

BUFx2_ASAP7_75t_L g4148 ( 
.A(n_3417),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3592),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_3901),
.B(n_2946),
.Y(n_4150)
);

NAND2xp5_ASAP7_75t_L g4151 ( 
.A(n_3498),
.B(n_2956),
.Y(n_4151)
);

XOR2x2_ASAP7_75t_L g4152 ( 
.A(n_3747),
.B(n_2633),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3502),
.B(n_2860),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3594),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_3594),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3603),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_3603),
.Y(n_4157)
);

INVxp67_ASAP7_75t_SL g4158 ( 
.A(n_3485),
.Y(n_4158)
);

AND2x2_ASAP7_75t_L g4159 ( 
.A(n_3502),
.B(n_2862),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_3568),
.B(n_2958),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3606),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3606),
.Y(n_4162)
);

XOR2xp5_ASAP7_75t_L g4163 ( 
.A(n_3409),
.B(n_2167),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3762),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3614),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3614),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3619),
.Y(n_4167)
);

AND2x2_ASAP7_75t_SL g4168 ( 
.A(n_3597),
.B(n_2912),
.Y(n_4168)
);

NOR2xp33_ASAP7_75t_L g4169 ( 
.A(n_3695),
.B(n_2867),
.Y(n_4169)
);

BUFx6f_ASAP7_75t_L g4170 ( 
.A(n_3769),
.Y(n_4170)
);

INVx2_ASAP7_75t_L g4171 ( 
.A(n_3765),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_3619),
.Y(n_4172)
);

NOR2xp33_ASAP7_75t_SL g4173 ( 
.A(n_3664),
.B(n_2817),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3626),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_3765),
.Y(n_4175)
);

INVx2_ASAP7_75t_SL g4176 ( 
.A(n_3911),
.Y(n_4176)
);

XOR2xp5_ASAP7_75t_L g4177 ( 
.A(n_3914),
.B(n_2180),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3626),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_3770),
.Y(n_4179)
);

INVxp67_ASAP7_75t_SL g4180 ( 
.A(n_3863),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3628),
.Y(n_4181)
);

NOR2x1p5_ASAP7_75t_L g4182 ( 
.A(n_3757),
.B(n_2470),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3628),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_3541),
.B(n_2870),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_SL g4185 ( 
.A(n_3664),
.B(n_2180),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3560),
.B(n_2962),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3635),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3635),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_3587),
.B(n_2872),
.Y(n_4189)
);

INVxp67_ASAP7_75t_SL g4190 ( 
.A(n_3740),
.Y(n_4190)
);

HB1xp67_ASAP7_75t_L g4191 ( 
.A(n_3754),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_3647),
.Y(n_4192)
);

OR2x2_ASAP7_75t_L g4193 ( 
.A(n_3612),
.B(n_2873),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3647),
.Y(n_4194)
);

BUFx3_ASAP7_75t_L g4195 ( 
.A(n_3757),
.Y(n_4195)
);

INVxp67_ASAP7_75t_SL g4196 ( 
.A(n_3787),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_3650),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3650),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_L g4199 ( 
.A(n_3623),
.B(n_3074),
.Y(n_4199)
);

CKINVDCx5p33_ASAP7_75t_R g4200 ( 
.A(n_3460),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_3823),
.B(n_3075),
.Y(n_4201)
);

CKINVDCx5p33_ASAP7_75t_R g4202 ( 
.A(n_3460),
.Y(n_4202)
);

XOR2xp5_ASAP7_75t_L g4203 ( 
.A(n_3374),
.B(n_2185),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3652),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3652),
.Y(n_4205)
);

BUFx2_ASAP7_75t_L g4206 ( 
.A(n_3748),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3653),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_3653),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_3655),
.Y(n_4209)
);

OAI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_3756),
.A2(n_3274),
.B(n_3328),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3655),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_3826),
.B(n_3085),
.Y(n_4212)
);

NOR2xp33_ASAP7_75t_L g4213 ( 
.A(n_3415),
.B(n_3931),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3661),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_3541),
.B(n_2790),
.Y(n_4215)
);

CKINVDCx5p33_ASAP7_75t_R g4216 ( 
.A(n_3460),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3661),
.Y(n_4217)
);

NAND2xp33_ASAP7_75t_R g4218 ( 
.A(n_3639),
.B(n_2519),
.Y(n_4218)
);

NOR2xp33_ASAP7_75t_L g4219 ( 
.A(n_3430),
.B(n_3107),
.Y(n_4219)
);

BUFx3_ASAP7_75t_L g4220 ( 
.A(n_3460),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3667),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3667),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3668),
.Y(n_4223)
);

BUFx2_ASAP7_75t_L g4224 ( 
.A(n_3748),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_3439),
.B(n_2811),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_3567),
.B(n_2612),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_L g4227 ( 
.A(n_3751),
.B(n_3119),
.Y(n_4227)
);

XOR2xp5_ASAP7_75t_L g4228 ( 
.A(n_3750),
.B(n_2185),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3668),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_3770),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3669),
.B(n_3058),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_3376),
.B(n_3125),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_3773),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3669),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_3773),
.Y(n_4235)
);

INVxp33_ASAP7_75t_L g4236 ( 
.A(n_3536),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3672),
.B(n_3068),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_3775),
.Y(n_4238)
);

XOR2xp5_ASAP7_75t_L g4239 ( 
.A(n_3750),
.B(n_2191),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_3591),
.B(n_2612),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3672),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3596),
.B(n_2612),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_3675),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_3561),
.B(n_3324),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_3675),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_3683),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_3602),
.B(n_3551),
.Y(n_4247)
);

NOR2xp33_ASAP7_75t_L g4248 ( 
.A(n_3376),
.B(n_3131),
.Y(n_4248)
);

INVx1_ASAP7_75t_SL g4249 ( 
.A(n_3612),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_3683),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_3687),
.Y(n_4251)
);

NOR2xp33_ASAP7_75t_L g4252 ( 
.A(n_3376),
.B(n_3139),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3687),
.Y(n_4253)
);

AND2x2_ASAP7_75t_L g4254 ( 
.A(n_3553),
.B(n_3376),
.Y(n_4254)
);

INVx2_ASAP7_75t_SL g4255 ( 
.A(n_3911),
.Y(n_4255)
);

CKINVDCx20_ASAP7_75t_R g4256 ( 
.A(n_3855),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_3429),
.B(n_2591),
.Y(n_4257)
);

NOR2xp33_ASAP7_75t_L g4258 ( 
.A(n_3662),
.B(n_3220),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3689),
.Y(n_4259)
);

AND2x6_ASAP7_75t_L g4260 ( 
.A(n_3611),
.B(n_3705),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_3610),
.B(n_1898),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_3689),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_3696),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_3696),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3698),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_3698),
.B(n_3076),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3701),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_3701),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3711),
.Y(n_4269)
);

INVx2_ASAP7_75t_L g4270 ( 
.A(n_3775),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_3779),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_3779),
.Y(n_4272)
);

XOR2xp5_ASAP7_75t_L g4273 ( 
.A(n_3690),
.B(n_2191),
.Y(n_4273)
);

AOI21xp5_ASAP7_75t_L g4274 ( 
.A1(n_3772),
.A2(n_2927),
.B(n_2904),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_3711),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3719),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_3719),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_3720),
.Y(n_4278)
);

NAND2xp33_ASAP7_75t_R g4279 ( 
.A(n_3639),
.B(n_2519),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_3720),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_3721),
.Y(n_4281)
);

AND2x4_ASAP7_75t_L g4282 ( 
.A(n_3917),
.B(n_3185),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3721),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_3726),
.Y(n_4284)
);

CKINVDCx20_ASAP7_75t_R g4285 ( 
.A(n_3514),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_3726),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_3791),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_SL g4288 ( 
.A(n_3664),
.B(n_2195),
.Y(n_4288)
);

AND2x2_ASAP7_75t_L g4289 ( 
.A(n_3663),
.B(n_1908),
.Y(n_4289)
);

CKINVDCx20_ASAP7_75t_R g4290 ( 
.A(n_3514),
.Y(n_4290)
);

BUFx6f_ASAP7_75t_L g4291 ( 
.A(n_3833),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_3733),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_3733),
.Y(n_4293)
);

BUFx5_ASAP7_75t_L g4294 ( 
.A(n_3576),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3734),
.B(n_3077),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_3734),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_3684),
.B(n_3792),
.Y(n_4297)
);

INVx2_ASAP7_75t_L g4298 ( 
.A(n_3791),
.Y(n_4298)
);

OR2x2_ASAP7_75t_L g4299 ( 
.A(n_3644),
.B(n_3870),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_3735),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_3735),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_3793),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_3793),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3752),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_3752),
.Y(n_4305)
);

INVx1_ASAP7_75t_L g4306 ( 
.A(n_3753),
.Y(n_4306)
);

OAI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_3772),
.A2(n_3328),
.B(n_3039),
.Y(n_4307)
);

XOR2xp5_ASAP7_75t_L g4308 ( 
.A(n_3617),
.B(n_2195),
.Y(n_4308)
);

INVx3_ASAP7_75t_L g4309 ( 
.A(n_3470),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_3753),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_3763),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_3763),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3767),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_3806),
.B(n_1908),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3767),
.Y(n_4315)
);

CKINVDCx20_ASAP7_75t_R g4316 ( 
.A(n_3514),
.Y(n_4316)
);

XNOR2xp5_ASAP7_75t_L g4317 ( 
.A(n_3812),
.B(n_2198),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_3794),
.Y(n_4318)
);

INVxp67_ASAP7_75t_L g4319 ( 
.A(n_3825),
.Y(n_4319)
);

OR2x2_ASAP7_75t_L g4320 ( 
.A(n_3644),
.B(n_2957),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3771),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_3890),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3771),
.Y(n_4323)
);

XOR2xp5_ASAP7_75t_L g4324 ( 
.A(n_3380),
.B(n_2198),
.Y(n_4324)
);

NAND2xp33_ASAP7_75t_R g4325 ( 
.A(n_3639),
.B(n_2633),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_3778),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_3778),
.Y(n_4327)
);

BUFx3_ASAP7_75t_L g4328 ( 
.A(n_3514),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3784),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3784),
.Y(n_4330)
);

NOR2xp33_ASAP7_75t_L g4331 ( 
.A(n_3853),
.B(n_3244),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_3566),
.B(n_1909),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_3788),
.Y(n_4333)
);

AND2x2_ASAP7_75t_L g4334 ( 
.A(n_3566),
.B(n_1909),
.Y(n_4334)
);

CKINVDCx5p33_ASAP7_75t_R g4335 ( 
.A(n_3831),
.Y(n_4335)
);

NOR2xp33_ASAP7_75t_L g4336 ( 
.A(n_3875),
.B(n_3325),
.Y(n_4336)
);

INVx2_ASAP7_75t_L g4337 ( 
.A(n_3794),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3788),
.Y(n_4338)
);

OR2x6_ASAP7_75t_L g4339 ( 
.A(n_3595),
.B(n_3715),
.Y(n_4339)
);

XOR2xp5_ASAP7_75t_L g4340 ( 
.A(n_3544),
.B(n_2236),
.Y(n_4340)
);

AND2x4_ASAP7_75t_L g4341 ( 
.A(n_3608),
.B(n_3186),
.Y(n_4341)
);

XOR2xp5_ASAP7_75t_L g4342 ( 
.A(n_3870),
.B(n_2236),
.Y(n_4342)
);

CKINVDCx20_ASAP7_75t_R g4343 ( 
.A(n_3855),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3789),
.Y(n_4344)
);

INVx1_ASAP7_75t_L g4345 ( 
.A(n_3789),
.Y(n_4345)
);

INVx2_ASAP7_75t_L g4346 ( 
.A(n_3800),
.Y(n_4346)
);

INVx1_ASAP7_75t_L g4347 ( 
.A(n_3797),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3797),
.B(n_3078),
.Y(n_4348)
);

AND2x6_ASAP7_75t_L g4349 ( 
.A(n_3611),
.B(n_2941),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_3809),
.B(n_3080),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_3800),
.Y(n_4351)
);

XNOR2x2_ASAP7_75t_L g4352 ( 
.A(n_3562),
.B(n_2842),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_3809),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_SL g4354 ( 
.A(n_3561),
.B(n_3598),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3813),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3813),
.Y(n_4356)
);

NOR2xp33_ASAP7_75t_L g4357 ( 
.A(n_3712),
.B(n_3349),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3817),
.Y(n_4358)
);

AOI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_3691),
.A2(n_2971),
.B(n_2932),
.Y(n_4359)
);

XOR2xp5_ASAP7_75t_L g4360 ( 
.A(n_3427),
.B(n_2238),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_3817),
.B(n_3082),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_3822),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_3608),
.B(n_3187),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_3822),
.Y(n_4364)
);

XOR2xp5_ASAP7_75t_L g4365 ( 
.A(n_3465),
.B(n_2238),
.Y(n_4365)
);

NOR2xp33_ASAP7_75t_L g4366 ( 
.A(n_3712),
.B(n_3356),
.Y(n_4366)
);

XOR2xp5_ASAP7_75t_L g4367 ( 
.A(n_3470),
.B(n_2251),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3828),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3828),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_3436),
.B(n_3093),
.Y(n_4370)
);

AND2x2_ASAP7_75t_L g4371 ( 
.A(n_3936),
.B(n_3639),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_3849),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3849),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_3852),
.Y(n_4374)
);

XNOR2x2_ASAP7_75t_L g4375 ( 
.A(n_3570),
.B(n_849),
.Y(n_4375)
);

CKINVDCx20_ASAP7_75t_R g4376 ( 
.A(n_3419),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_3852),
.Y(n_4377)
);

INVx2_ASAP7_75t_SL g4378 ( 
.A(n_3812),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_3884),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_3884),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_3892),
.Y(n_4381)
);

HB1xp67_ASAP7_75t_L g4382 ( 
.A(n_3869),
.Y(n_4382)
);

INVx2_ASAP7_75t_SL g4383 ( 
.A(n_3867),
.Y(n_4383)
);

XOR2xp5_ASAP7_75t_L g4384 ( 
.A(n_3470),
.B(n_2251),
.Y(n_4384)
);

INVxp67_ASAP7_75t_SL g4385 ( 
.A(n_3833),
.Y(n_4385)
);

AND2x2_ASAP7_75t_L g4386 ( 
.A(n_3639),
.B(n_1912),
.Y(n_4386)
);

BUFx6f_ASAP7_75t_SL g4387 ( 
.A(n_3608),
.Y(n_4387)
);

XOR2xp5_ASAP7_75t_L g4388 ( 
.A(n_3656),
.B(n_2252),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_3858),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_3867),
.B(n_1912),
.Y(n_4390)
);

XNOR2xp5_ASAP7_75t_L g4391 ( 
.A(n_3608),
.B(n_2252),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_3858),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_3864),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_3864),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_3882),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_3920),
.B(n_1913),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_3831),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_3882),
.Y(n_4398)
);

BUFx6f_ASAP7_75t_L g4399 ( 
.A(n_3833),
.Y(n_4399)
);

XOR2xp5_ASAP7_75t_L g4400 ( 
.A(n_3903),
.B(n_2258),
.Y(n_4400)
);

CKINVDCx16_ASAP7_75t_R g4401 ( 
.A(n_3831),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_3883),
.Y(n_4402)
);

XNOR2xp5_ASAP7_75t_L g4403 ( 
.A(n_3608),
.B(n_2258),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_3883),
.Y(n_4404)
);

BUFx2_ASAP7_75t_L g4405 ( 
.A(n_3458),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_3888),
.Y(n_4406)
);

OR2x2_ASAP7_75t_L g4407 ( 
.A(n_3910),
.B(n_2957),
.Y(n_4407)
);

OR2x6_ASAP7_75t_L g4408 ( 
.A(n_3595),
.B(n_3366),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_3624),
.B(n_3098),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_3888),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_3893),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_3893),
.Y(n_4412)
);

NOR2xp33_ASAP7_75t_L g4413 ( 
.A(n_3462),
.B(n_2566),
.Y(n_4413)
);

NOR2xp33_ASAP7_75t_L g4414 ( 
.A(n_3755),
.B(n_2566),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_3896),
.Y(n_4415)
);

AND2x2_ASAP7_75t_L g4416 ( 
.A(n_3744),
.B(n_1917),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_3896),
.Y(n_4417)
);

BUFx2_ASAP7_75t_L g4418 ( 
.A(n_3458),
.Y(n_4418)
);

NOR2xp33_ASAP7_75t_L g4419 ( 
.A(n_3786),
.B(n_3790),
.Y(n_4419)
);

XOR2xp5_ASAP7_75t_L g4420 ( 
.A(n_3903),
.B(n_2260),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3900),
.Y(n_4421)
);

CKINVDCx20_ASAP7_75t_R g4422 ( 
.A(n_3458),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_3744),
.B(n_1917),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_3900),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_3902),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_3902),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_3905),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_L g4428 ( 
.A(n_3631),
.B(n_3102),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_3905),
.Y(n_4429)
);

CKINVDCx16_ASAP7_75t_R g4430 ( 
.A(n_3845),
.Y(n_4430)
);

XOR2xp5_ASAP7_75t_L g4431 ( 
.A(n_3390),
.B(n_2260),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_3906),
.Y(n_4432)
);

INVxp33_ASAP7_75t_SL g4433 ( 
.A(n_3438),
.Y(n_4433)
);

BUFx8_ASAP7_75t_L g4434 ( 
.A(n_3845),
.Y(n_4434)
);

CKINVDCx5p33_ASAP7_75t_R g4435 ( 
.A(n_3845),
.Y(n_4435)
);

XOR2xp5_ASAP7_75t_L g4436 ( 
.A(n_3785),
.B(n_2265),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_3906),
.Y(n_4437)
);

BUFx6f_ASAP7_75t_L g4438 ( 
.A(n_3833),
.Y(n_4438)
);

OAI21xp5_ASAP7_75t_L g4439 ( 
.A1(n_3397),
.A2(n_3039),
.B(n_3037),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_3907),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_3744),
.B(n_1930),
.Y(n_4441)
);

AOI21x1_ASAP7_75t_L g4442 ( 
.A1(n_3924),
.A2(n_3330),
.B(n_2948),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_3638),
.B(n_3106),
.Y(n_4443)
);

XNOR2xp5_ASAP7_75t_L g4444 ( 
.A(n_3880),
.B(n_2265),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_3907),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_3946),
.Y(n_4446)
);

OR2x2_ASAP7_75t_L g4447 ( 
.A(n_4299),
.B(n_3593),
.Y(n_4447)
);

INVx2_ASAP7_75t_L g4448 ( 
.A(n_3948),
.Y(n_4448)
);

OAI221xp5_ASAP7_75t_L g4449 ( 
.A1(n_4056),
.A2(n_3351),
.B1(n_3280),
.B2(n_3630),
.C(n_3625),
.Y(n_4449)
);

O2A1O1Ixp33_ASAP7_75t_L g4450 ( 
.A1(n_4049),
.A2(n_3682),
.B(n_3708),
.C(n_3702),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_3970),
.Y(n_4451)
);

INVx2_ASAP7_75t_L g4452 ( 
.A(n_4001),
.Y(n_4452)
);

AOI22xp33_ASAP7_75t_L g4453 ( 
.A1(n_4076),
.A2(n_3785),
.B1(n_3654),
.B2(n_3515),
.Y(n_4453)
);

NOR2xp33_ASAP7_75t_L g4454 ( 
.A(n_3966),
.B(n_2268),
.Y(n_4454)
);

AOI22xp33_ASAP7_75t_L g4455 ( 
.A1(n_3954),
.A2(n_3500),
.B1(n_3651),
.B2(n_3497),
.Y(n_4455)
);

INVxp33_ASAP7_75t_L g4456 ( 
.A(n_4273),
.Y(n_4456)
);

NOR2xp33_ASAP7_75t_L g4457 ( 
.A(n_3966),
.B(n_2268),
.Y(n_4457)
);

INVxp67_ASAP7_75t_L g4458 ( 
.A(n_4148),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4049),
.B(n_3550),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_SL g4460 ( 
.A(n_4247),
.B(n_3744),
.Y(n_4460)
);

INVx2_ASAP7_75t_SL g4461 ( 
.A(n_4434),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4056),
.B(n_3552),
.Y(n_4462)
);

NAND2xp5_ASAP7_75t_L g4463 ( 
.A(n_3980),
.B(n_2825),
.Y(n_4463)
);

AOI221xp5_ASAP7_75t_L g4464 ( 
.A1(n_4081),
.A2(n_1288),
.B1(n_980),
.B2(n_1002),
.C(n_978),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_3980),
.B(n_2825),
.Y(n_4465)
);

INVx3_ASAP7_75t_L g4466 ( 
.A(n_3977),
.Y(n_4466)
);

INVx1_ASAP7_75t_SL g4467 ( 
.A(n_4249),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_3988),
.B(n_2825),
.Y(n_4468)
);

INVx2_ASAP7_75t_SL g4469 ( 
.A(n_4434),
.Y(n_4469)
);

AOI22xp33_ASAP7_75t_L g4470 ( 
.A1(n_4030),
.A2(n_3486),
.B1(n_3731),
.B2(n_3108),
.Y(n_4470)
);

OAI21xp5_ASAP7_75t_L g4471 ( 
.A1(n_4081),
.A2(n_3442),
.B(n_3440),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_SL g4472 ( 
.A(n_4254),
.B(n_3891),
.Y(n_4472)
);

INVxp67_ASAP7_75t_L g4473 ( 
.A(n_3990),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_SL g4474 ( 
.A(n_4213),
.B(n_3891),
.Y(n_4474)
);

INVx2_ASAP7_75t_SL g4475 ( 
.A(n_3967),
.Y(n_4475)
);

NOR2xp33_ASAP7_75t_L g4476 ( 
.A(n_3951),
.B(n_3816),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_4213),
.B(n_3891),
.Y(n_4477)
);

BUFx6f_ASAP7_75t_SL g4478 ( 
.A(n_3978),
.Y(n_4478)
);

INVx2_ASAP7_75t_L g4479 ( 
.A(n_4043),
.Y(n_4479)
);

NOR2xp33_ASAP7_75t_L g4480 ( 
.A(n_4046),
.B(n_2271),
.Y(n_4480)
);

O2A1O1Ixp33_ASAP7_75t_L g4481 ( 
.A1(n_3951),
.A2(n_3554),
.B(n_3601),
.C(n_3798),
.Y(n_4481)
);

NOR2xp33_ASAP7_75t_L g4482 ( 
.A(n_4046),
.B(n_3454),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_4078),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_3988),
.B(n_2434),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4123),
.B(n_2982),
.Y(n_4485)
);

INVx3_ASAP7_75t_L g4486 ( 
.A(n_3977),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_3950),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_L g4488 ( 
.A(n_4089),
.B(n_3820),
.Y(n_4488)
);

AOI22xp5_ASAP7_75t_L g4489 ( 
.A1(n_4212),
.A2(n_2719),
.B1(n_2434),
.B2(n_3782),
.Y(n_4489)
);

NOR2x1_ASAP7_75t_R g4490 ( 
.A(n_4071),
.B(n_2764),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_3995),
.B(n_2434),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_3995),
.B(n_2719),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_L g4493 ( 
.A(n_4089),
.B(n_3821),
.Y(n_4493)
);

NAND3xp33_ASAP7_75t_L g4494 ( 
.A(n_4212),
.B(n_3935),
.C(n_2719),
.Y(n_4494)
);

NAND2xp33_ASAP7_75t_L g4495 ( 
.A(n_4260),
.B(n_3703),
.Y(n_4495)
);

AOI22xp33_ASAP7_75t_L g4496 ( 
.A1(n_4436),
.A2(n_3109),
.B1(n_3116),
.B2(n_3110),
.Y(n_4496)
);

OAI22xp5_ASAP7_75t_L g4497 ( 
.A1(n_4006),
.A2(n_3450),
.B1(n_3741),
.B2(n_3705),
.Y(n_4497)
);

INVx2_ASAP7_75t_SL g4498 ( 
.A(n_3967),
.Y(n_4498)
);

NOR2xp33_ASAP7_75t_L g4499 ( 
.A(n_4006),
.B(n_3836),
.Y(n_4499)
);

NOR2xp33_ASAP7_75t_L g4500 ( 
.A(n_4236),
.B(n_3918),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_3968),
.B(n_1933),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_SL g4502 ( 
.A(n_4087),
.B(n_3891),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4080),
.Y(n_4503)
);

AOI22xp33_ASAP7_75t_L g4504 ( 
.A1(n_4324),
.A2(n_3118),
.B1(n_3126),
.B2(n_3123),
.Y(n_4504)
);

NAND2xp5_ASAP7_75t_L g4505 ( 
.A(n_4040),
.B(n_1933),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_3964),
.Y(n_4506)
);

INVx2_ASAP7_75t_L g4507 ( 
.A(n_4147),
.Y(n_4507)
);

NOR2xp33_ASAP7_75t_L g4508 ( 
.A(n_4236),
.B(n_3918),
.Y(n_4508)
);

NAND2x1p5_ASAP7_75t_L g4509 ( 
.A(n_4168),
.B(n_3918),
.Y(n_4509)
);

NOR2xp33_ASAP7_75t_L g4510 ( 
.A(n_4040),
.B(n_3918),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_SL g4511 ( 
.A(n_4087),
.B(n_3375),
.Y(n_4511)
);

INVx2_ASAP7_75t_SL g4512 ( 
.A(n_3967),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_3990),
.Y(n_4513)
);

NOR3xp33_ASAP7_75t_L g4514 ( 
.A(n_4227),
.B(n_3854),
.C(n_3840),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_SL g4515 ( 
.A(n_4028),
.B(n_3375),
.Y(n_4515)
);

INVx2_ASAP7_75t_L g4516 ( 
.A(n_4164),
.Y(n_4516)
);

O2A1O1Ixp33_ASAP7_75t_L g4517 ( 
.A1(n_4227),
.A2(n_3725),
.B(n_3466),
.C(n_3543),
.Y(n_4517)
);

INVx4_ASAP7_75t_L g4518 ( 
.A(n_3983),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4189),
.B(n_1935),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_SL g4520 ( 
.A(n_4034),
.B(n_3375),
.Y(n_4520)
);

INVxp67_ASAP7_75t_L g4521 ( 
.A(n_4142),
.Y(n_4521)
);

INVx2_ASAP7_75t_L g4522 ( 
.A(n_4171),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_SL g4523 ( 
.A(n_4169),
.B(n_3375),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_4342),
.B(n_3519),
.Y(n_4524)
);

INVx2_ASAP7_75t_L g4525 ( 
.A(n_4175),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_3961),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4372),
.Y(n_4527)
);

OR2x6_ASAP7_75t_L g4528 ( 
.A(n_4339),
.B(n_3595),
.Y(n_4528)
);

NOR2xp67_ASAP7_75t_L g4529 ( 
.A(n_4041),
.B(n_3284),
.Y(n_4529)
);

INVx3_ASAP7_75t_L g4530 ( 
.A(n_4309),
.Y(n_4530)
);

OAI22xp33_ASAP7_75t_L g4531 ( 
.A1(n_4218),
.A2(n_3741),
.B1(n_3856),
.B2(n_3780),
.Y(n_4531)
);

AOI21xp5_ASAP7_75t_L g4532 ( 
.A1(n_4023),
.A2(n_3706),
.B(n_3549),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4189),
.B(n_1935),
.Y(n_4533)
);

BUFx6f_ASAP7_75t_L g4534 ( 
.A(n_3945),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_4179),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4373),
.Y(n_4536)
);

INVx2_ASAP7_75t_L g4537 ( 
.A(n_4230),
.Y(n_4537)
);

NAND2x1_ASAP7_75t_L g4538 ( 
.A(n_4339),
.B(n_3382),
.Y(n_4538)
);

BUFx2_ASAP7_75t_L g4539 ( 
.A(n_3972),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_3953),
.B(n_1939),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4057),
.B(n_2982),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_SL g4542 ( 
.A(n_4169),
.B(n_3375),
.Y(n_4542)
);

BUFx12f_ASAP7_75t_L g4543 ( 
.A(n_4121),
.Y(n_4543)
);

OR2x2_ASAP7_75t_L g4544 ( 
.A(n_4193),
.B(n_3458),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_SL g4545 ( 
.A(n_4336),
.B(n_3381),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4233),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_L g4547 ( 
.A(n_4226),
.B(n_1939),
.Y(n_4547)
);

INVx2_ASAP7_75t_L g4548 ( 
.A(n_4235),
.Y(n_4548)
);

INVx2_ASAP7_75t_SL g4549 ( 
.A(n_3987),
.Y(n_4549)
);

NOR2xp67_ASAP7_75t_L g4550 ( 
.A(n_4378),
.B(n_3286),
.Y(n_4550)
);

OR2x6_ASAP7_75t_L g4551 ( 
.A(n_4339),
.B(n_3715),
.Y(n_4551)
);

NAND3xp33_ASAP7_75t_L g4552 ( 
.A(n_4336),
.B(n_3183),
.C(n_2983),
.Y(n_4552)
);

INVxp67_ASAP7_75t_SL g4553 ( 
.A(n_4190),
.Y(n_4553)
);

NOR2xp67_ASAP7_75t_L g4554 ( 
.A(n_4383),
.B(n_3301),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_4240),
.B(n_4242),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4238),
.Y(n_4556)
);

NOR2xp33_ASAP7_75t_L g4557 ( 
.A(n_4225),
.B(n_3449),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4374),
.Y(n_4558)
);

AND2x4_ASAP7_75t_L g4559 ( 
.A(n_3945),
.B(n_3458),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4396),
.B(n_1940),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_3989),
.B(n_1940),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_3989),
.B(n_1946),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4270),
.Y(n_4563)
);

AOI22xp5_ASAP7_75t_L g4564 ( 
.A1(n_4340),
.A2(n_2782),
.B1(n_2794),
.B2(n_2764),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4377),
.Y(n_4565)
);

INVxp33_ASAP7_75t_SL g4566 ( 
.A(n_3974),
.Y(n_4566)
);

AOI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_4104),
.A2(n_4400),
.B1(n_4420),
.B2(n_4203),
.Y(n_4567)
);

AOI22xp33_ASAP7_75t_L g4568 ( 
.A1(n_4163),
.A2(n_3162),
.B1(n_3168),
.B2(n_3163),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_SL g4569 ( 
.A(n_4433),
.B(n_4168),
.Y(n_4569)
);

AOI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4138),
.A2(n_2794),
.B1(n_2782),
.B2(n_3183),
.Y(n_4570)
);

INVx2_ASAP7_75t_L g4571 ( 
.A(n_4271),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4272),
.Y(n_4572)
);

INVx3_ASAP7_75t_L g4573 ( 
.A(n_4309),
.Y(n_4573)
);

NAND2xp5_ASAP7_75t_L g4574 ( 
.A(n_4199),
.B(n_1946),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4389),
.Y(n_4575)
);

INVx8_ASAP7_75t_L g4576 ( 
.A(n_4003),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4199),
.B(n_1951),
.Y(n_4577)
);

AOI22xp33_ASAP7_75t_L g4578 ( 
.A1(n_4388),
.A2(n_3766),
.B1(n_3897),
.B2(n_3837),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_SL g4579 ( 
.A(n_4219),
.B(n_3381),
.Y(n_4579)
);

INVx3_ASAP7_75t_L g4580 ( 
.A(n_3949),
.Y(n_4580)
);

INVx8_ASAP7_75t_L g4581 ( 
.A(n_4003),
.Y(n_4581)
);

BUFx6f_ASAP7_75t_L g4582 ( 
.A(n_3962),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4083),
.B(n_1951),
.Y(n_4583)
);

NOR2xp67_ASAP7_75t_SL g4584 ( 
.A(n_4146),
.B(n_2693),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4392),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4319),
.B(n_1952),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4319),
.B(n_1952),
.Y(n_4587)
);

A2O1A1Ixp33_ASAP7_75t_L g4588 ( 
.A1(n_4357),
.A2(n_3856),
.B(n_3780),
.C(n_3660),
.Y(n_4588)
);

NAND2xp33_ASAP7_75t_L g4589 ( 
.A(n_4260),
.B(n_3703),
.Y(n_4589)
);

INVx1_ASAP7_75t_L g4590 ( 
.A(n_4393),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_3973),
.B(n_1953),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4394),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_SL g4593 ( 
.A(n_4219),
.B(n_3381),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4395),
.Y(n_4594)
);

AND2x6_ASAP7_75t_SL g4595 ( 
.A(n_4142),
.B(n_4261),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_3993),
.B(n_1953),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4398),
.Y(n_4597)
);

INVxp67_ASAP7_75t_L g4598 ( 
.A(n_4016),
.Y(n_4598)
);

NOR2xp33_ASAP7_75t_L g4599 ( 
.A(n_4018),
.B(n_3461),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_3999),
.B(n_1954),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4287),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4027),
.B(n_1954),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_SL g4603 ( 
.A(n_4341),
.B(n_3381),
.Y(n_4603)
);

AOI22xp33_ASAP7_75t_L g4604 ( 
.A1(n_4431),
.A2(n_3766),
.B1(n_3897),
.B2(n_3837),
.Y(n_4604)
);

HB1xp67_ASAP7_75t_L g4605 ( 
.A(n_4018),
.Y(n_4605)
);

NOR2xp33_ASAP7_75t_L g4606 ( 
.A(n_4320),
.B(n_2693),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4033),
.B(n_1955),
.Y(n_4607)
);

NOR2xp33_ASAP7_75t_L g4608 ( 
.A(n_3962),
.B(n_3899),
.Y(n_4608)
);

NAND2xp33_ASAP7_75t_L g4609 ( 
.A(n_4260),
.B(n_3727),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4402),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4039),
.B(n_2982),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4404),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4159),
.B(n_1963),
.Y(n_4613)
);

AO22x1_ASAP7_75t_L g4614 ( 
.A1(n_4335),
.A2(n_2794),
.B1(n_2782),
.B2(n_3183),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4406),
.Y(n_4615)
);

NOR2xp33_ASAP7_75t_L g4616 ( 
.A(n_4201),
.B(n_3909),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4184),
.B(n_1963),
.Y(n_4617)
);

INVxp67_ASAP7_75t_L g4618 ( 
.A(n_4016),
.Y(n_4618)
);

NOR2xp67_ASAP7_75t_L g4619 ( 
.A(n_4176),
.B(n_2999),
.Y(n_4619)
);

AND2x2_ASAP7_75t_SL g4620 ( 
.A(n_4173),
.B(n_3597),
.Y(n_4620)
);

NOR2xp33_ASAP7_75t_L g4621 ( 
.A(n_4000),
.B(n_3362),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4215),
.B(n_4257),
.Y(n_4622)
);

NAND2xp5_ASAP7_75t_SL g4623 ( 
.A(n_4341),
.B(n_3381),
.Y(n_4623)
);

A2O1A1Ixp33_ASAP7_75t_L g4624 ( 
.A1(n_4357),
.A2(n_4366),
.B(n_4201),
.C(n_4331),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_4410),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4297),
.B(n_1967),
.Y(n_4626)
);

INVx2_ASAP7_75t_SL g4627 ( 
.A(n_4255),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_L g4628 ( 
.A(n_3986),
.B(n_1968),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_3986),
.B(n_1968),
.Y(n_4629)
);

AND2x6_ASAP7_75t_L g4630 ( 
.A(n_4363),
.B(n_3576),
.Y(n_4630)
);

NOR2xp33_ASAP7_75t_L g4631 ( 
.A(n_4010),
.B(n_3362),
.Y(n_4631)
);

AOI22xp5_ASAP7_75t_L g4632 ( 
.A1(n_4218),
.A2(n_3362),
.B1(n_1978),
.B2(n_1979),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_SL g4633 ( 
.A(n_4363),
.B(n_3424),
.Y(n_4633)
);

INVx1_ASAP7_75t_L g4634 ( 
.A(n_4411),
.Y(n_4634)
);

NOR2xp33_ASAP7_75t_L g4635 ( 
.A(n_4228),
.B(n_1971),
.Y(n_4635)
);

AND2x6_ASAP7_75t_SL g4636 ( 
.A(n_4390),
.B(n_1378),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4032),
.B(n_1971),
.Y(n_4637)
);

NOR2xp67_ASAP7_75t_L g4638 ( 
.A(n_4045),
.B(n_2999),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4032),
.B(n_1979),
.Y(n_4639)
);

OAI21xp5_ASAP7_75t_L g4640 ( 
.A1(n_4258),
.A2(n_3510),
.B(n_3717),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_4289),
.B(n_1996),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4412),
.Y(n_4642)
);

NOR2xp33_ASAP7_75t_L g4643 ( 
.A(n_4239),
.B(n_1996),
.Y(n_4643)
);

AOI21xp5_ASAP7_75t_L g4644 ( 
.A1(n_4023),
.A2(n_3549),
.B(n_3533),
.Y(n_4644)
);

NOR3xp33_ASAP7_75t_L g4645 ( 
.A(n_4366),
.B(n_4091),
.C(n_4258),
.Y(n_4645)
);

AND2x2_ASAP7_75t_L g4646 ( 
.A(n_4153),
.B(n_2999),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4415),
.Y(n_4647)
);

NOR2xp33_ASAP7_75t_L g4648 ( 
.A(n_3956),
.B(n_1997),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4314),
.B(n_1997),
.Y(n_4649)
);

NOR2xp33_ASAP7_75t_L g4650 ( 
.A(n_4079),
.B(n_3929),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4417),
.Y(n_4651)
);

INVx2_ASAP7_75t_L g4652 ( 
.A(n_4298),
.Y(n_4652)
);

NAND3xp33_ASAP7_75t_L g4653 ( 
.A(n_4331),
.B(n_3002),
.C(n_3467),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4302),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4136),
.B(n_1999),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4143),
.B(n_1999),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4303),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4421),
.Y(n_4658)
);

AND2x2_ASAP7_75t_L g4659 ( 
.A(n_4115),
.B(n_4127),
.Y(n_4659)
);

NOR2xp33_ASAP7_75t_R g4660 ( 
.A(n_4031),
.B(n_3400),
.Y(n_4660)
);

NAND2xp5_ASAP7_75t_SL g4661 ( 
.A(n_4232),
.B(n_3424),
.Y(n_4661)
);

NAND2xp5_ASAP7_75t_L g4662 ( 
.A(n_4186),
.B(n_3189),
.Y(n_4662)
);

AOI22xp5_ASAP7_75t_L g4663 ( 
.A1(n_4279),
.A2(n_3410),
.B1(n_3406),
.B2(n_3400),
.Y(n_4663)
);

INVx2_ASAP7_75t_SL g4664 ( 
.A(n_4195),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4186),
.B(n_3192),
.Y(n_4665)
);

INVx2_ASAP7_75t_L g4666 ( 
.A(n_4318),
.Y(n_4666)
);

AOI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_4097),
.A2(n_3549),
.B(n_3533),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4424),
.Y(n_4668)
);

NOR2xp67_ASAP7_75t_L g4669 ( 
.A(n_4391),
.B(n_3040),
.Y(n_4669)
);

BUFx6f_ASAP7_75t_L g4670 ( 
.A(n_4013),
.Y(n_4670)
);

OAI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4091),
.A2(n_3399),
.B1(n_3382),
.B2(n_3597),
.Y(n_4671)
);

NAND2xp5_ASAP7_75t_L g4672 ( 
.A(n_4191),
.B(n_3199),
.Y(n_4672)
);

INVx2_ASAP7_75t_L g4673 ( 
.A(n_4337),
.Y(n_4673)
);

NOR2xp33_ASAP7_75t_L g4674 ( 
.A(n_4103),
.B(n_3040),
.Y(n_4674)
);

AND2x4_ASAP7_75t_SL g4675 ( 
.A(n_4003),
.B(n_3382),
.Y(n_4675)
);

INVxp67_ASAP7_75t_L g4676 ( 
.A(n_4322),
.Y(n_4676)
);

AND2x2_ASAP7_75t_L g4677 ( 
.A(n_4129),
.B(n_3040),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_L g4678 ( 
.A(n_4191),
.B(n_3204),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4346),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4425),
.Y(n_4680)
);

CKINVDCx5p33_ASAP7_75t_R g4681 ( 
.A(n_3959),
.Y(n_4681)
);

INVx4_ASAP7_75t_L g4682 ( 
.A(n_4120),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_SL g4683 ( 
.A(n_4232),
.B(n_3424),
.Y(n_4683)
);

INVx1_ASAP7_75t_L g4684 ( 
.A(n_4426),
.Y(n_4684)
);

AOI22xp5_ASAP7_75t_L g4685 ( 
.A1(n_4279),
.A2(n_3837),
.B1(n_3727),
.B2(n_3399),
.Y(n_4685)
);

AOI22xp33_ASAP7_75t_L g4686 ( 
.A1(n_4360),
.A2(n_3766),
.B1(n_3897),
.B2(n_3837),
.Y(n_4686)
);

INVx1_ASAP7_75t_L g4687 ( 
.A(n_4427),
.Y(n_4687)
);

NOR2x1p5_ASAP7_75t_L g4688 ( 
.A(n_4200),
.B(n_3492),
.Y(n_4688)
);

INVx3_ASAP7_75t_L g4689 ( 
.A(n_3949),
.Y(n_4689)
);

INVx5_ASAP7_75t_L g4690 ( 
.A(n_4120),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_SL g4691 ( 
.A(n_4248),
.B(n_4252),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4429),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_SL g4693 ( 
.A(n_4248),
.B(n_3424),
.Y(n_4693)
);

INVx2_ASAP7_75t_L g4694 ( 
.A(n_4351),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4332),
.B(n_3209),
.Y(n_4695)
);

INVx2_ASAP7_75t_L g4696 ( 
.A(n_4379),
.Y(n_4696)
);

INVx2_ASAP7_75t_L g4697 ( 
.A(n_4380),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4432),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_4029),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_4334),
.B(n_3213),
.Y(n_4700)
);

CKINVDCx5p33_ASAP7_75t_R g4701 ( 
.A(n_4029),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4158),
.B(n_3216),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4437),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4440),
.Y(n_4704)
);

CKINVDCx20_ASAP7_75t_R g4705 ( 
.A(n_4026),
.Y(n_4705)
);

NOR2xp33_ASAP7_75t_L g4706 ( 
.A(n_4117),
.B(n_3474),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4158),
.B(n_3218),
.Y(n_4707)
);

INVx2_ASAP7_75t_L g4708 ( 
.A(n_4381),
.Y(n_4708)
);

AOI22xp33_ASAP7_75t_L g4709 ( 
.A1(n_4365),
.A2(n_3837),
.B1(n_3457),
.B2(n_2741),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_SL g4710 ( 
.A(n_4252),
.B(n_3965),
.Y(n_4710)
);

NAND2xp5_ASAP7_75t_L g4711 ( 
.A(n_4180),
.B(n_4160),
.Y(n_4711)
);

NOR2xp33_ASAP7_75t_L g4712 ( 
.A(n_4407),
.B(n_3479),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_3952),
.Y(n_4713)
);

HB1xp67_ASAP7_75t_L g4714 ( 
.A(n_4382),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4445),
.Y(n_4715)
);

AND2x2_ASAP7_75t_L g4716 ( 
.A(n_4067),
.B(n_2626),
.Y(n_4716)
);

O2A1O1Ixp5_ASAP7_75t_L g4717 ( 
.A1(n_4069),
.A2(n_3904),
.B(n_3692),
.C(n_3760),
.Y(n_4717)
);

NOR2xp33_ASAP7_75t_L g4718 ( 
.A(n_4099),
.B(n_3942),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4180),
.B(n_4160),
.Y(n_4719)
);

INVx2_ASAP7_75t_L g4720 ( 
.A(n_3955),
.Y(n_4720)
);

AND2x4_ASAP7_75t_L g4721 ( 
.A(n_3965),
.B(n_3492),
.Y(n_4721)
);

INVx2_ASAP7_75t_L g4722 ( 
.A(n_3957),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4282),
.B(n_3222),
.Y(n_4723)
);

OR2x2_ASAP7_75t_L g4724 ( 
.A(n_3947),
.B(n_3225),
.Y(n_4724)
);

AOI22xp5_ASAP7_75t_L g4725 ( 
.A1(n_4177),
.A2(n_3837),
.B1(n_3727),
.B2(n_3399),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_L g4726 ( 
.A(n_4282),
.B(n_3235),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4190),
.B(n_3237),
.Y(n_4727)
);

NOR3xp33_ASAP7_75t_L g4728 ( 
.A(n_4141),
.B(n_1288),
.C(n_947),
.Y(n_4728)
);

NAND2xp5_ASAP7_75t_L g4729 ( 
.A(n_4196),
.B(n_3239),
.Y(n_4729)
);

INVx2_ASAP7_75t_SL g4730 ( 
.A(n_4182),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_SL g4731 ( 
.A(n_4386),
.B(n_3424),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_SL g4732 ( 
.A(n_4416),
.B(n_3481),
.Y(n_4732)
);

NOR2xp33_ASAP7_75t_SL g4733 ( 
.A(n_4185),
.B(n_3660),
.Y(n_4733)
);

INVx1_ASAP7_75t_L g4734 ( 
.A(n_3960),
.Y(n_4734)
);

INVx3_ASAP7_75t_L g4735 ( 
.A(n_3997),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_L g4736 ( 
.A(n_4196),
.B(n_3240),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_3963),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4151),
.B(n_3243),
.Y(n_4738)
);

INVx2_ASAP7_75t_L g4739 ( 
.A(n_3971),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4151),
.B(n_3245),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_3975),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4382),
.B(n_3248),
.Y(n_4742)
);

NOR2xp67_ASAP7_75t_SL g4743 ( 
.A(n_4202),
.B(n_4216),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4423),
.B(n_3257),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4441),
.B(n_4135),
.Y(n_4745)
);

AOI22xp33_ASAP7_75t_L g4746 ( 
.A1(n_3969),
.A2(n_3837),
.B1(n_3457),
.B2(n_3369),
.Y(n_4746)
);

AOI22xp5_ASAP7_75t_L g4747 ( 
.A1(n_4031),
.A2(n_3727),
.B1(n_3382),
.B2(n_3399),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4371),
.B(n_2626),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4141),
.B(n_3367),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_3976),
.B(n_2586),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_SL g4751 ( 
.A(n_4413),
.B(n_4092),
.Y(n_4751)
);

OR2x6_ASAP7_75t_L g4752 ( 
.A(n_4120),
.B(n_3715),
.Y(n_4752)
);

NAND2x1_ASAP7_75t_L g4753 ( 
.A(n_4408),
.B(n_3382),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_3979),
.B(n_2641),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_3981),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_3982),
.B(n_2641),
.Y(n_4756)
);

OR2x2_ASAP7_75t_L g4757 ( 
.A(n_4206),
.B(n_2641),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_SL g4758 ( 
.A(n_4413),
.B(n_3481),
.Y(n_4758)
);

AOI221xp5_ASAP7_75t_L g4759 ( 
.A1(n_4308),
.A2(n_980),
.B1(n_1002),
.B2(n_978),
.C(n_849),
.Y(n_4759)
);

INVx2_ASAP7_75t_SL g4760 ( 
.A(n_4397),
.Y(n_4760)
);

AND2x2_ASAP7_75t_L g4761 ( 
.A(n_4224),
.B(n_2626),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_3984),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_SL g4763 ( 
.A(n_4092),
.B(n_4108),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_3985),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4367),
.B(n_2627),
.Y(n_4765)
);

OAI221xp5_ASAP7_75t_L g4766 ( 
.A1(n_3996),
.A2(n_2618),
.B1(n_2643),
.B2(n_2622),
.C(n_2617),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_3991),
.B(n_2649),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_3992),
.Y(n_4768)
);

OAI22xp5_ASAP7_75t_SL g4769 ( 
.A1(n_4317),
.A2(n_1231),
.B1(n_1301),
.B2(n_1132),
.Y(n_4769)
);

NOR2xp33_ASAP7_75t_SL g4770 ( 
.A(n_4288),
.B(n_3660),
.Y(n_4770)
);

INVxp33_ASAP7_75t_L g4771 ( 
.A(n_4384),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_3994),
.B(n_2649),
.Y(n_4772)
);

BUFx3_ASAP7_75t_L g4773 ( 
.A(n_4343),
.Y(n_4773)
);

O2A1O1Ixp5_ASAP7_75t_L g4774 ( 
.A1(n_4274),
.A2(n_3760),
.B(n_3768),
.C(n_3700),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_SL g4775 ( 
.A(n_4108),
.B(n_3481),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_3998),
.B(n_4002),
.Y(n_4776)
);

CKINVDCx20_ASAP7_75t_R g4777 ( 
.A(n_4285),
.Y(n_4777)
);

AND2x2_ASAP7_75t_L g4778 ( 
.A(n_4403),
.B(n_4014),
.Y(n_4778)
);

INVx2_ASAP7_75t_L g4779 ( 
.A(n_4004),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4005),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4007),
.B(n_4008),
.Y(n_4781)
);

A2O1A1Ixp33_ASAP7_75t_L g4782 ( 
.A1(n_4419),
.A2(n_3944),
.B(n_3715),
.C(n_3312),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4009),
.Y(n_4783)
);

NOR2xp33_ASAP7_75t_L g4784 ( 
.A(n_4150),
.B(n_3399),
.Y(n_4784)
);

AOI22xp33_ASAP7_75t_L g4785 ( 
.A1(n_4260),
.A2(n_4375),
.B1(n_4152),
.B2(n_4352),
.Y(n_4785)
);

AND2x2_ASAP7_75t_L g4786 ( 
.A(n_4401),
.B(n_2627),
.Y(n_4786)
);

INVx2_ASAP7_75t_L g4787 ( 
.A(n_4020),
.Y(n_4787)
);

AND2x6_ASAP7_75t_SL g4788 ( 
.A(n_4094),
.B(n_1390),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4021),
.B(n_2649),
.Y(n_4789)
);

OR2x6_ASAP7_75t_L g4790 ( 
.A(n_3997),
.B(n_3715),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4430),
.B(n_2627),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4024),
.B(n_2686),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4025),
.B(n_2686),
.Y(n_4793)
);

AND2x6_ASAP7_75t_SL g4794 ( 
.A(n_4098),
.B(n_1390),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4035),
.B(n_2686),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4037),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4038),
.B(n_2645),
.Y(n_4797)
);

OAI22xp33_ASAP7_75t_L g4798 ( 
.A1(n_4011),
.A2(n_1231),
.B1(n_1301),
.B2(n_1132),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_SL g4799 ( 
.A(n_4150),
.B(n_3481),
.Y(n_4799)
);

NOR2xp33_ASAP7_75t_L g4800 ( 
.A(n_4107),
.B(n_2497),
.Y(n_4800)
);

AOI22xp33_ASAP7_75t_L g4801 ( 
.A1(n_4260),
.A2(n_3457),
.B1(n_2726),
.B2(n_2737),
.Y(n_4801)
);

NOR2xp33_ASAP7_75t_L g4802 ( 
.A(n_4113),
.B(n_2497),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4042),
.B(n_2650),
.Y(n_4803)
);

AOI22xp33_ASAP7_75t_L g4804 ( 
.A1(n_4011),
.A2(n_2726),
.B1(n_2737),
.B2(n_2729),
.Y(n_4804)
);

NOR2xp33_ASAP7_75t_L g4805 ( 
.A(n_4414),
.B(n_2522),
.Y(n_4805)
);

INVx8_ASAP7_75t_L g4806 ( 
.A(n_4387),
.Y(n_4806)
);

AND2x2_ASAP7_75t_L g4807 ( 
.A(n_4093),
.B(n_944),
.Y(n_4807)
);

AND2x2_ASAP7_75t_L g4808 ( 
.A(n_3958),
.B(n_1160),
.Y(n_4808)
);

O2A1O1Ixp5_ASAP7_75t_L g4809 ( 
.A1(n_4274),
.A2(n_3760),
.B(n_3768),
.C(n_3700),
.Y(n_4809)
);

BUFx5_ASAP7_75t_L g4810 ( 
.A(n_4017),
.Y(n_4810)
);

NOR2xp33_ASAP7_75t_L g4811 ( 
.A(n_4414),
.B(n_2522),
.Y(n_4811)
);

AND2x2_ASAP7_75t_L g4812 ( 
.A(n_4061),
.B(n_1160),
.Y(n_4812)
);

OAI22xp5_ASAP7_75t_L g4813 ( 
.A1(n_4376),
.A2(n_3533),
.B1(n_3585),
.B2(n_3549),
.Y(n_4813)
);

INVx2_ASAP7_75t_L g4814 ( 
.A(n_4044),
.Y(n_4814)
);

OAI21xp5_ASAP7_75t_L g4815 ( 
.A1(n_4439),
.A2(n_3727),
.B(n_3420),
.Y(n_4815)
);

AND2x2_ASAP7_75t_L g4816 ( 
.A(n_4256),
.B(n_1160),
.Y(n_4816)
);

NOR2xp33_ASAP7_75t_L g4817 ( 
.A(n_4290),
.B(n_2543),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_SL g4818 ( 
.A(n_4294),
.B(n_3481),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4047),
.Y(n_4819)
);

NOR3xp33_ASAP7_75t_L g4820 ( 
.A(n_4419),
.B(n_947),
.C(n_932),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_SL g4821 ( 
.A(n_4294),
.B(n_3507),
.Y(n_4821)
);

NOR2xp33_ASAP7_75t_L g4822 ( 
.A(n_4316),
.B(n_2543),
.Y(n_4822)
);

INVx2_ASAP7_75t_L g4823 ( 
.A(n_4048),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4050),
.B(n_2661),
.Y(n_4824)
);

OAI21xp5_ASAP7_75t_L g4825 ( 
.A1(n_4439),
.A2(n_3727),
.B(n_3312),
.Y(n_4825)
);

INVxp67_ASAP7_75t_L g4826 ( 
.A(n_4051),
.Y(n_4826)
);

INVx1_ASAP7_75t_L g4827 ( 
.A(n_4052),
.Y(n_4827)
);

BUFx3_ASAP7_75t_L g4828 ( 
.A(n_4256),
.Y(n_4828)
);

AND2x2_ASAP7_75t_L g4829 ( 
.A(n_4435),
.B(n_1160),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4053),
.Y(n_4830)
);

INVx2_ASAP7_75t_SL g4831 ( 
.A(n_4220),
.Y(n_4831)
);

NAND2xp5_ASAP7_75t_L g4832 ( 
.A(n_4054),
.B(n_4055),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_SL g4833 ( 
.A(n_4294),
.B(n_3507),
.Y(n_4833)
);

NOR2xp33_ASAP7_75t_L g4834 ( 
.A(n_4409),
.B(n_3492),
.Y(n_4834)
);

NOR2xp33_ASAP7_75t_L g4835 ( 
.A(n_4409),
.B(n_3509),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_SL g4836 ( 
.A(n_4294),
.B(n_3507),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4058),
.B(n_2663),
.Y(n_4837)
);

AOI22xp33_ASAP7_75t_L g4838 ( 
.A1(n_4012),
.A2(n_2729),
.B1(n_2743),
.B2(n_2737),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_4059),
.B(n_2680),
.Y(n_4839)
);

NAND3xp33_ASAP7_75t_L g4840 ( 
.A(n_4051),
.B(n_2737),
.C(n_2729),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_SL g4841 ( 
.A(n_4294),
.B(n_3507),
.Y(n_4841)
);

NOR2xp67_ASAP7_75t_L g4842 ( 
.A(n_4444),
.B(n_3441),
.Y(n_4842)
);

INVx2_ASAP7_75t_SL g4843 ( 
.A(n_4328),
.Y(n_4843)
);

INVx2_ASAP7_75t_L g4844 ( 
.A(n_4060),
.Y(n_4844)
);

AOI22xp5_ASAP7_75t_L g4845 ( 
.A1(n_4349),
.A2(n_3727),
.B1(n_3848),
.B2(n_2959),
.Y(n_4845)
);

AOI22xp5_ASAP7_75t_L g4846 ( 
.A1(n_4349),
.A2(n_3848),
.B1(n_2959),
.B2(n_2985),
.Y(n_4846)
);

INVx2_ASAP7_75t_L g4847 ( 
.A(n_4062),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_SL g4848 ( 
.A(n_4294),
.B(n_3507),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4063),
.Y(n_4849)
);

OAI21xp33_ASAP7_75t_L g4850 ( 
.A1(n_4370),
.A2(n_957),
.B(n_953),
.Y(n_4850)
);

BUFx3_ASAP7_75t_L g4851 ( 
.A(n_4422),
.Y(n_4851)
);

INVx2_ASAP7_75t_L g4852 ( 
.A(n_4064),
.Y(n_4852)
);

INVx2_ASAP7_75t_L g4853 ( 
.A(n_4065),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_L g4854 ( 
.A(n_4066),
.B(n_2682),
.Y(n_4854)
);

NAND2xp5_ASAP7_75t_L g4855 ( 
.A(n_4068),
.B(n_2689),
.Y(n_4855)
);

NOR2xp33_ASAP7_75t_L g4856 ( 
.A(n_4428),
.B(n_3509),
.Y(n_4856)
);

NAND2x1p5_ASAP7_75t_L g4857 ( 
.A(n_4405),
.B(n_3509),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4070),
.B(n_2695),
.Y(n_4858)
);

NOR3xp33_ASAP7_75t_L g4859 ( 
.A(n_4359),
.B(n_954),
.C(n_932),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4072),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4073),
.B(n_2708),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4074),
.B(n_2711),
.Y(n_4862)
);

NAND2xp5_ASAP7_75t_SL g4863 ( 
.A(n_4013),
.B(n_3574),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4075),
.B(n_2718),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4082),
.B(n_2721),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4085),
.B(n_2724),
.Y(n_4866)
);

INVx4_ASAP7_75t_L g4867 ( 
.A(n_4013),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_L g4868 ( 
.A(n_4086),
.B(n_2732),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4088),
.B(n_2747),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_SL g4870 ( 
.A(n_4468),
.B(n_4013),
.Y(n_4870)
);

INVx2_ASAP7_75t_L g4871 ( 
.A(n_4448),
.Y(n_4871)
);

AO22x1_ASAP7_75t_L g4872 ( 
.A1(n_4484),
.A2(n_4077),
.B1(n_4118),
.B2(n_4012),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4451),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_SL g4874 ( 
.A(n_4463),
.B(n_4465),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4711),
.B(n_4090),
.Y(n_4875)
);

INVx1_ASAP7_75t_L g4876 ( 
.A(n_4713),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4462),
.B(n_4459),
.Y(n_4877)
);

BUFx12f_ASAP7_75t_SL g4878 ( 
.A(n_4518),
.Y(n_4878)
);

HB1xp67_ASAP7_75t_L g4879 ( 
.A(n_4513),
.Y(n_4879)
);

AOI22xp33_ASAP7_75t_SL g4880 ( 
.A1(n_4769),
.A2(n_4118),
.B1(n_4077),
.B2(n_4387),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4521),
.B(n_4095),
.Y(n_4881)
);

NOR3xp33_ASAP7_75t_SL g4882 ( 
.A(n_4681),
.B(n_964),
.C(n_963),
.Y(n_4882)
);

INVx4_ASAP7_75t_L g4883 ( 
.A(n_4478),
.Y(n_4883)
);

INVx2_ASAP7_75t_L g4884 ( 
.A(n_4452),
.Y(n_4884)
);

NAND2xp5_ASAP7_75t_L g4885 ( 
.A(n_4521),
.B(n_4096),
.Y(n_4885)
);

NAND2x1p5_ASAP7_75t_L g4886 ( 
.A(n_4690),
.B(n_4418),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4720),
.Y(n_4887)
);

AND2x4_ASAP7_75t_L g4888 ( 
.A(n_4559),
.B(n_4422),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4722),
.Y(n_4889)
);

NOR2xp33_ASAP7_75t_L g4890 ( 
.A(n_4454),
.B(n_1331),
.Y(n_4890)
);

OAI22xp33_ASAP7_75t_L g4891 ( 
.A1(n_4491),
.A2(n_4325),
.B1(n_3915),
.B2(n_3818),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4719),
.B(n_4100),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4624),
.B(n_4101),
.Y(n_4893)
);

AND2x4_ASAP7_75t_L g4894 ( 
.A(n_4559),
.B(n_4102),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4737),
.Y(n_4895)
);

BUFx6f_ASAP7_75t_L g4896 ( 
.A(n_4534),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_SL g4897 ( 
.A(n_4492),
.B(n_4015),
.Y(n_4897)
);

CKINVDCx5p33_ASAP7_75t_R g4898 ( 
.A(n_4478),
.Y(n_4898)
);

NOR2xp33_ASAP7_75t_R g4899 ( 
.A(n_4699),
.B(n_4325),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_SL g4900 ( 
.A(n_4616),
.B(n_4015),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4553),
.B(n_4105),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_L g4902 ( 
.A(n_4553),
.B(n_4106),
.Y(n_4902)
);

INVx2_ASAP7_75t_L g4903 ( 
.A(n_4479),
.Y(n_4903)
);

BUFx3_ASAP7_75t_L g4904 ( 
.A(n_4543),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4739),
.Y(n_4905)
);

INVx1_ASAP7_75t_L g4906 ( 
.A(n_4779),
.Y(n_4906)
);

AOI21xp5_ASAP7_75t_L g4907 ( 
.A1(n_4609),
.A2(n_4532),
.B(n_4667),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4645),
.B(n_4109),
.Y(n_4908)
);

AND2x4_ASAP7_75t_L g4909 ( 
.A(n_4690),
.B(n_4110),
.Y(n_4909)
);

INVx5_ASAP7_75t_L g4910 ( 
.A(n_4630),
.Y(n_4910)
);

INVx2_ASAP7_75t_SL g4911 ( 
.A(n_4688),
.Y(n_4911)
);

NOR3xp33_ASAP7_75t_L g4912 ( 
.A(n_4464),
.B(n_979),
.C(n_954),
.Y(n_4912)
);

NOR3xp33_ASAP7_75t_SL g4913 ( 
.A(n_4701),
.B(n_970),
.C(n_965),
.Y(n_4913)
);

BUFx12f_ASAP7_75t_SL g4914 ( 
.A(n_4518),
.Y(n_4914)
);

NOR2xp67_ASAP7_75t_L g4915 ( 
.A(n_4552),
.B(n_3700),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4659),
.B(n_1331),
.Y(n_4916)
);

BUFx4f_ASAP7_75t_L g4917 ( 
.A(n_4620),
.Y(n_4917)
);

NAND2xp5_ASAP7_75t_SL g4918 ( 
.A(n_4616),
.B(n_4015),
.Y(n_4918)
);

AOI22xp5_ASAP7_75t_L g4919 ( 
.A1(n_4480),
.A2(n_4349),
.B1(n_4019),
.B2(n_4017),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4787),
.Y(n_4920)
);

AOI22xp33_ASAP7_75t_SL g4921 ( 
.A1(n_4449),
.A2(n_4349),
.B1(n_4019),
.B2(n_4017),
.Y(n_4921)
);

INVx2_ASAP7_75t_L g4922 ( 
.A(n_4483),
.Y(n_4922)
);

BUFx2_ASAP7_75t_L g4923 ( 
.A(n_4458),
.Y(n_4923)
);

INVx2_ASAP7_75t_SL g4924 ( 
.A(n_4773),
.Y(n_4924)
);

INVx2_ASAP7_75t_L g4925 ( 
.A(n_4503),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4814),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4819),
.Y(n_4927)
);

INVx2_ASAP7_75t_L g4928 ( 
.A(n_4507),
.Y(n_4928)
);

INVx1_ASAP7_75t_L g4929 ( 
.A(n_4823),
.Y(n_4929)
);

INVx2_ASAP7_75t_L g4930 ( 
.A(n_4516),
.Y(n_4930)
);

BUFx6f_ASAP7_75t_L g4931 ( 
.A(n_4534),
.Y(n_4931)
);

NAND2xp5_ASAP7_75t_SL g4932 ( 
.A(n_4510),
.B(n_4489),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4598),
.B(n_4618),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4844),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4522),
.Y(n_4935)
);

AOI21xp5_ASAP7_75t_L g4936 ( 
.A1(n_4532),
.A2(n_4354),
.B(n_4097),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4598),
.B(n_4618),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_SL g4938 ( 
.A(n_4510),
.B(n_4015),
.Y(n_4938)
);

AND2x4_ASAP7_75t_L g4939 ( 
.A(n_4690),
.B(n_4111),
.Y(n_4939)
);

INVx2_ASAP7_75t_L g4940 ( 
.A(n_4525),
.Y(n_4940)
);

AND2x6_ASAP7_75t_SL g4941 ( 
.A(n_4621),
.B(n_1408),
.Y(n_4941)
);

HB1xp67_ASAP7_75t_L g4942 ( 
.A(n_4513),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4535),
.Y(n_4943)
);

INVx2_ASAP7_75t_L g4944 ( 
.A(n_4537),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4847),
.Y(n_4945)
);

A2O1A1Ixp33_ASAP7_75t_L g4946 ( 
.A1(n_4519),
.A2(n_4359),
.B(n_4443),
.C(n_4428),
.Y(n_4946)
);

INVx2_ASAP7_75t_L g4947 ( 
.A(n_4546),
.Y(n_4947)
);

INVx1_ASAP7_75t_L g4948 ( 
.A(n_4852),
.Y(n_4948)
);

BUFx3_ASAP7_75t_L g4949 ( 
.A(n_4664),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4645),
.B(n_4112),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4853),
.Y(n_4951)
);

INVx3_ASAP7_75t_L g4952 ( 
.A(n_4534),
.Y(n_4952)
);

OAI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_4476),
.A2(n_4116),
.B1(n_4119),
.B2(n_4114),
.Y(n_4953)
);

AOI21xp33_ASAP7_75t_L g4954 ( 
.A1(n_4481),
.A2(n_4370),
.B(n_4443),
.Y(n_4954)
);

CKINVDCx8_ASAP7_75t_R g4955 ( 
.A(n_4636),
.Y(n_4955)
);

AND2x4_ASAP7_75t_L g4956 ( 
.A(n_4690),
.B(n_4124),
.Y(n_4956)
);

A2O1A1Ixp33_ASAP7_75t_L g4957 ( 
.A1(n_4533),
.A2(n_4126),
.B(n_4128),
.C(n_4125),
.Y(n_4957)
);

NOR2xp33_ASAP7_75t_L g4958 ( 
.A(n_4457),
.B(n_1440),
.Y(n_4958)
);

INVx2_ASAP7_75t_L g4959 ( 
.A(n_4548),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4527),
.Y(n_4960)
);

INVx1_ASAP7_75t_SL g4961 ( 
.A(n_4605),
.Y(n_4961)
);

INVx2_ASAP7_75t_L g4962 ( 
.A(n_4556),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4563),
.Y(n_4963)
);

OAI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4640),
.A2(n_4137),
.B(n_4307),
.Y(n_4964)
);

BUFx3_ASAP7_75t_L g4965 ( 
.A(n_4777),
.Y(n_4965)
);

O2A1O1Ixp33_ASAP7_75t_L g4966 ( 
.A1(n_4505),
.A2(n_1440),
.B(n_979),
.C(n_996),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4536),
.Y(n_4967)
);

BUFx6f_ASAP7_75t_L g4968 ( 
.A(n_4582),
.Y(n_4968)
);

NOR2xp33_ASAP7_75t_L g4969 ( 
.A(n_4566),
.B(n_1214),
.Y(n_4969)
);

INVx5_ASAP7_75t_L g4970 ( 
.A(n_4630),
.Y(n_4970)
);

BUFx2_ASAP7_75t_L g4971 ( 
.A(n_4458),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_SL g4972 ( 
.A(n_4826),
.B(n_4022),
.Y(n_4972)
);

INVx1_ASAP7_75t_L g4973 ( 
.A(n_4558),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4565),
.Y(n_4974)
);

A2O1A1Ixp33_ASAP7_75t_L g4975 ( 
.A1(n_4464),
.A2(n_4131),
.B(n_4132),
.C(n_4130),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4834),
.B(n_4835),
.Y(n_4976)
);

AND2x2_ASAP7_75t_L g4977 ( 
.A(n_4541),
.B(n_1178),
.Y(n_4977)
);

AND2x4_ASAP7_75t_L g4978 ( 
.A(n_4721),
.B(n_4133),
.Y(n_4978)
);

NOR2xp33_ASAP7_75t_L g4979 ( 
.A(n_4648),
.B(n_4635),
.Y(n_4979)
);

A2O1A1Ixp33_ASAP7_75t_L g4980 ( 
.A1(n_4785),
.A2(n_4139),
.B(n_4140),
.C(n_4134),
.Y(n_4980)
);

NOR2xp33_ASAP7_75t_R g4981 ( 
.A(n_4705),
.B(n_4022),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4622),
.B(n_4144),
.Y(n_4982)
);

INVx1_ASAP7_75t_SL g4983 ( 
.A(n_4605),
.Y(n_4983)
);

BUFx6f_ASAP7_75t_L g4984 ( 
.A(n_4582),
.Y(n_4984)
);

NAND2xp5_ASAP7_75t_L g4985 ( 
.A(n_4482),
.B(n_4145),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4571),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4575),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4473),
.B(n_4149),
.Y(n_4988)
);

INVx2_ASAP7_75t_L g4989 ( 
.A(n_4572),
.Y(n_4989)
);

NOR2xp33_ASAP7_75t_R g4990 ( 
.A(n_4549),
.B(n_4022),
.Y(n_4990)
);

BUFx2_ASAP7_75t_L g4991 ( 
.A(n_4676),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4601),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4476),
.B(n_4154),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_4834),
.B(n_4155),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4585),
.Y(n_4995)
);

NAND2xp5_ASAP7_75t_L g4996 ( 
.A(n_4835),
.B(n_4156),
.Y(n_4996)
);

HB1xp67_ASAP7_75t_L g4997 ( 
.A(n_4473),
.Y(n_4997)
);

INVx3_ASAP7_75t_L g4998 ( 
.A(n_4582),
.Y(n_4998)
);

AOI22xp33_ASAP7_75t_L g4999 ( 
.A1(n_4567),
.A2(n_2743),
.B1(n_2757),
.B2(n_2729),
.Y(n_4999)
);

AND2x4_ASAP7_75t_L g5000 ( 
.A(n_4721),
.B(n_4157),
.Y(n_5000)
);

AO22x1_ASAP7_75t_L g5001 ( 
.A1(n_4820),
.A2(n_974),
.B1(n_984),
.B2(n_983),
.Y(n_5001)
);

OR2x2_ASAP7_75t_SL g5002 ( 
.A(n_4494),
.B(n_1408),
.Y(n_5002)
);

INVx2_ASAP7_75t_SL g5003 ( 
.A(n_4806),
.Y(n_5003)
);

INVx1_ASAP7_75t_L g5004 ( 
.A(n_4590),
.Y(n_5004)
);

OR2x6_ASAP7_75t_SL g5005 ( 
.A(n_4574),
.B(n_987),
.Y(n_5005)
);

AND2x6_ASAP7_75t_L g5006 ( 
.A(n_4685),
.B(n_4161),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4592),
.Y(n_5007)
);

CKINVDCx5p33_ASAP7_75t_R g5008 ( 
.A(n_4788),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_SL g5009 ( 
.A(n_4826),
.B(n_4022),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4594),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4856),
.B(n_4162),
.Y(n_5011)
);

AOI22xp5_ASAP7_75t_L g5012 ( 
.A1(n_4643),
.A2(n_4349),
.B1(n_4019),
.B2(n_4017),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_4749),
.B(n_4165),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_SL g5014 ( 
.A(n_4805),
.B(n_4084),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4526),
.B(n_4166),
.Y(n_5015)
);

INVx2_ASAP7_75t_L g5016 ( 
.A(n_4652),
.Y(n_5016)
);

NOR2xp33_ASAP7_75t_R g5017 ( 
.A(n_4461),
.B(n_4084),
.Y(n_5017)
);

CKINVDCx14_ASAP7_75t_R g5018 ( 
.A(n_4539),
.Y(n_5018)
);

BUFx6f_ASAP7_75t_L g5019 ( 
.A(n_4806),
.Y(n_5019)
);

NOR2xp33_ASAP7_75t_L g5020 ( 
.A(n_4456),
.B(n_1215),
.Y(n_5020)
);

BUFx2_ASAP7_75t_L g5021 ( 
.A(n_4676),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4597),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4856),
.B(n_4763),
.Y(n_5023)
);

INVx2_ASAP7_75t_L g5024 ( 
.A(n_4654),
.Y(n_5024)
);

AND2x4_ASAP7_75t_L g5025 ( 
.A(n_4752),
.B(n_4682),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_L g5026 ( 
.A(n_4506),
.B(n_4714),
.Y(n_5026)
);

INVx2_ASAP7_75t_L g5027 ( 
.A(n_4657),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4610),
.Y(n_5028)
);

NAND2xp5_ASAP7_75t_L g5029 ( 
.A(n_4727),
.B(n_4167),
.Y(n_5029)
);

AOI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_4667),
.A2(n_4354),
.B(n_4385),
.Y(n_5030)
);

INVx2_ASAP7_75t_L g5031 ( 
.A(n_4666),
.Y(n_5031)
);

NOR2xp33_ASAP7_75t_L g5032 ( 
.A(n_4577),
.B(n_1218),
.Y(n_5032)
);

AND3x1_ASAP7_75t_L g5033 ( 
.A(n_4728),
.B(n_990),
.C(n_952),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_SL g5034 ( 
.A(n_4811),
.B(n_4084),
.Y(n_5034)
);

AOI22xp33_ASAP7_75t_L g5035 ( 
.A1(n_4567),
.A2(n_4496),
.B1(n_4785),
.B2(n_4759),
.Y(n_5035)
);

INVx2_ASAP7_75t_SL g5036 ( 
.A(n_4806),
.Y(n_5036)
);

AND2x6_ASAP7_75t_SL g5037 ( 
.A(n_4631),
.B(n_1410),
.Y(n_5037)
);

O2A1O1Ixp33_ASAP7_75t_L g5038 ( 
.A1(n_4728),
.A2(n_996),
.B(n_1000),
.C(n_992),
.Y(n_5038)
);

INVx1_ASAP7_75t_L g5039 ( 
.A(n_4612),
.Y(n_5039)
);

AOI22xp5_ASAP7_75t_L g5040 ( 
.A1(n_4820),
.A2(n_4019),
.B1(n_4017),
.B2(n_2624),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4615),
.Y(n_5041)
);

AOI21xp5_ASAP7_75t_L g5042 ( 
.A1(n_4644),
.A2(n_4385),
.B(n_4137),
.Y(n_5042)
);

INVx1_ASAP7_75t_L g5043 ( 
.A(n_4625),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_SL g5044 ( 
.A(n_4471),
.B(n_4084),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4634),
.Y(n_5045)
);

AOI22xp33_ASAP7_75t_L g5046 ( 
.A1(n_4496),
.A2(n_2757),
.B1(n_2743),
.B2(n_2570),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4642),
.Y(n_5047)
);

INVx1_ASAP7_75t_L g5048 ( 
.A(n_4647),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4673),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_SL g5050 ( 
.A(n_4725),
.B(n_4170),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_4679),
.Y(n_5051)
);

OAI21xp5_ASAP7_75t_L g5052 ( 
.A1(n_4859),
.A2(n_4307),
.B(n_4210),
.Y(n_5052)
);

NOR2xp33_ASAP7_75t_L g5053 ( 
.A(n_4560),
.B(n_1225),
.Y(n_5053)
);

INVx1_ASAP7_75t_L g5054 ( 
.A(n_4651),
.Y(n_5054)
);

OAI22xp5_ASAP7_75t_L g5055 ( 
.A1(n_4531),
.A2(n_4588),
.B1(n_4846),
.B2(n_4756),
.Y(n_5055)
);

NOR3xp33_ASAP7_75t_SL g5056 ( 
.A(n_4583),
.B(n_999),
.C(n_994),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_4714),
.B(n_4172),
.Y(n_5057)
);

BUFx8_ASAP7_75t_L g5058 ( 
.A(n_4469),
.Y(n_5058)
);

INVx3_ASAP7_75t_L g5059 ( 
.A(n_4682),
.Y(n_5059)
);

NAND2x1p5_ASAP7_75t_L g5060 ( 
.A(n_4753),
.B(n_4538),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4694),
.Y(n_5061)
);

BUFx2_ASAP7_75t_L g5062 ( 
.A(n_4828),
.Y(n_5062)
);

BUFx2_ASAP7_75t_L g5063 ( 
.A(n_4851),
.Y(n_5063)
);

AND2x4_ASAP7_75t_L g5064 ( 
.A(n_4752),
.B(n_4174),
.Y(n_5064)
);

BUFx3_ASAP7_75t_L g5065 ( 
.A(n_4760),
.Y(n_5065)
);

NAND2xp5_ASAP7_75t_SL g5066 ( 
.A(n_4620),
.B(n_4170),
.Y(n_5066)
);

NOR2xp33_ASAP7_75t_L g5067 ( 
.A(n_4691),
.B(n_1228),
.Y(n_5067)
);

INVx1_ASAP7_75t_SL g5068 ( 
.A(n_4515),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4658),
.Y(n_5069)
);

NOR2xp33_ASAP7_75t_L g5070 ( 
.A(n_4540),
.B(n_1241),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4668),
.Y(n_5071)
);

AOI22xp5_ASAP7_75t_L g5072 ( 
.A1(n_4674),
.A2(n_4019),
.B1(n_2624),
.B2(n_2630),
.Y(n_5072)
);

BUFx3_ASAP7_75t_L g5073 ( 
.A(n_4467),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4680),
.Y(n_5074)
);

OR2x2_ASAP7_75t_L g5075 ( 
.A(n_4544),
.B(n_4724),
.Y(n_5075)
);

NAND2xp5_ASAP7_75t_SL g5076 ( 
.A(n_4632),
.B(n_4170),
.Y(n_5076)
);

AND2x4_ASAP7_75t_L g5077 ( 
.A(n_4752),
.B(n_4178),
.Y(n_5077)
);

BUFx10_ASAP7_75t_L g5078 ( 
.A(n_4817),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_SL g5079 ( 
.A(n_4729),
.B(n_4170),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4736),
.B(n_4181),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4684),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_SL g5082 ( 
.A(n_4702),
.B(n_4291),
.Y(n_5082)
);

OAI22xp33_ASAP7_75t_L g5083 ( 
.A1(n_4564),
.A2(n_3915),
.B1(n_3818),
.B2(n_4408),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4687),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_4707),
.B(n_4183),
.Y(n_5085)
);

BUFx3_ASAP7_75t_L g5086 ( 
.A(n_4730),
.Y(n_5086)
);

AOI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4674),
.A2(n_2624),
.B1(n_2630),
.B2(n_2604),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_SL g5088 ( 
.A(n_4747),
.B(n_4291),
.Y(n_5088)
);

INVx2_ASAP7_75t_SL g5089 ( 
.A(n_4831),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4692),
.Y(n_5090)
);

OAI22xp5_ASAP7_75t_SL g5091 ( 
.A1(n_4568),
.A2(n_1000),
.B1(n_1009),
.B2(n_992),
.Y(n_5091)
);

INVx3_ASAP7_75t_L g5092 ( 
.A(n_4630),
.Y(n_5092)
);

A2O1A1Ixp33_ASAP7_75t_L g5093 ( 
.A1(n_4481),
.A2(n_4188),
.B(n_4192),
.C(n_4187),
.Y(n_5093)
);

INVx2_ASAP7_75t_SL g5094 ( 
.A(n_4843),
.Y(n_5094)
);

AOI22xp5_ASAP7_75t_L g5095 ( 
.A1(n_4606),
.A2(n_2624),
.B1(n_2630),
.B2(n_2604),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_4698),
.Y(n_5096)
);

INVx5_ASAP7_75t_L g5097 ( 
.A(n_4630),
.Y(n_5097)
);

AOI22xp33_ASAP7_75t_L g5098 ( 
.A1(n_4759),
.A2(n_2757),
.B1(n_2743),
.B2(n_2570),
.Y(n_5098)
);

INVx1_ASAP7_75t_L g5099 ( 
.A(n_4703),
.Y(n_5099)
);

INVx1_ASAP7_75t_L g5100 ( 
.A(n_4704),
.Y(n_5100)
);

INVxp67_ASAP7_75t_L g5101 ( 
.A(n_4488),
.Y(n_5101)
);

NOR2xp33_ASAP7_75t_L g5102 ( 
.A(n_4745),
.B(n_1243),
.Y(n_5102)
);

HB1xp67_ASAP7_75t_L g5103 ( 
.A(n_4599),
.Y(n_5103)
);

NAND3xp33_ASAP7_75t_L g5104 ( 
.A(n_4859),
.B(n_990),
.C(n_952),
.Y(n_5104)
);

BUFx4f_ASAP7_75t_SL g5105 ( 
.A(n_4627),
.Y(n_5105)
);

NAND2xp33_ASAP7_75t_L g5106 ( 
.A(n_4561),
.B(n_4291),
.Y(n_5106)
);

INVx2_ASAP7_75t_SL g5107 ( 
.A(n_4475),
.Y(n_5107)
);

NAND2xp5_ASAP7_75t_L g5108 ( 
.A(n_4628),
.B(n_4194),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4715),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_4629),
.B(n_4197),
.Y(n_5110)
);

NAND2x1p5_ASAP7_75t_L g5111 ( 
.A(n_4580),
.B(n_3576),
.Y(n_5111)
);

NAND2xp5_ASAP7_75t_SL g5112 ( 
.A(n_4520),
.B(n_4291),
.Y(n_5112)
);

BUFx6f_ASAP7_75t_L g5113 ( 
.A(n_4576),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4734),
.Y(n_5114)
);

INVx1_ASAP7_75t_L g5115 ( 
.A(n_4741),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4755),
.Y(n_5116)
);

AND2x4_ASAP7_75t_L g5117 ( 
.A(n_4675),
.B(n_4198),
.Y(n_5117)
);

CKINVDCx5p33_ASAP7_75t_R g5118 ( 
.A(n_4794),
.Y(n_5118)
);

BUFx8_ASAP7_75t_L g5119 ( 
.A(n_4816),
.Y(n_5119)
);

INVx5_ASAP7_75t_L g5120 ( 
.A(n_4630),
.Y(n_5120)
);

NOR2xp33_ASAP7_75t_R g5121 ( 
.A(n_4498),
.B(n_4399),
.Y(n_5121)
);

INVx1_ASAP7_75t_L g5122 ( 
.A(n_4762),
.Y(n_5122)
);

CKINVDCx5p33_ASAP7_75t_R g5123 ( 
.A(n_4595),
.Y(n_5123)
);

NAND2xp5_ASAP7_75t_L g5124 ( 
.A(n_4784),
.B(n_4204),
.Y(n_5124)
);

AOI22xp33_ASAP7_75t_L g5125 ( 
.A1(n_4568),
.A2(n_2757),
.B1(n_2570),
.B2(n_2571),
.Y(n_5125)
);

BUFx3_ASAP7_75t_L g5126 ( 
.A(n_4512),
.Y(n_5126)
);

HB1xp67_ASAP7_75t_L g5127 ( 
.A(n_4599),
.Y(n_5127)
);

AOI22xp5_ASAP7_75t_L g5128 ( 
.A1(n_4606),
.A2(n_2630),
.B1(n_2604),
.B2(n_1006),
.Y(n_5128)
);

NAND2xp5_ASAP7_75t_L g5129 ( 
.A(n_4695),
.B(n_4205),
.Y(n_5129)
);

BUFx8_ASAP7_75t_SL g5130 ( 
.A(n_4591),
.Y(n_5130)
);

NOR2xp33_ASAP7_75t_L g5131 ( 
.A(n_4637),
.B(n_1246),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_SL g5132 ( 
.A(n_4813),
.B(n_4399),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_4764),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_4768),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4780),
.Y(n_5135)
);

AOI22xp5_ASAP7_75t_L g5136 ( 
.A1(n_4800),
.A2(n_2630),
.B1(n_2604),
.B2(n_1007),
.Y(n_5136)
);

AND2x4_ASAP7_75t_L g5137 ( 
.A(n_4528),
.B(n_4207),
.Y(n_5137)
);

BUFx3_ASAP7_75t_L g5138 ( 
.A(n_4786),
.Y(n_5138)
);

INVx1_ASAP7_75t_L g5139 ( 
.A(n_4783),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_4485),
.B(n_1178),
.Y(n_5140)
);

AOI22xp5_ASAP7_75t_L g5141 ( 
.A1(n_4802),
.A2(n_4557),
.B1(n_4524),
.B2(n_4499),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_4784),
.B(n_4208),
.Y(n_5142)
);

NAND2xp5_ASAP7_75t_L g5143 ( 
.A(n_4662),
.B(n_4209),
.Y(n_5143)
);

OR2x4_ASAP7_75t_L g5144 ( 
.A(n_4822),
.B(n_4211),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_4796),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_SL g5146 ( 
.A(n_4671),
.B(n_4399),
.Y(n_5146)
);

AND2x6_ASAP7_75t_L g5147 ( 
.A(n_4845),
.B(n_4214),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4827),
.Y(n_5148)
);

CKINVDCx5p33_ASAP7_75t_R g5149 ( 
.A(n_4614),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4830),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4849),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_4665),
.B(n_4217),
.Y(n_5152)
);

BUFx12f_ASAP7_75t_L g5153 ( 
.A(n_4791),
.Y(n_5153)
);

NAND2xp5_ASAP7_75t_L g5154 ( 
.A(n_4738),
.B(n_4221),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_4860),
.Y(n_5155)
);

AOI22xp5_ASAP7_75t_L g5156 ( 
.A1(n_4499),
.A2(n_2604),
.B1(n_1010),
.B2(n_1016),
.Y(n_5156)
);

INVx3_ASAP7_75t_L g5157 ( 
.A(n_4867),
.Y(n_5157)
);

AND2x4_ASAP7_75t_L g5158 ( 
.A(n_4528),
.B(n_4551),
.Y(n_5158)
);

INVx1_ASAP7_75t_L g5159 ( 
.A(n_4446),
.Y(n_5159)
);

INVx1_ASAP7_75t_L g5160 ( 
.A(n_4487),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_4740),
.B(n_4222),
.Y(n_5161)
);

INVx2_ASAP7_75t_L g5162 ( 
.A(n_4696),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_4751),
.B(n_4223),
.Y(n_5163)
);

AND2x6_ASAP7_75t_L g5164 ( 
.A(n_4580),
.B(n_4229),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_4776),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_SL g5166 ( 
.A(n_4562),
.B(n_4399),
.Y(n_5166)
);

NOR2xp33_ASAP7_75t_L g5167 ( 
.A(n_4639),
.B(n_1250),
.Y(n_5167)
);

INVx1_ASAP7_75t_L g5168 ( 
.A(n_4781),
.Y(n_5168)
);

NAND2xp5_ASAP7_75t_L g5169 ( 
.A(n_4832),
.B(n_4234),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_SL g5170 ( 
.A(n_4466),
.B(n_4438),
.Y(n_5170)
);

BUFx3_ASAP7_75t_L g5171 ( 
.A(n_4576),
.Y(n_5171)
);

AOI22xp33_ASAP7_75t_L g5172 ( 
.A1(n_4453),
.A2(n_2570),
.B1(n_2571),
.B2(n_2509),
.Y(n_5172)
);

INVx2_ASAP7_75t_SL g5173 ( 
.A(n_4576),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_L g5174 ( 
.A(n_4523),
.B(n_4542),
.Y(n_5174)
);

AOI22xp33_ASAP7_75t_SL g5175 ( 
.A1(n_4812),
.A2(n_1220),
.B1(n_1178),
.B2(n_1034),
.Y(n_5175)
);

INVx3_ASAP7_75t_L g5176 ( 
.A(n_4867),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_SL g5177 ( 
.A(n_4466),
.B(n_4438),
.Y(n_5177)
);

AOI22xp5_ASAP7_75t_L g5178 ( 
.A1(n_4488),
.A2(n_1048),
.B1(n_1053),
.B2(n_1003),
.Y(n_5178)
);

INVx3_ASAP7_75t_L g5179 ( 
.A(n_4670),
.Y(n_5179)
);

BUFx4f_ASAP7_75t_L g5180 ( 
.A(n_4581),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_4697),
.Y(n_5181)
);

INVxp67_ASAP7_75t_SL g5182 ( 
.A(n_4672),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_L g5183 ( 
.A(n_4700),
.B(n_4241),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_4708),
.Y(n_5184)
);

BUFx3_ASAP7_75t_L g5185 ( 
.A(n_4581),
.Y(n_5185)
);

NAND2xp5_ASAP7_75t_L g5186 ( 
.A(n_4798),
.B(n_4243),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_4742),
.Y(n_5187)
);

BUFx12f_ASAP7_75t_L g5188 ( 
.A(n_4829),
.Y(n_5188)
);

NAND2xp5_ASAP7_75t_SL g5189 ( 
.A(n_4486),
.B(n_4438),
.Y(n_5189)
);

INVx2_ASAP7_75t_L g5190 ( 
.A(n_4797),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_4798),
.B(n_4245),
.Y(n_5191)
);

NAND2x1p5_ASAP7_75t_L g5192 ( 
.A(n_4689),
.B(n_3599),
.Y(n_5192)
);

OAI22xp5_ASAP7_75t_SL g5193 ( 
.A1(n_4570),
.A2(n_4453),
.B1(n_4493),
.B2(n_4771),
.Y(n_5193)
);

AOI22xp5_ASAP7_75t_L g5194 ( 
.A1(n_4531),
.A2(n_4493),
.B1(n_4508),
.B2(n_4500),
.Y(n_5194)
);

BUFx3_ASAP7_75t_L g5195 ( 
.A(n_4581),
.Y(n_5195)
);

NAND2xp5_ASAP7_75t_SL g5196 ( 
.A(n_4486),
.B(n_4438),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_4511),
.B(n_4718),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_4718),
.B(n_4246),
.Y(n_5198)
);

AOI21xp5_ASAP7_75t_L g5199 ( 
.A1(n_4644),
.A2(n_4244),
.B(n_4036),
.Y(n_5199)
);

INVx2_ASAP7_75t_L g5200 ( 
.A(n_4803),
.Y(n_5200)
);

INVx1_ASAP7_75t_L g5201 ( 
.A(n_4678),
.Y(n_5201)
);

NAND2xp5_ASAP7_75t_L g5202 ( 
.A(n_4578),
.B(n_4250),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_4578),
.B(n_4251),
.Y(n_5203)
);

INVx2_ASAP7_75t_SL g5204 ( 
.A(n_4660),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_4447),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4824),
.Y(n_5206)
);

NAND2xp5_ASAP7_75t_SL g5207 ( 
.A(n_4555),
.B(n_3574),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_4837),
.Y(n_5208)
);

INVx2_ASAP7_75t_L g5209 ( 
.A(n_4839),
.Y(n_5209)
);

HB1xp67_ASAP7_75t_L g5210 ( 
.A(n_4650),
.Y(n_5210)
);

INVx1_ASAP7_75t_L g5211 ( 
.A(n_4854),
.Y(n_5211)
);

BUFx3_ASAP7_75t_L g5212 ( 
.A(n_4857),
.Y(n_5212)
);

AOI22xp5_ASAP7_75t_L g5213 ( 
.A1(n_4500),
.A2(n_1071),
.B1(n_1077),
.B2(n_1058),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_4855),
.Y(n_5214)
);

NOR2xp33_ASAP7_75t_L g5215 ( 
.A(n_4596),
.B(n_1253),
.Y(n_5215)
);

NOR2xp33_ASAP7_75t_R g5216 ( 
.A(n_4733),
.B(n_3511),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_4858),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_4861),
.Y(n_5218)
);

AOI22xp5_ASAP7_75t_L g5219 ( 
.A1(n_4508),
.A2(n_1082),
.B1(n_1086),
.B2(n_1079),
.Y(n_5219)
);

NOR3xp33_ASAP7_75t_SL g5220 ( 
.A(n_4641),
.B(n_1094),
.C(n_1093),
.Y(n_5220)
);

HB1xp67_ASAP7_75t_L g5221 ( 
.A(n_4650),
.Y(n_5221)
);

NAND2xp5_ASAP7_75t_L g5222 ( 
.A(n_4744),
.B(n_4253),
.Y(n_5222)
);

INVx1_ASAP7_75t_L g5223 ( 
.A(n_4862),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_SL g5224 ( 
.A(n_4514),
.B(n_3574),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_4723),
.B(n_4259),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_4726),
.B(n_4262),
.Y(n_5226)
);

AOI22xp5_ASAP7_75t_L g5227 ( 
.A1(n_4807),
.A2(n_1103),
.B1(n_1110),
.B2(n_1095),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_4864),
.Y(n_5228)
);

AOI22xp33_ASAP7_75t_L g5229 ( 
.A1(n_4709),
.A2(n_2571),
.B1(n_2572),
.B2(n_2509),
.Y(n_5229)
);

NAND2xp5_ASAP7_75t_SL g5230 ( 
.A(n_4514),
.B(n_3574),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4626),
.B(n_4263),
.Y(n_5231)
);

BUFx3_ASAP7_75t_L g5232 ( 
.A(n_4857),
.Y(n_5232)
);

XNOR2xp5_ASAP7_75t_L g5233 ( 
.A(n_4778),
.B(n_1111),
.Y(n_5233)
);

NAND2xp5_ASAP7_75t_SL g5234 ( 
.A(n_4840),
.B(n_3574),
.Y(n_5234)
);

AND2x4_ASAP7_75t_L g5235 ( 
.A(n_4528),
.B(n_4264),
.Y(n_5235)
);

AOI22xp5_ASAP7_75t_L g5236 ( 
.A1(n_4677),
.A2(n_1127),
.B1(n_1138),
.B2(n_1122),
.Y(n_5236)
);

INVx2_ASAP7_75t_SL g5237 ( 
.A(n_4761),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_4501),
.B(n_4265),
.Y(n_5238)
);

NAND2xp33_ASAP7_75t_SL g5239 ( 
.A(n_4743),
.B(n_3833),
.Y(n_5239)
);

BUFx12f_ASAP7_75t_L g5240 ( 
.A(n_4757),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_4865),
.Y(n_5241)
);

OAI21xp5_ASAP7_75t_L g5242 ( 
.A1(n_4717),
.A2(n_4210),
.B(n_4231),
.Y(n_5242)
);

BUFx3_ASAP7_75t_L g5243 ( 
.A(n_4670),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_L g5244 ( 
.A(n_4547),
.B(n_4267),
.Y(n_5244)
);

INVx3_ASAP7_75t_L g5245 ( 
.A(n_4670),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_4866),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_SL g5247 ( 
.A(n_4663),
.B(n_4231),
.Y(n_5247)
);

INVx3_ASAP7_75t_L g5248 ( 
.A(n_4509),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_4868),
.Y(n_5249)
);

OR2x2_ASAP7_75t_L g5250 ( 
.A(n_4710),
.B(n_4268),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_4646),
.B(n_4269),
.Y(n_5251)
);

INVx1_ASAP7_75t_L g5252 ( 
.A(n_4869),
.Y(n_5252)
);

HB1xp67_ASAP7_75t_L g5253 ( 
.A(n_4712),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4750),
.Y(n_5254)
);

INVx1_ASAP7_75t_L g5255 ( 
.A(n_4545),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_4716),
.B(n_4275),
.Y(n_5256)
);

INVx3_ASAP7_75t_L g5257 ( 
.A(n_4509),
.Y(n_5257)
);

INVx2_ASAP7_75t_SL g5258 ( 
.A(n_4530),
.Y(n_5258)
);

AOI22xp33_ASAP7_75t_L g5259 ( 
.A1(n_4709),
.A2(n_4504),
.B1(n_4686),
.B2(n_4808),
.Y(n_5259)
);

INVx2_ASAP7_75t_L g5260 ( 
.A(n_4775),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_SL g5261 ( 
.A(n_4502),
.B(n_4770),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_4754),
.Y(n_5262)
);

INVx2_ASAP7_75t_L g5263 ( 
.A(n_4799),
.Y(n_5263)
);

AOI22xp5_ASAP7_75t_L g5264 ( 
.A1(n_4706),
.A2(n_1151),
.B1(n_1153),
.B2(n_1140),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_SL g5265 ( 
.A(n_4529),
.B(n_4237),
.Y(n_5265)
);

INVx5_ASAP7_75t_L g5266 ( 
.A(n_4551),
.Y(n_5266)
);

INVx2_ASAP7_75t_L g5267 ( 
.A(n_4748),
.Y(n_5267)
);

NOR2xp33_ASAP7_75t_L g5268 ( 
.A(n_4600),
.B(n_1260),
.Y(n_5268)
);

AOI21xp33_ASAP7_75t_L g5269 ( 
.A1(n_4517),
.A2(n_4266),
.B(n_4237),
.Y(n_5269)
);

NOR2xp33_ASAP7_75t_R g5270 ( 
.A(n_4495),
.B(n_3511),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_4746),
.B(n_4347),
.Y(n_5271)
);

A2O1A1Ixp33_ASAP7_75t_L g5272 ( 
.A1(n_4450),
.A2(n_4276),
.B(n_4278),
.C(n_4277),
.Y(n_5272)
);

A2O1A1Ixp33_ASAP7_75t_SL g5273 ( 
.A1(n_4766),
.A2(n_2748),
.B(n_2767),
.C(n_2759),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_4746),
.B(n_4362),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_SL g5275 ( 
.A(n_4450),
.B(n_4266),
.Y(n_5275)
);

AOI22xp33_ASAP7_75t_SL g5276 ( 
.A1(n_4765),
.A2(n_1220),
.B1(n_1178),
.B2(n_1164),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_4767),
.Y(n_5277)
);

BUFx4f_ASAP7_75t_L g5278 ( 
.A(n_4551),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_4772),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4789),
.Y(n_5280)
);

INVx2_ASAP7_75t_L g5281 ( 
.A(n_4731),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_4792),
.Y(n_5282)
);

INVx2_ASAP7_75t_L g5283 ( 
.A(n_4793),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4795),
.Y(n_5284)
);

NAND2xp5_ASAP7_75t_L g5285 ( 
.A(n_4686),
.B(n_4369),
.Y(n_5285)
);

NOR2xp33_ASAP7_75t_L g5286 ( 
.A(n_4602),
.B(n_1261),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_4579),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_4815),
.A2(n_4244),
.B(n_4036),
.Y(n_5288)
);

AND2x2_ASAP7_75t_L g5289 ( 
.A(n_4611),
.B(n_1220),
.Y(n_5289)
);

INVx1_ASAP7_75t_SL g5290 ( 
.A(n_4593),
.Y(n_5290)
);

AOI22xp33_ASAP7_75t_L g5291 ( 
.A1(n_4504),
.A2(n_4604),
.B1(n_4470),
.B2(n_4455),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_4607),
.B(n_1220),
.Y(n_5292)
);

BUFx2_ASAP7_75t_L g5293 ( 
.A(n_4530),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_4613),
.B(n_4280),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_4617),
.B(n_4281),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_4586),
.B(n_4283),
.Y(n_5296)
);

AND2x4_ASAP7_75t_L g5297 ( 
.A(n_4603),
.B(n_4284),
.Y(n_5297)
);

AND2x4_ASAP7_75t_L g5298 ( 
.A(n_4623),
.B(n_4286),
.Y(n_5298)
);

AO21x2_ASAP7_75t_L g5299 ( 
.A1(n_4825),
.A2(n_4442),
.B(n_3924),
.Y(n_5299)
);

AOI22xp33_ASAP7_75t_L g5300 ( 
.A1(n_4604),
.A2(n_2572),
.B1(n_2575),
.B2(n_2571),
.Y(n_5300)
);

BUFx10_ASAP7_75t_L g5301 ( 
.A(n_4608),
.Y(n_5301)
);

INVx2_ASAP7_75t_SL g5302 ( 
.A(n_4573),
.Y(n_5302)
);

HB1xp67_ASAP7_75t_L g5303 ( 
.A(n_4712),
.Y(n_5303)
);

HB1xp67_ASAP7_75t_L g5304 ( 
.A(n_4633),
.Y(n_5304)
);

OR2x6_ASAP7_75t_L g5305 ( 
.A(n_4790),
.B(n_4408),
.Y(n_5305)
);

BUFx6f_ASAP7_75t_L g5306 ( 
.A(n_4790),
.Y(n_5306)
);

INVx2_ASAP7_75t_L g5307 ( 
.A(n_4732),
.Y(n_5307)
);

INVx2_ASAP7_75t_L g5308 ( 
.A(n_4871),
.Y(n_5308)
);

INVx3_ASAP7_75t_L g5309 ( 
.A(n_5064),
.Y(n_5309)
);

BUFx3_ASAP7_75t_L g5310 ( 
.A(n_5073),
.Y(n_5310)
);

AOI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_4907),
.A2(n_4589),
.B(n_4782),
.Y(n_5311)
);

OR2x2_ASAP7_75t_L g5312 ( 
.A(n_4961),
.B(n_4983),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_5210),
.B(n_5221),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_4873),
.Y(n_5314)
);

AOI21xp5_ASAP7_75t_L g5315 ( 
.A1(n_5052),
.A2(n_4809),
.B(n_4774),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_4879),
.Y(n_5316)
);

AOI22x1_ASAP7_75t_L g5317 ( 
.A1(n_5293),
.A2(n_1165),
.B1(n_1168),
.B2(n_1157),
.Y(n_5317)
);

OAI21xp5_ASAP7_75t_L g5318 ( 
.A1(n_4890),
.A2(n_4653),
.B(n_4587),
.Y(n_5318)
);

AOI21xp5_ASAP7_75t_L g5319 ( 
.A1(n_5052),
.A2(n_4809),
.B(n_4774),
.Y(n_5319)
);

AOI21xp5_ASAP7_75t_L g5320 ( 
.A1(n_4964),
.A2(n_4821),
.B(n_4818),
.Y(n_5320)
);

OAI21xp5_ASAP7_75t_L g5321 ( 
.A1(n_4958),
.A2(n_4979),
.B(n_5032),
.Y(n_5321)
);

AOI21xp5_ASAP7_75t_L g5322 ( 
.A1(n_4964),
.A2(n_4836),
.B(n_4833),
.Y(n_5322)
);

NAND2x1p5_ASAP7_75t_L g5323 ( 
.A(n_4910),
.B(n_4661),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_4942),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_4877),
.B(n_4292),
.Y(n_5325)
);

AOI21x1_ASAP7_75t_L g5326 ( 
.A1(n_4932),
.A2(n_4693),
.B(n_4683),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_4960),
.Y(n_5327)
);

INVx3_ASAP7_75t_L g5328 ( 
.A(n_5064),
.Y(n_5328)
);

INVx1_ASAP7_75t_L g5329 ( 
.A(n_4967),
.Y(n_5329)
);

NAND2xp5_ASAP7_75t_L g5330 ( 
.A(n_5182),
.B(n_4293),
.Y(n_5330)
);

BUFx3_ASAP7_75t_L g5331 ( 
.A(n_5105),
.Y(n_5331)
);

A2O1A1Ixp33_ASAP7_75t_L g5332 ( 
.A1(n_4966),
.A2(n_4850),
.B(n_4669),
.C(n_4517),
.Y(n_5332)
);

O2A1O1Ixp33_ASAP7_75t_L g5333 ( 
.A1(n_5038),
.A2(n_4649),
.B(n_4474),
.C(n_4477),
.Y(n_5333)
);

AOI22x1_ASAP7_75t_L g5334 ( 
.A1(n_4997),
.A2(n_1169),
.B1(n_1175),
.B2(n_1166),
.Y(n_5334)
);

NAND2x1p5_ASAP7_75t_L g5335 ( 
.A(n_4910),
.B(n_4758),
.Y(n_5335)
);

BUFx6f_ASAP7_75t_L g5336 ( 
.A(n_5180),
.Y(n_5336)
);

OAI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_5131),
.A2(n_4656),
.B(n_4655),
.Y(n_5337)
);

AOI22xp5_ASAP7_75t_L g5338 ( 
.A1(n_5035),
.A2(n_4470),
.B1(n_4497),
.B2(n_4455),
.Y(n_5338)
);

CKINVDCx8_ASAP7_75t_R g5339 ( 
.A(n_4941),
.Y(n_5339)
);

AND2x2_ASAP7_75t_L g5340 ( 
.A(n_5103),
.B(n_4608),
.Y(n_5340)
);

O2A1O1Ixp5_ASAP7_75t_L g5341 ( 
.A1(n_5224),
.A2(n_4460),
.B(n_4472),
.C(n_4848),
.Y(n_5341)
);

NOR3xp33_ASAP7_75t_L g5342 ( 
.A(n_5001),
.B(n_1032),
.C(n_1009),
.Y(n_5342)
);

NOR3xp33_ASAP7_75t_L g5343 ( 
.A(n_4874),
.B(n_1033),
.C(n_1032),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_4933),
.B(n_4296),
.Y(n_5344)
);

HB1xp67_ASAP7_75t_L g5345 ( 
.A(n_4961),
.Y(n_5345)
);

AOI21xp5_ASAP7_75t_L g5346 ( 
.A1(n_5042),
.A2(n_5275),
.B(n_4936),
.Y(n_5346)
);

OAI21x1_ASAP7_75t_L g5347 ( 
.A1(n_5030),
.A2(n_5199),
.B(n_4717),
.Y(n_5347)
);

AOI21xp5_ASAP7_75t_L g5348 ( 
.A1(n_4921),
.A2(n_4841),
.B(n_4863),
.Y(n_5348)
);

AOI21xp5_ASAP7_75t_L g5349 ( 
.A1(n_5242),
.A2(n_4801),
.B(n_4348),
.Y(n_5349)
);

OAI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_5167),
.A2(n_4554),
.B(n_4550),
.Y(n_5350)
);

AOI21xp5_ASAP7_75t_L g5351 ( 
.A1(n_5242),
.A2(n_4801),
.B(n_4348),
.Y(n_5351)
);

NAND2xp5_ASAP7_75t_L g5352 ( 
.A(n_4937),
.B(n_4300),
.Y(n_5352)
);

NOR2xp33_ASAP7_75t_L g5353 ( 
.A(n_4969),
.B(n_4490),
.Y(n_5353)
);

O2A1O1Ixp33_ASAP7_75t_L g5354 ( 
.A1(n_4946),
.A2(n_1041),
.B(n_1051),
.C(n_1033),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_4884),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_5055),
.A2(n_4350),
.B(n_4295),
.Y(n_5356)
);

NOR2xp33_ASAP7_75t_L g5357 ( 
.A(n_5130),
.B(n_4569),
.Y(n_5357)
);

HB1xp67_ASAP7_75t_SL g5358 ( 
.A(n_4955),
.Y(n_5358)
);

OA22x2_ASAP7_75t_L g5359 ( 
.A1(n_5193),
.A2(n_4301),
.B1(n_4305),
.B2(n_4304),
.Y(n_5359)
);

NOR2xp33_ASAP7_75t_L g5360 ( 
.A(n_5005),
.B(n_4584),
.Y(n_5360)
);

AOI21xp5_ASAP7_75t_L g5361 ( 
.A1(n_5055),
.A2(n_4361),
.B(n_4350),
.Y(n_5361)
);

NOR2xp33_ASAP7_75t_SL g5362 ( 
.A(n_4910),
.B(n_4810),
.Y(n_5362)
);

OAI21xp5_ASAP7_75t_L g5363 ( 
.A1(n_5104),
.A2(n_4638),
.B(n_4619),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_SL g5364 ( 
.A(n_4917),
.B(n_4810),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_SL g5365 ( 
.A(n_4917),
.B(n_4810),
.Y(n_5365)
);

AOI21xp5_ASAP7_75t_L g5366 ( 
.A1(n_5040),
.A2(n_4361),
.B(n_4295),
.Y(n_5366)
);

AND2x2_ASAP7_75t_L g5367 ( 
.A(n_5127),
.B(n_4810),
.Y(n_5367)
);

NOR2xp33_ASAP7_75t_L g5368 ( 
.A(n_4965),
.B(n_4573),
.Y(n_5368)
);

AOI21xp5_ASAP7_75t_L g5369 ( 
.A1(n_5269),
.A2(n_3915),
.B(n_3818),
.Y(n_5369)
);

NAND2xp5_ASAP7_75t_L g5370 ( 
.A(n_5187),
.B(n_4306),
.Y(n_5370)
);

INVxp67_ASAP7_75t_L g5371 ( 
.A(n_4923),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_4973),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_5201),
.B(n_4310),
.Y(n_5373)
);

OR2x2_ASAP7_75t_L g5374 ( 
.A(n_4983),
.B(n_4804),
.Y(n_5374)
);

AOI21xp5_ASAP7_75t_L g5375 ( 
.A1(n_5269),
.A2(n_3915),
.B(n_3818),
.Y(n_5375)
);

OAI22xp5_ASAP7_75t_L g5376 ( 
.A1(n_4919),
.A2(n_4838),
.B1(n_4804),
.B2(n_4311),
.Y(n_5376)
);

AOI22xp33_ASAP7_75t_L g5377 ( 
.A1(n_5291),
.A2(n_4842),
.B1(n_4810),
.B2(n_2575),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_SL g5378 ( 
.A(n_5270),
.B(n_4810),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_5253),
.B(n_4312),
.Y(n_5379)
);

O2A1O1Ixp33_ASAP7_75t_L g5380 ( 
.A1(n_5273),
.A2(n_1060),
.B(n_1061),
.C(n_1041),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_4974),
.Y(n_5381)
);

AOI21x1_ASAP7_75t_L g5382 ( 
.A1(n_5014),
.A2(n_3832),
.B(n_3697),
.Y(n_5382)
);

AND2x2_ASAP7_75t_L g5383 ( 
.A(n_5303),
.B(n_4313),
.Y(n_5383)
);

NAND2xp5_ASAP7_75t_L g5384 ( 
.A(n_4993),
.B(n_4315),
.Y(n_5384)
);

NAND2xp5_ASAP7_75t_L g5385 ( 
.A(n_5198),
.B(n_4321),
.Y(n_5385)
);

OAI21xp5_ASAP7_75t_L g5386 ( 
.A1(n_5104),
.A2(n_4838),
.B(n_1060),
.Y(n_5386)
);

CKINVDCx5p33_ASAP7_75t_R g5387 ( 
.A(n_5058),
.Y(n_5387)
);

NOR2xp33_ASAP7_75t_L g5388 ( 
.A(n_5018),
.B(n_1262),
.Y(n_5388)
);

OAI21xp5_ASAP7_75t_L g5389 ( 
.A1(n_5067),
.A2(n_5053),
.B(n_4954),
.Y(n_5389)
);

INVx2_ASAP7_75t_L g5390 ( 
.A(n_4903),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5237),
.B(n_4894),
.Y(n_5391)
);

NAND2xp5_ASAP7_75t_L g5392 ( 
.A(n_5198),
.B(n_4323),
.Y(n_5392)
);

BUFx3_ASAP7_75t_L g5393 ( 
.A(n_4949),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_4985),
.B(n_4326),
.Y(n_5394)
);

NOR3xp33_ASAP7_75t_L g5395 ( 
.A(n_4870),
.B(n_1061),
.C(n_1051),
.Y(n_5395)
);

INVx2_ASAP7_75t_L g5396 ( 
.A(n_4922),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_L g5397 ( 
.A(n_4976),
.B(n_4327),
.Y(n_5397)
);

HB1xp67_ASAP7_75t_L g5398 ( 
.A(n_5026),
.Y(n_5398)
);

AND2x2_ASAP7_75t_L g5399 ( 
.A(n_4894),
.B(n_4329),
.Y(n_5399)
);

AOI21xp5_ASAP7_75t_L g5400 ( 
.A1(n_4901),
.A2(n_3915),
.B(n_3818),
.Y(n_5400)
);

OAI22xp5_ASAP7_75t_L g5401 ( 
.A1(n_5012),
.A2(n_4368),
.B1(n_4330),
.B2(n_4338),
.Y(n_5401)
);

A2O1A1Ixp33_ASAP7_75t_L g5402 ( 
.A1(n_5128),
.A2(n_1414),
.B(n_1415),
.C(n_1410),
.Y(n_5402)
);

NAND2xp5_ASAP7_75t_L g5403 ( 
.A(n_4976),
.B(n_4333),
.Y(n_5403)
);

NOR2xp33_ASAP7_75t_L g5404 ( 
.A(n_5101),
.B(n_1275),
.Y(n_5404)
);

NOR2xp33_ASAP7_75t_L g5405 ( 
.A(n_5078),
.B(n_1280),
.Y(n_5405)
);

OAI22xp5_ASAP7_75t_L g5406 ( 
.A1(n_5072),
.A2(n_4344),
.B1(n_4353),
.B2(n_4345),
.Y(n_5406)
);

HB1xp67_ASAP7_75t_L g5407 ( 
.A(n_4971),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_4987),
.Y(n_5408)
);

OAI22xp5_ASAP7_75t_L g5409 ( 
.A1(n_5141),
.A2(n_5095),
.B1(n_5087),
.B2(n_5156),
.Y(n_5409)
);

BUFx2_ASAP7_75t_L g5410 ( 
.A(n_4990),
.Y(n_5410)
);

NAND2xp5_ASAP7_75t_L g5411 ( 
.A(n_5165),
.B(n_4355),
.Y(n_5411)
);

OAI21xp5_ASAP7_75t_L g5412 ( 
.A1(n_4954),
.A2(n_1075),
.B(n_1066),
.Y(n_5412)
);

NAND2xp5_ASAP7_75t_SL g5413 ( 
.A(n_4953),
.B(n_5078),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_SL g5414 ( 
.A(n_4953),
.B(n_4689),
.Y(n_5414)
);

NAND2xp5_ASAP7_75t_L g5415 ( 
.A(n_5168),
.B(n_4356),
.Y(n_5415)
);

AOI21xp5_ASAP7_75t_L g5416 ( 
.A1(n_4901),
.A2(n_3915),
.B(n_3818),
.Y(n_5416)
);

AOI21xp5_ASAP7_75t_L g5417 ( 
.A1(n_4902),
.A2(n_3598),
.B(n_3561),
.Y(n_5417)
);

AND2x6_ASAP7_75t_L g5418 ( 
.A(n_5092),
.B(n_4735),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_4995),
.Y(n_5419)
);

BUFx12f_ASAP7_75t_L g5420 ( 
.A(n_4898),
.Y(n_5420)
);

OR2x6_ASAP7_75t_SL g5421 ( 
.A(n_5123),
.B(n_1177),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_4925),
.Y(n_5422)
);

AO32x1_ASAP7_75t_L g5423 ( 
.A1(n_5255),
.A2(n_4364),
.A3(n_4358),
.B1(n_3737),
.B2(n_3743),
.Y(n_5423)
);

OAI22xp5_ASAP7_75t_L g5424 ( 
.A1(n_5033),
.A2(n_4122),
.B1(n_3393),
.B2(n_3405),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_L g5425 ( 
.A(n_5254),
.B(n_4881),
.Y(n_5425)
);

AOI21xp5_ASAP7_75t_L g5426 ( 
.A1(n_4902),
.A2(n_3598),
.B(n_3561),
.Y(n_5426)
);

BUFx6f_ASAP7_75t_L g5427 ( 
.A(n_5180),
.Y(n_5427)
);

AND2x2_ASAP7_75t_L g5428 ( 
.A(n_4991),
.B(n_1066),
.Y(n_5428)
);

BUFx6f_ASAP7_75t_L g5429 ( 
.A(n_5113),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_SL g5430 ( 
.A(n_4915),
.B(n_4981),
.Y(n_5430)
);

OAI21x1_ASAP7_75t_L g5431 ( 
.A1(n_5234),
.A2(n_3832),
.B(n_3697),
.Y(n_5431)
);

O2A1O1Ixp33_ASAP7_75t_L g5432 ( 
.A1(n_4912),
.A2(n_1085),
.B(n_1099),
.C(n_1090),
.Y(n_5432)
);

AOI21xp5_ASAP7_75t_L g5433 ( 
.A1(n_5239),
.A2(n_3598),
.B(n_3561),
.Y(n_5433)
);

NAND2xp5_ASAP7_75t_L g5434 ( 
.A(n_4885),
.B(n_5190),
.Y(n_5434)
);

AOI21xp5_ASAP7_75t_L g5435 ( 
.A1(n_5132),
.A2(n_3642),
.B(n_3598),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_4928),
.Y(n_5436)
);

AOI22xp5_ASAP7_75t_L g5437 ( 
.A1(n_5091),
.A2(n_1085),
.B1(n_1090),
.B2(n_1075),
.Y(n_5437)
);

INVx2_ASAP7_75t_L g5438 ( 
.A(n_4930),
.Y(n_5438)
);

NOR2xp33_ASAP7_75t_L g5439 ( 
.A(n_5188),
.B(n_5065),
.Y(n_5439)
);

NAND2xp5_ASAP7_75t_L g5440 ( 
.A(n_5200),
.B(n_5209),
.Y(n_5440)
);

OAI22xp5_ASAP7_75t_L g5441 ( 
.A1(n_5033),
.A2(n_5136),
.B1(n_5194),
.B2(n_5193),
.Y(n_5441)
);

AOI21x1_ASAP7_75t_L g5442 ( 
.A1(n_5034),
.A2(n_1643),
.B(n_1642),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_L g5443 ( 
.A(n_5214),
.B(n_4735),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_4994),
.B(n_3912),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_4935),
.Y(n_5445)
);

AO21x1_ASAP7_75t_L g5446 ( 
.A1(n_5186),
.A2(n_1415),
.B(n_1414),
.Y(n_5446)
);

OAI21xp5_ASAP7_75t_L g5447 ( 
.A1(n_5264),
.A2(n_1107),
.B(n_1099),
.Y(n_5447)
);

AOI21xp5_ASAP7_75t_L g5448 ( 
.A1(n_5230),
.A2(n_3642),
.B(n_3598),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_4994),
.B(n_3912),
.Y(n_5449)
);

AOI21xp5_ASAP7_75t_L g5450 ( 
.A1(n_5093),
.A2(n_4893),
.B(n_5106),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_4996),
.B(n_3921),
.Y(n_5451)
);

OAI22xp5_ASAP7_75t_L g5452 ( 
.A1(n_5002),
.A2(n_4122),
.B1(n_3393),
.B2(n_3405),
.Y(n_5452)
);

O2A1O1Ixp33_ASAP7_75t_L g5453 ( 
.A1(n_5215),
.A2(n_1113),
.B(n_1120),
.C(n_1115),
.Y(n_5453)
);

OR2x6_ASAP7_75t_SL g5454 ( 
.A(n_5149),
.B(n_1183),
.Y(n_5454)
);

NAND2xp5_ASAP7_75t_L g5455 ( 
.A(n_4996),
.B(n_3921),
.Y(n_5455)
);

NOR2xp33_ASAP7_75t_SL g5456 ( 
.A(n_4970),
.B(n_4790),
.Y(n_5456)
);

INVx2_ASAP7_75t_L g5457 ( 
.A(n_4940),
.Y(n_5457)
);

AOI21xp5_ASAP7_75t_L g5458 ( 
.A1(n_4893),
.A2(n_3670),
.B(n_3642),
.Y(n_5458)
);

BUFx6f_ASAP7_75t_L g5459 ( 
.A(n_5113),
.Y(n_5459)
);

NOR2xp33_ASAP7_75t_L g5460 ( 
.A(n_4924),
.B(n_1282),
.Y(n_5460)
);

NOR2xp33_ASAP7_75t_L g5461 ( 
.A(n_5020),
.B(n_1284),
.Y(n_5461)
);

OR2x2_ASAP7_75t_L g5462 ( 
.A(n_5075),
.B(n_1648),
.Y(n_5462)
);

AOI21xp5_ASAP7_75t_L g5463 ( 
.A1(n_5288),
.A2(n_5272),
.B(n_5011),
.Y(n_5463)
);

NAND2xp5_ASAP7_75t_SL g5464 ( 
.A(n_4970),
.B(n_3857),
.Y(n_5464)
);

NOR3xp33_ASAP7_75t_L g5465 ( 
.A(n_4897),
.B(n_1113),
.C(n_1107),
.Y(n_5465)
);

NAND2xp5_ASAP7_75t_L g5466 ( 
.A(n_5011),
.B(n_3927),
.Y(n_5466)
);

OAI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_5091),
.A2(n_3393),
.B1(n_3405),
.B2(n_3383),
.Y(n_5467)
);

OAI21xp33_ASAP7_75t_SL g5468 ( 
.A1(n_4950),
.A2(n_1120),
.B(n_1115),
.Y(n_5468)
);

NAND2xp5_ASAP7_75t_L g5469 ( 
.A(n_5206),
.B(n_3927),
.Y(n_5469)
);

INVx8_ASAP7_75t_L g5470 ( 
.A(n_5164),
.Y(n_5470)
);

INVxp67_ASAP7_75t_L g5471 ( 
.A(n_5021),
.Y(n_5471)
);

AO21x1_ASAP7_75t_L g5472 ( 
.A1(n_5191),
.A2(n_1449),
.B(n_1421),
.Y(n_5472)
);

AOI21xp5_ASAP7_75t_L g5473 ( 
.A1(n_5143),
.A2(n_3670),
.B(n_3642),
.Y(n_5473)
);

AOI21xp5_ASAP7_75t_L g5474 ( 
.A1(n_5143),
.A2(n_5154),
.B(n_5152),
.Y(n_5474)
);

AOI22xp5_ASAP7_75t_L g5475 ( 
.A1(n_5259),
.A2(n_5098),
.B1(n_4999),
.B2(n_5233),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5004),
.Y(n_5476)
);

OAI21xp5_ASAP7_75t_L g5477 ( 
.A1(n_5268),
.A2(n_1125),
.B(n_1121),
.Y(n_5477)
);

HB1xp67_ASAP7_75t_L g5478 ( 
.A(n_4908),
.Y(n_5478)
);

AOI21xp5_ASAP7_75t_L g5479 ( 
.A1(n_5152),
.A2(n_3670),
.B(n_3642),
.Y(n_5479)
);

NAND2xp5_ASAP7_75t_L g5480 ( 
.A(n_5208),
.B(n_3930),
.Y(n_5480)
);

HB1xp67_ASAP7_75t_L g5481 ( 
.A(n_4908),
.Y(n_5481)
);

AOI22xp5_ASAP7_75t_L g5482 ( 
.A1(n_5197),
.A2(n_1125),
.B1(n_1128),
.B2(n_1121),
.Y(n_5482)
);

OAI21xp5_ASAP7_75t_L g5483 ( 
.A1(n_5286),
.A2(n_1137),
.B(n_1128),
.Y(n_5483)
);

NAND2xp5_ASAP7_75t_L g5484 ( 
.A(n_5211),
.B(n_3930),
.Y(n_5484)
);

NOR2xp33_ASAP7_75t_SL g5485 ( 
.A(n_4883),
.B(n_3700),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5007),
.Y(n_5486)
);

OAI22xp5_ASAP7_75t_L g5487 ( 
.A1(n_5178),
.A2(n_3393),
.B1(n_3405),
.B2(n_3383),
.Y(n_5487)
);

AOI21xp5_ASAP7_75t_L g5488 ( 
.A1(n_5154),
.A2(n_3670),
.B(n_3642),
.Y(n_5488)
);

AOI21xp5_ASAP7_75t_L g5489 ( 
.A1(n_5161),
.A2(n_3670),
.B(n_3437),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_5217),
.B(n_3934),
.Y(n_5490)
);

NAND2xp5_ASAP7_75t_L g5491 ( 
.A(n_5218),
.B(n_3934),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_SL g5492 ( 
.A(n_4970),
.B(n_3857),
.Y(n_5492)
);

NOR2xp33_ASAP7_75t_SL g5493 ( 
.A(n_5097),
.B(n_3760),
.Y(n_5493)
);

AOI22xp5_ASAP7_75t_L g5494 ( 
.A1(n_5197),
.A2(n_1145),
.B1(n_1146),
.B2(n_1137),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5010),
.Y(n_5495)
);

BUFx3_ASAP7_75t_L g5496 ( 
.A(n_5086),
.Y(n_5496)
);

HB1xp67_ASAP7_75t_L g5497 ( 
.A(n_4988),
.Y(n_5497)
);

AO21x1_ASAP7_75t_L g5498 ( 
.A1(n_5265),
.A2(n_1449),
.B(n_1421),
.Y(n_5498)
);

NOR2xp33_ASAP7_75t_SL g5499 ( 
.A(n_4883),
.B(n_3768),
.Y(n_5499)
);

NAND2xp5_ASAP7_75t_L g5500 ( 
.A(n_5223),
.B(n_1145),
.Y(n_5500)
);

OA22x2_ASAP7_75t_L g5501 ( 
.A1(n_5227),
.A2(n_1458),
.B1(n_1457),
.B2(n_1649),
.Y(n_5501)
);

NAND2x1p5_ASAP7_75t_L g5502 ( 
.A(n_5097),
.B(n_3926),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_5161),
.A2(n_3670),
.B(n_3437),
.Y(n_5503)
);

AOI21xp5_ASAP7_75t_L g5504 ( 
.A1(n_5044),
.A2(n_3388),
.B(n_3857),
.Y(n_5504)
);

NOR3xp33_ASAP7_75t_L g5505 ( 
.A(n_5166),
.B(n_1170),
.C(n_1146),
.Y(n_5505)
);

OR2x6_ASAP7_75t_L g5506 ( 
.A(n_4872),
.B(n_3737),
.Y(n_5506)
);

NAND2xp5_ASAP7_75t_L g5507 ( 
.A(n_5228),
.B(n_1170),
.Y(n_5507)
);

AND2x2_ASAP7_75t_L g5508 ( 
.A(n_4978),
.B(n_1221),
.Y(n_5508)
);

AOI21xp5_ASAP7_75t_L g5509 ( 
.A1(n_5278),
.A2(n_5080),
.B(n_5029),
.Y(n_5509)
);

INVx2_ASAP7_75t_L g5510 ( 
.A(n_4943),
.Y(n_5510)
);

AOI21xp5_ASAP7_75t_L g5511 ( 
.A1(n_5278),
.A2(n_3388),
.B(n_3857),
.Y(n_5511)
);

OAI21x1_ASAP7_75t_L g5512 ( 
.A1(n_5060),
.A2(n_3737),
.B(n_3738),
.Y(n_5512)
);

AOI21xp5_ASAP7_75t_L g5513 ( 
.A1(n_5029),
.A2(n_3916),
.B(n_3857),
.Y(n_5513)
);

OAI22xp5_ASAP7_75t_L g5514 ( 
.A1(n_5213),
.A2(n_3484),
.B1(n_3489),
.B2(n_3383),
.Y(n_5514)
);

NAND2xp5_ASAP7_75t_L g5515 ( 
.A(n_5241),
.B(n_1221),
.Y(n_5515)
);

NAND2xp5_ASAP7_75t_L g5516 ( 
.A(n_5246),
.B(n_1222),
.Y(n_5516)
);

BUFx2_ASAP7_75t_L g5517 ( 
.A(n_5144),
.Y(n_5517)
);

NAND2xp5_ASAP7_75t_L g5518 ( 
.A(n_5249),
.B(n_1222),
.Y(n_5518)
);

NAND2xp5_ASAP7_75t_SL g5519 ( 
.A(n_5097),
.B(n_3916),
.Y(n_5519)
);

INVxp67_ASAP7_75t_L g5520 ( 
.A(n_4916),
.Y(n_5520)
);

A2O1A1Ixp33_ASAP7_75t_SL g5521 ( 
.A1(n_5070),
.A2(n_1230),
.B(n_1235),
.C(n_1229),
.Y(n_5521)
);

NAND2xp5_ASAP7_75t_L g5522 ( 
.A(n_5252),
.B(n_1229),
.Y(n_5522)
);

NAND2xp5_ASAP7_75t_L g5523 ( 
.A(n_5013),
.B(n_1230),
.Y(n_5523)
);

BUFx4f_ASAP7_75t_L g5524 ( 
.A(n_5019),
.Y(n_5524)
);

INVx2_ASAP7_75t_L g5525 ( 
.A(n_4944),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5022),
.Y(n_5526)
);

OA22x2_ASAP7_75t_L g5527 ( 
.A1(n_4977),
.A2(n_1458),
.B1(n_1457),
.B2(n_1652),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_5023),
.B(n_1235),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_5023),
.B(n_1237),
.Y(n_5529)
);

OAI21xp33_ASAP7_75t_L g5530 ( 
.A1(n_5219),
.A2(n_990),
.B(n_952),
.Y(n_5530)
);

NAND2xp5_ASAP7_75t_L g5531 ( 
.A(n_5222),
.B(n_1237),
.Y(n_5531)
);

AOI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_5080),
.A2(n_3916),
.B(n_3585),
.Y(n_5532)
);

NAND2xp5_ASAP7_75t_L g5533 ( 
.A(n_5124),
.B(n_5142),
.Y(n_5533)
);

INVx5_ASAP7_75t_L g5534 ( 
.A(n_5120),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5028),
.Y(n_5535)
);

NAND2xp5_ASAP7_75t_L g5536 ( 
.A(n_5124),
.B(n_1245),
.Y(n_5536)
);

INVxp67_ASAP7_75t_L g5537 ( 
.A(n_5063),
.Y(n_5537)
);

NAND2xp5_ASAP7_75t_L g5538 ( 
.A(n_5142),
.B(n_1245),
.Y(n_5538)
);

OR2x6_ASAP7_75t_L g5539 ( 
.A(n_5305),
.B(n_3673),
.Y(n_5539)
);

INVx2_ASAP7_75t_L g5540 ( 
.A(n_4947),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5039),
.Y(n_5541)
);

INVx3_ASAP7_75t_L g5542 ( 
.A(n_5077),
.Y(n_5542)
);

INVx11_ASAP7_75t_L g5543 ( 
.A(n_5058),
.Y(n_5543)
);

NOR2xp33_ASAP7_75t_SL g5544 ( 
.A(n_5120),
.B(n_3768),
.Y(n_5544)
);

NAND2xp5_ASAP7_75t_L g5545 ( 
.A(n_5225),
.B(n_1252),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_L g5546 ( 
.A(n_5226),
.B(n_1252),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_4959),
.Y(n_5547)
);

AND2x2_ASAP7_75t_L g5548 ( 
.A(n_4978),
.B(n_1256),
.Y(n_5548)
);

INVxp67_ASAP7_75t_L g5549 ( 
.A(n_5089),
.Y(n_5549)
);

NAND2xp5_ASAP7_75t_L g5550 ( 
.A(n_5129),
.B(n_5183),
.Y(n_5550)
);

AOI22xp5_ASAP7_75t_L g5551 ( 
.A1(n_5172),
.A2(n_1265),
.B1(n_1271),
.B2(n_1256),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5041),
.Y(n_5552)
);

OAI21xp5_ASAP7_75t_L g5553 ( 
.A1(n_4957),
.A2(n_1271),
.B(n_1265),
.Y(n_5553)
);

AOI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_5085),
.A2(n_3916),
.B(n_3585),
.Y(n_5554)
);

A2O1A1Ixp33_ASAP7_75t_L g5555 ( 
.A1(n_5102),
.A2(n_1185),
.B(n_1193),
.C(n_1184),
.Y(n_5555)
);

AOI21xp33_ASAP7_75t_L g5556 ( 
.A1(n_5247),
.A2(n_3330),
.B(n_3363),
.Y(n_5556)
);

NOR3xp33_ASAP7_75t_L g5557 ( 
.A(n_5076),
.B(n_1276),
.C(n_1273),
.Y(n_5557)
);

NAND3xp33_ASAP7_75t_L g5558 ( 
.A(n_4980),
.B(n_1276),
.C(n_1273),
.Y(n_5558)
);

NOR2xp33_ASAP7_75t_L g5559 ( 
.A(n_4878),
.B(n_1291),
.Y(n_5559)
);

AOI21xp5_ASAP7_75t_L g5560 ( 
.A1(n_5085),
.A2(n_3916),
.B(n_3585),
.Y(n_5560)
);

AOI22xp33_ASAP7_75t_L g5561 ( 
.A1(n_4880),
.A2(n_5267),
.B1(n_5140),
.B2(n_5292),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_4962),
.Y(n_5562)
);

AOI21xp5_ASAP7_75t_L g5563 ( 
.A1(n_4900),
.A2(n_3586),
.B(n_3533),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_5000),
.B(n_1278),
.Y(n_5564)
);

INVx1_ASAP7_75t_L g5565 ( 
.A(n_5043),
.Y(n_5565)
);

AOI21xp5_ASAP7_75t_L g5566 ( 
.A1(n_4918),
.A2(n_3629),
.B(n_3586),
.Y(n_5566)
);

AND2x2_ASAP7_75t_L g5567 ( 
.A(n_5000),
.B(n_1278),
.Y(n_5567)
);

NAND3xp33_ASAP7_75t_L g5568 ( 
.A(n_5287),
.B(n_1321),
.C(n_1286),
.Y(n_5568)
);

CKINVDCx16_ASAP7_75t_R g5569 ( 
.A(n_4899),
.Y(n_5569)
);

AOI22xp5_ASAP7_75t_L g5570 ( 
.A1(n_5289),
.A2(n_1321),
.B1(n_1326),
.B2(n_1286),
.Y(n_5570)
);

OA21x2_ASAP7_75t_L g5571 ( 
.A1(n_5202),
.A2(n_3743),
.B(n_3738),
.Y(n_5571)
);

CKINVDCx10_ASAP7_75t_R g5572 ( 
.A(n_4914),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_SL g5573 ( 
.A(n_5120),
.B(n_5301),
.Y(n_5573)
);

NAND2xp5_ASAP7_75t_L g5574 ( 
.A(n_4982),
.B(n_1326),
.Y(n_5574)
);

AOI21xp5_ASAP7_75t_L g5575 ( 
.A1(n_5169),
.A2(n_3629),
.B(n_3586),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_5057),
.B(n_5262),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_5277),
.B(n_1332),
.Y(n_5577)
);

AOI21xp5_ASAP7_75t_L g5578 ( 
.A1(n_5169),
.A2(n_4892),
.B(n_4875),
.Y(n_5578)
);

BUFx2_ASAP7_75t_L g5579 ( 
.A(n_5144),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_5279),
.B(n_1332),
.Y(n_5580)
);

INVx2_ASAP7_75t_L g5581 ( 
.A(n_4963),
.Y(n_5581)
);

NAND2xp5_ASAP7_75t_SL g5582 ( 
.A(n_5301),
.B(n_3839),
.Y(n_5582)
);

AOI22xp33_ASAP7_75t_L g5583 ( 
.A1(n_5006),
.A2(n_2575),
.B1(n_2583),
.B2(n_2572),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5280),
.B(n_1340),
.Y(n_5584)
);

AOI22x1_ASAP7_75t_L g5585 ( 
.A1(n_5157),
.A2(n_1200),
.B1(n_1202),
.B2(n_1186),
.Y(n_5585)
);

AND2x2_ASAP7_75t_L g5586 ( 
.A(n_5138),
.B(n_1340),
.Y(n_5586)
);

AOI21x1_ASAP7_75t_L g5587 ( 
.A1(n_5261),
.A2(n_1654),
.B(n_1653),
.Y(n_5587)
);

NAND2xp5_ASAP7_75t_L g5588 ( 
.A(n_5282),
.B(n_1341),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_5045),
.Y(n_5589)
);

BUFx6f_ASAP7_75t_L g5590 ( 
.A(n_5113),
.Y(n_5590)
);

NAND2xp33_ASAP7_75t_SL g5591 ( 
.A(n_5017),
.B(n_3839),
.Y(n_5591)
);

AOI221xp5_ASAP7_75t_SL g5592 ( 
.A1(n_5108),
.A2(n_1357),
.B1(n_1372),
.B2(n_1355),
.C(n_1341),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5284),
.B(n_5205),
.Y(n_5593)
);

O2A1O1Ixp33_ASAP7_75t_L g5594 ( 
.A1(n_4975),
.A2(n_1357),
.B(n_1372),
.C(n_1355),
.Y(n_5594)
);

A2O1A1Ixp33_ASAP7_75t_L g5595 ( 
.A1(n_5220),
.A2(n_1210),
.B(n_1212),
.C(n_1198),
.Y(n_5595)
);

NAND2xp5_ASAP7_75t_L g5596 ( 
.A(n_5283),
.B(n_1381),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_5047),
.Y(n_5597)
);

NAND2xp5_ASAP7_75t_L g5598 ( 
.A(n_5251),
.B(n_5256),
.Y(n_5598)
);

AOI21xp5_ASAP7_75t_L g5599 ( 
.A1(n_4875),
.A2(n_3629),
.B(n_3586),
.Y(n_5599)
);

AND2x4_ASAP7_75t_L g5600 ( 
.A(n_5158),
.B(n_3673),
.Y(n_5600)
);

OAI22xp5_ASAP7_75t_L g5601 ( 
.A1(n_5236),
.A2(n_5110),
.B1(n_5056),
.B2(n_5294),
.Y(n_5601)
);

AND2x4_ASAP7_75t_L g5602 ( 
.A(n_5158),
.B(n_3673),
.Y(n_5602)
);

OAI21xp5_ASAP7_75t_L g5603 ( 
.A1(n_5296),
.A2(n_1384),
.B(n_1381),
.Y(n_5603)
);

AND2x2_ASAP7_75t_L g5604 ( 
.A(n_5077),
.B(n_1384),
.Y(n_5604)
);

CKINVDCx8_ASAP7_75t_R g5605 ( 
.A(n_4941),
.Y(n_5605)
);

NAND3xp33_ASAP7_75t_L g5606 ( 
.A(n_5174),
.B(n_1393),
.C(n_1385),
.Y(n_5606)
);

OAI21xp5_ASAP7_75t_L g5607 ( 
.A1(n_5079),
.A2(n_5082),
.B(n_5231),
.Y(n_5607)
);

NAND3xp33_ASAP7_75t_L g5608 ( 
.A(n_5174),
.B(n_1393),
.C(n_1385),
.Y(n_5608)
);

INVx2_ASAP7_75t_L g5609 ( 
.A(n_4986),
.Y(n_5609)
);

AND2x4_ASAP7_75t_L g5610 ( 
.A(n_5266),
.B(n_3783),
.Y(n_5610)
);

BUFx6f_ASAP7_75t_L g5611 ( 
.A(n_4896),
.Y(n_5611)
);

AOI21xp5_ASAP7_75t_L g5612 ( 
.A1(n_4892),
.A2(n_3629),
.B(n_3604),
.Y(n_5612)
);

INVx2_ASAP7_75t_L g5613 ( 
.A(n_4989),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_SL g5614 ( 
.A(n_5059),
.B(n_3839),
.Y(n_5614)
);

A2O1A1Ixp33_ASAP7_75t_L g5615 ( 
.A1(n_5271),
.A2(n_1226),
.B(n_1232),
.C(n_1227),
.Y(n_5615)
);

AOI22x1_ASAP7_75t_L g5616 ( 
.A1(n_5157),
.A2(n_1233),
.B1(n_1238),
.B2(n_1234),
.Y(n_5616)
);

NAND2xp5_ASAP7_75t_L g5617 ( 
.A(n_5244),
.B(n_5238),
.Y(n_5617)
);

O2A1O1Ixp33_ASAP7_75t_L g5618 ( 
.A1(n_5295),
.A2(n_1401),
.B(n_1413),
.C(n_1397),
.Y(n_5618)
);

A2O1A1Ixp33_ASAP7_75t_L g5619 ( 
.A1(n_5271),
.A2(n_1242),
.B(n_1247),
.C(n_1244),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_5015),
.B(n_1397),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5163),
.B(n_1401),
.Y(n_5621)
);

BUFx6f_ASAP7_75t_L g5622 ( 
.A(n_4896),
.Y(n_5622)
);

NOR2xp33_ASAP7_75t_SL g5623 ( 
.A(n_5083),
.B(n_5266),
.Y(n_5623)
);

NAND2xp5_ASAP7_75t_SL g5624 ( 
.A(n_5059),
.B(n_4891),
.Y(n_5624)
);

OA22x2_ASAP7_75t_L g5625 ( 
.A1(n_5008),
.A2(n_1657),
.B1(n_1655),
.B2(n_2559),
.Y(n_5625)
);

O2A1O1Ixp33_ASAP7_75t_SL g5626 ( 
.A1(n_4911),
.A2(n_1417),
.B(n_1419),
.C(n_1413),
.Y(n_5626)
);

INVx11_ASAP7_75t_L g5627 ( 
.A(n_5119),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_5048),
.Y(n_5628)
);

AOI21xp5_ASAP7_75t_L g5629 ( 
.A1(n_5066),
.A2(n_3604),
.B(n_3582),
.Y(n_5629)
);

AOI21xp5_ASAP7_75t_L g5630 ( 
.A1(n_5146),
.A2(n_3609),
.B(n_3582),
.Y(n_5630)
);

BUFx2_ASAP7_75t_L g5631 ( 
.A(n_5121),
.Y(n_5631)
);

AND2x4_ASAP7_75t_L g5632 ( 
.A(n_5266),
.B(n_3783),
.Y(n_5632)
);

BUFx12f_ASAP7_75t_L g5633 ( 
.A(n_5119),
.Y(n_5633)
);

BUFx2_ASAP7_75t_L g5634 ( 
.A(n_5240),
.Y(n_5634)
);

NOR2xp33_ASAP7_75t_L g5635 ( 
.A(n_5062),
.B(n_1298),
.Y(n_5635)
);

INVx2_ASAP7_75t_L g5636 ( 
.A(n_4992),
.Y(n_5636)
);

AOI21xp5_ASAP7_75t_L g5637 ( 
.A1(n_4938),
.A2(n_3609),
.B(n_3839),
.Y(n_5637)
);

AOI21xp5_ASAP7_75t_L g5638 ( 
.A1(n_5305),
.A2(n_3886),
.B(n_3871),
.Y(n_5638)
);

NAND2xp5_ASAP7_75t_L g5639 ( 
.A(n_5163),
.B(n_1417),
.Y(n_5639)
);

NOR2xp33_ASAP7_75t_L g5640 ( 
.A(n_5126),
.B(n_1300),
.Y(n_5640)
);

OAI21x1_ASAP7_75t_L g5641 ( 
.A1(n_5060),
.A2(n_3842),
.B(n_3838),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_5054),
.B(n_1419),
.Y(n_5642)
);

NAND2x1p5_ASAP7_75t_L g5643 ( 
.A(n_5092),
.B(n_3783),
.Y(n_5643)
);

NAND2xp5_ASAP7_75t_L g5644 ( 
.A(n_5069),
.B(n_1426),
.Y(n_5644)
);

INVx1_ASAP7_75t_L g5645 ( 
.A(n_5071),
.Y(n_5645)
);

NOR2xp33_ASAP7_75t_L g5646 ( 
.A(n_5094),
.B(n_1304),
.Y(n_5646)
);

AOI21xp5_ASAP7_75t_L g5647 ( 
.A1(n_5305),
.A2(n_3886),
.B(n_3871),
.Y(n_5647)
);

A2O1A1Ixp33_ASAP7_75t_L g5648 ( 
.A1(n_5274),
.A2(n_1248),
.B(n_1281),
.C(n_1268),
.Y(n_5648)
);

AOI22xp33_ASAP7_75t_L g5649 ( 
.A1(n_5006),
.A2(n_2575),
.B1(n_2583),
.B2(n_2572),
.Y(n_5649)
);

AOI21xp5_ASAP7_75t_L g5650 ( 
.A1(n_5170),
.A2(n_3886),
.B(n_3871),
.Y(n_5650)
);

AOI21xp5_ASAP7_75t_L g5651 ( 
.A1(n_5177),
.A2(n_3886),
.B(n_3871),
.Y(n_5651)
);

O2A1O1Ixp33_ASAP7_75t_L g5652 ( 
.A1(n_5207),
.A2(n_1428),
.B(n_1429),
.C(n_1426),
.Y(n_5652)
);

AND2x2_ASAP7_75t_L g5653 ( 
.A(n_5137),
.B(n_1428),
.Y(n_5653)
);

AO21x1_ASAP7_75t_L g5654 ( 
.A1(n_5297),
.A2(n_1431),
.B(n_1429),
.Y(n_5654)
);

NOR2xp33_ASAP7_75t_L g5655 ( 
.A(n_5107),
.B(n_1311),
.Y(n_5655)
);

AOI22xp33_ASAP7_75t_L g5656 ( 
.A1(n_5006),
.A2(n_5202),
.B1(n_5285),
.B2(n_5203),
.Y(n_5656)
);

CKINVDCx10_ASAP7_75t_R g5657 ( 
.A(n_5118),
.Y(n_5657)
);

AOI21xp5_ASAP7_75t_L g5658 ( 
.A1(n_5189),
.A2(n_3922),
.B(n_3889),
.Y(n_5658)
);

AOI21xp5_ASAP7_75t_L g5659 ( 
.A1(n_5196),
.A2(n_3922),
.B(n_3889),
.Y(n_5659)
);

AOI21xp5_ASAP7_75t_L g5660 ( 
.A1(n_5088),
.A2(n_3922),
.B(n_3889),
.Y(n_5660)
);

AOI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_4972),
.A2(n_3922),
.B(n_3889),
.Y(n_5661)
);

NAND2xp5_ASAP7_75t_L g5662 ( 
.A(n_5074),
.B(n_1431),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_5016),
.Y(n_5663)
);

NAND2xp5_ASAP7_75t_L g5664 ( 
.A(n_5081),
.B(n_1444),
.Y(n_5664)
);

NAND2xp5_ASAP7_75t_L g5665 ( 
.A(n_5084),
.B(n_1444),
.Y(n_5665)
);

BUFx6f_ASAP7_75t_L g5666 ( 
.A(n_4896),
.Y(n_5666)
);

INVx2_ASAP7_75t_L g5667 ( 
.A(n_5024),
.Y(n_5667)
);

AOI21xp5_ASAP7_75t_L g5668 ( 
.A1(n_5009),
.A2(n_3411),
.B(n_3389),
.Y(n_5668)
);

AOI21xp5_ASAP7_75t_L g5669 ( 
.A1(n_5050),
.A2(n_3411),
.B(n_3389),
.Y(n_5669)
);

AOI22xp33_ASAP7_75t_L g5670 ( 
.A1(n_5006),
.A2(n_2601),
.B1(n_2628),
.B2(n_2583),
.Y(n_5670)
);

NAND2xp5_ASAP7_75t_L g5671 ( 
.A(n_5090),
.B(n_1454),
.Y(n_5671)
);

AO32x1_ASAP7_75t_L g5672 ( 
.A1(n_5307),
.A2(n_3843),
.A3(n_3842),
.B1(n_3838),
.B2(n_3862),
.Y(n_5672)
);

NOR2xp33_ASAP7_75t_SL g5673 ( 
.A(n_5164),
.B(n_3807),
.Y(n_5673)
);

INVx1_ASAP7_75t_L g5674 ( 
.A(n_5096),
.Y(n_5674)
);

NAND2xp5_ASAP7_75t_SL g5675 ( 
.A(n_4909),
.B(n_3383),
.Y(n_5675)
);

NAND3xp33_ASAP7_75t_L g5676 ( 
.A(n_5281),
.B(n_1461),
.C(n_1454),
.Y(n_5676)
);

NAND2xp5_ASAP7_75t_L g5677 ( 
.A(n_5099),
.B(n_1461),
.Y(n_5677)
);

AO22x1_ASAP7_75t_L g5678 ( 
.A1(n_5164),
.A2(n_1462),
.B1(n_1004),
.B2(n_1027),
.Y(n_5678)
);

AOI21xp5_ASAP7_75t_L g5679 ( 
.A1(n_5137),
.A2(n_3411),
.B(n_3389),
.Y(n_5679)
);

AOI21xp5_ASAP7_75t_L g5680 ( 
.A1(n_5235),
.A2(n_3411),
.B(n_3389),
.Y(n_5680)
);

OR2x2_ASAP7_75t_L g5681 ( 
.A(n_5100),
.B(n_1462),
.Y(n_5681)
);

NAND2xp5_ASAP7_75t_L g5682 ( 
.A(n_5109),
.B(n_1224),
.Y(n_5682)
);

INVxp67_ASAP7_75t_L g5683 ( 
.A(n_5304),
.Y(n_5683)
);

AO32x1_ASAP7_75t_L g5684 ( 
.A1(n_5260),
.A2(n_5263),
.A3(n_5302),
.B1(n_5258),
.B2(n_5116),
.Y(n_5684)
);

NOR3xp33_ASAP7_75t_L g5685 ( 
.A(n_5175),
.B(n_1027),
.C(n_1022),
.Y(n_5685)
);

NAND2xp5_ASAP7_75t_L g5686 ( 
.A(n_5114),
.B(n_1283),
.Y(n_5686)
);

A2O1A1Ixp33_ASAP7_75t_L g5687 ( 
.A1(n_5274),
.A2(n_1292),
.B(n_1293),
.C(n_1290),
.Y(n_5687)
);

OAI22xp5_ASAP7_75t_L g5688 ( 
.A1(n_5125),
.A2(n_3489),
.B1(n_3521),
.B2(n_3484),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_5115),
.Y(n_5689)
);

NOR2xp33_ASAP7_75t_L g5690 ( 
.A(n_5003),
.B(n_1313),
.Y(n_5690)
);

AOI22xp5_ASAP7_75t_L g5691 ( 
.A1(n_5147),
.A2(n_1439),
.B1(n_1423),
.B2(n_1297),
.Y(n_5691)
);

AOI21xp5_ASAP7_75t_L g5692 ( 
.A1(n_5235),
.A2(n_3488),
.B(n_3425),
.Y(n_5692)
);

AND2x2_ASAP7_75t_L g5693 ( 
.A(n_4888),
.B(n_1004),
.Y(n_5693)
);

AOI22xp5_ASAP7_75t_L g5694 ( 
.A1(n_5147),
.A2(n_1350),
.B1(n_1399),
.B2(n_1338),
.Y(n_5694)
);

AOI21xp5_ASAP7_75t_L g5695 ( 
.A1(n_5112),
.A2(n_3488),
.B(n_3425),
.Y(n_5695)
);

AND2x2_ASAP7_75t_L g5696 ( 
.A(n_4888),
.B(n_1004),
.Y(n_5696)
);

CKINVDCx20_ASAP7_75t_R g5697 ( 
.A(n_4904),
.Y(n_5697)
);

NAND2xp5_ASAP7_75t_L g5698 ( 
.A(n_5122),
.B(n_1294),
.Y(n_5698)
);

OAI21x1_ASAP7_75t_L g5699 ( 
.A1(n_5176),
.A2(n_3843),
.B(n_3862),
.Y(n_5699)
);

OR2x2_ASAP7_75t_L g5700 ( 
.A(n_5133),
.B(n_1022),
.Y(n_5700)
);

AO22x1_ASAP7_75t_L g5701 ( 
.A1(n_5164),
.A2(n_5204),
.B1(n_5019),
.B2(n_5147),
.Y(n_5701)
);

AOI21xp5_ASAP7_75t_L g5702 ( 
.A1(n_5299),
.A2(n_3488),
.B(n_3425),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_5027),
.Y(n_5703)
);

AOI21xp5_ASAP7_75t_L g5704 ( 
.A1(n_5299),
.A2(n_3488),
.B(n_3425),
.Y(n_5704)
);

OA22x2_ASAP7_75t_L g5705 ( 
.A1(n_5117),
.A2(n_2769),
.B1(n_2772),
.B2(n_2768),
.Y(n_5705)
);

NAND3xp33_ASAP7_75t_L g5706 ( 
.A(n_5297),
.B(n_1027),
.C(n_1022),
.Y(n_5706)
);

AND2x2_ASAP7_75t_L g5707 ( 
.A(n_5159),
.B(n_1037),
.Y(n_5707)
);

AO21x1_ASAP7_75t_L g5708 ( 
.A1(n_5298),
.A2(n_1049),
.B(n_1037),
.Y(n_5708)
);

AOI21xp5_ASAP7_75t_L g5709 ( 
.A1(n_4909),
.A2(n_4956),
.B(n_4939),
.Y(n_5709)
);

AOI21xp5_ASAP7_75t_L g5710 ( 
.A1(n_4939),
.A2(n_3658),
.B(n_3645),
.Y(n_5710)
);

NOR2xp33_ASAP7_75t_L g5711 ( 
.A(n_5036),
.B(n_1315),
.Y(n_5711)
);

AOI221xp5_ASAP7_75t_L g5712 ( 
.A1(n_5276),
.A2(n_1322),
.B1(n_1333),
.B2(n_1309),
.C(n_1307),
.Y(n_5712)
);

AOI21xp5_ASAP7_75t_L g5713 ( 
.A1(n_4956),
.A2(n_3658),
.B(n_3645),
.Y(n_5713)
);

OAI22xp5_ASAP7_75t_L g5714 ( 
.A1(n_5046),
.A2(n_3489),
.B1(n_3521),
.B2(n_3484),
.Y(n_5714)
);

OAI22x1_ASAP7_75t_L g5715 ( 
.A1(n_5160),
.A2(n_1344),
.B1(n_1348),
.B2(n_1339),
.Y(n_5715)
);

BUFx6f_ASAP7_75t_L g5716 ( 
.A(n_4931),
.Y(n_5716)
);

OAI22xp5_ASAP7_75t_L g5717 ( 
.A1(n_5229),
.A2(n_3489),
.B1(n_3521),
.B2(n_3484),
.Y(n_5717)
);

OAI21x1_ASAP7_75t_L g5718 ( 
.A1(n_5176),
.A2(n_3872),
.B(n_3866),
.Y(n_5718)
);

NAND2xp5_ASAP7_75t_SL g5719 ( 
.A(n_5025),
.B(n_3521),
.Y(n_5719)
);

NAND2xp5_ASAP7_75t_L g5720 ( 
.A(n_5134),
.B(n_1354),
.Y(n_5720)
);

OAI22xp5_ASAP7_75t_L g5721 ( 
.A1(n_5250),
.A2(n_3531),
.B1(n_3558),
.B2(n_3529),
.Y(n_5721)
);

NOR3xp33_ASAP7_75t_L g5722 ( 
.A(n_5179),
.B(n_1054),
.C(n_1049),
.Y(n_5722)
);

CKINVDCx8_ASAP7_75t_R g5723 ( 
.A(n_5037),
.Y(n_5723)
);

AOI22xp33_ASAP7_75t_SL g5724 ( 
.A1(n_5147),
.A2(n_1363),
.B1(n_1364),
.B2(n_1359),
.Y(n_5724)
);

NAND2xp5_ASAP7_75t_SL g5725 ( 
.A(n_5025),
.B(n_3529),
.Y(n_5725)
);

INVx3_ASAP7_75t_L g5726 ( 
.A(n_5212),
.Y(n_5726)
);

NAND2xp5_ASAP7_75t_L g5727 ( 
.A(n_5135),
.B(n_1374),
.Y(n_5727)
);

NAND2xp5_ASAP7_75t_L g5728 ( 
.A(n_5139),
.B(n_1379),
.Y(n_5728)
);

NOR2xp33_ASAP7_75t_SL g5729 ( 
.A(n_5019),
.B(n_3807),
.Y(n_5729)
);

AOI22xp5_ASAP7_75t_L g5730 ( 
.A1(n_5298),
.A2(n_1438),
.B1(n_1383),
.B2(n_1388),
.Y(n_5730)
);

INVx4_ASAP7_75t_L g5731 ( 
.A(n_5179),
.Y(n_5731)
);

NAND2xp5_ASAP7_75t_SL g5732 ( 
.A(n_4931),
.B(n_4968),
.Y(n_5732)
);

NAND2x1p5_ASAP7_75t_L g5733 ( 
.A(n_5306),
.B(n_3898),
.Y(n_5733)
);

AOI21xp5_ASAP7_75t_L g5734 ( 
.A1(n_5290),
.A2(n_3759),
.B(n_3688),
.Y(n_5734)
);

A2O1A1Ixp33_ASAP7_75t_L g5735 ( 
.A1(n_5203),
.A2(n_1389),
.B(n_1404),
.C(n_1380),
.Y(n_5735)
);

AOI21xp5_ASAP7_75t_L g5736 ( 
.A1(n_5290),
.A2(n_3759),
.B(n_3688),
.Y(n_5736)
);

INVx1_ASAP7_75t_L g5737 ( 
.A(n_5145),
.Y(n_5737)
);

NAND2xp5_ASAP7_75t_L g5738 ( 
.A(n_5148),
.B(n_1416),
.Y(n_5738)
);

NAND2xp5_ASAP7_75t_L g5739 ( 
.A(n_5150),
.B(n_1435),
.Y(n_5739)
);

NAND2xp5_ASAP7_75t_L g5740 ( 
.A(n_5151),
.B(n_1436),
.Y(n_5740)
);

NAND2xp5_ASAP7_75t_L g5741 ( 
.A(n_5155),
.B(n_1441),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5031),
.Y(n_5742)
);

AOI21xp5_ASAP7_75t_L g5743 ( 
.A1(n_5285),
.A2(n_3859),
.B(n_3801),
.Y(n_5743)
);

AOI21xp5_ASAP7_75t_L g5744 ( 
.A1(n_5117),
.A2(n_3859),
.B(n_3801),
.Y(n_5744)
);

INVx1_ASAP7_75t_SL g5745 ( 
.A(n_5153),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_4876),
.Y(n_5746)
);

A2O1A1Ixp33_ASAP7_75t_L g5747 ( 
.A1(n_4913),
.A2(n_1445),
.B(n_1456),
.C(n_1450),
.Y(n_5747)
);

NAND2xp5_ASAP7_75t_L g5748 ( 
.A(n_4887),
.B(n_4889),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5049),
.Y(n_5749)
);

AOI21xp5_ASAP7_75t_L g5750 ( 
.A1(n_5245),
.A2(n_3925),
.B(n_3874),
.Y(n_5750)
);

AOI21x1_ASAP7_75t_L g5751 ( 
.A1(n_5173),
.A2(n_3330),
.B(n_3866),
.Y(n_5751)
);

O2A1O1Ixp33_ASAP7_75t_SL g5752 ( 
.A1(n_5068),
.A2(n_1049),
.B(n_1054),
.C(n_1037),
.Y(n_5752)
);

AOI21xp5_ASAP7_75t_L g5753 ( 
.A1(n_5245),
.A2(n_3925),
.B(n_3874),
.Y(n_5753)
);

OAI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_4882),
.A2(n_1191),
.B(n_1054),
.Y(n_5754)
);

AOI21x1_ASAP7_75t_L g5755 ( 
.A1(n_4895),
.A2(n_3873),
.B(n_3872),
.Y(n_5755)
);

AOI21x1_ASAP7_75t_L g5756 ( 
.A1(n_4905),
.A2(n_4920),
.B(n_4906),
.Y(n_5756)
);

BUFx6f_ASAP7_75t_L g5757 ( 
.A(n_4931),
.Y(n_5757)
);

AND2x2_ASAP7_75t_L g5758 ( 
.A(n_5243),
.B(n_1191),
.Y(n_5758)
);

BUFx2_ASAP7_75t_L g5759 ( 
.A(n_5232),
.Y(n_5759)
);

INVx1_ASAP7_75t_L g5760 ( 
.A(n_5327),
.Y(n_5760)
);

AND2x2_ASAP7_75t_L g5761 ( 
.A(n_5497),
.B(n_5068),
.Y(n_5761)
);

BUFx3_ASAP7_75t_L g5762 ( 
.A(n_5331),
.Y(n_5762)
);

AND2x2_ASAP7_75t_L g5763 ( 
.A(n_5398),
.B(n_4952),
.Y(n_5763)
);

OR2x2_ASAP7_75t_L g5764 ( 
.A(n_5312),
.B(n_4926),
.Y(n_5764)
);

OAI21xp5_ASAP7_75t_L g5765 ( 
.A1(n_5321),
.A2(n_5300),
.B(n_1236),
.Y(n_5765)
);

INVxp67_ASAP7_75t_L g5766 ( 
.A(n_5407),
.Y(n_5766)
);

AOI21x1_ASAP7_75t_L g5767 ( 
.A1(n_5413),
.A2(n_4929),
.B(n_4927),
.Y(n_5767)
);

BUFx2_ASAP7_75t_L g5768 ( 
.A(n_5345),
.Y(n_5768)
);

NAND2xp5_ASAP7_75t_L g5769 ( 
.A(n_5478),
.B(n_4934),
.Y(n_5769)
);

CKINVDCx5p33_ASAP7_75t_R g5770 ( 
.A(n_5572),
.Y(n_5770)
);

OAI21x1_ASAP7_75t_L g5771 ( 
.A1(n_5347),
.A2(n_4886),
.B(n_5111),
.Y(n_5771)
);

AO21x2_ASAP7_75t_L g5772 ( 
.A1(n_5751),
.A2(n_5694),
.B(n_5691),
.Y(n_5772)
);

OAI21xp5_ASAP7_75t_L g5773 ( 
.A1(n_5691),
.A2(n_1236),
.B(n_1191),
.Y(n_5773)
);

AOI21xp5_ASAP7_75t_L g5774 ( 
.A1(n_5311),
.A2(n_3885),
.B(n_3807),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5329),
.Y(n_5775)
);

OAI21x1_ASAP7_75t_L g5776 ( 
.A1(n_5346),
.A2(n_4886),
.B(n_5111),
.Y(n_5776)
);

AOI21xp33_ASAP7_75t_L g5777 ( 
.A1(n_5441),
.A2(n_4948),
.B(n_4945),
.Y(n_5777)
);

AOI21xp5_ASAP7_75t_L g5778 ( 
.A1(n_5356),
.A2(n_3898),
.B(n_3885),
.Y(n_5778)
);

OAI21x1_ASAP7_75t_L g5779 ( 
.A1(n_5315),
.A2(n_5192),
.B(n_4951),
.Y(n_5779)
);

NAND2xp5_ASAP7_75t_L g5780 ( 
.A(n_5481),
.B(n_4952),
.Y(n_5780)
);

INVx2_ASAP7_75t_L g5781 ( 
.A(n_5746),
.Y(n_5781)
);

O2A1O1Ixp33_ASAP7_75t_L g5782 ( 
.A1(n_5389),
.A2(n_1455),
.B(n_1254),
.C(n_1285),
.Y(n_5782)
);

AOI21xp5_ASAP7_75t_L g5783 ( 
.A1(n_5361),
.A2(n_3898),
.B(n_3885),
.Y(n_5783)
);

NOR2xp33_ASAP7_75t_L g5784 ( 
.A(n_5393),
.B(n_5037),
.Y(n_5784)
);

AOI21xp5_ASAP7_75t_L g5785 ( 
.A1(n_5463),
.A2(n_3926),
.B(n_3632),
.Y(n_5785)
);

AOI21xp5_ASAP7_75t_L g5786 ( 
.A1(n_5450),
.A2(n_3926),
.B(n_3632),
.Y(n_5786)
);

AOI221xp5_ASAP7_75t_L g5787 ( 
.A1(n_5453),
.A2(n_1464),
.B1(n_1467),
.B2(n_1460),
.C(n_1442),
.Y(n_5787)
);

OAI21x1_ASAP7_75t_L g5788 ( 
.A1(n_5319),
.A2(n_5192),
.B(n_5248),
.Y(n_5788)
);

NOR2x1_ASAP7_75t_L g5789 ( 
.A(n_5410),
.B(n_5171),
.Y(n_5789)
);

AOI21x1_ASAP7_75t_L g5790 ( 
.A1(n_5701),
.A2(n_5184),
.B(n_5181),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5372),
.Y(n_5791)
);

AO31x2_ASAP7_75t_L g5792 ( 
.A1(n_5349),
.A2(n_5061),
.A3(n_5162),
.B(n_5051),
.Y(n_5792)
);

NAND2x1p5_ASAP7_75t_L g5793 ( 
.A(n_5534),
.B(n_5306),
.Y(n_5793)
);

A2O1A1Ixp33_ASAP7_75t_L g5794 ( 
.A1(n_5694),
.A2(n_1254),
.B(n_1285),
.C(n_1236),
.Y(n_5794)
);

NAND2xp5_ASAP7_75t_L g5795 ( 
.A(n_5533),
.B(n_4998),
.Y(n_5795)
);

BUFx6f_ASAP7_75t_L g5796 ( 
.A(n_5336),
.Y(n_5796)
);

AOI21xp5_ASAP7_75t_L g5797 ( 
.A1(n_5433),
.A2(n_3632),
.B(n_3599),
.Y(n_5797)
);

A2O1A1Ixp33_ASAP7_75t_L g5798 ( 
.A1(n_5332),
.A2(n_1285),
.B(n_1347),
.C(n_1254),
.Y(n_5798)
);

OR2x6_ASAP7_75t_L g5799 ( 
.A(n_5470),
.B(n_5306),
.Y(n_5799)
);

AOI21xp5_ASAP7_75t_L g5800 ( 
.A1(n_5366),
.A2(n_3599),
.B(n_3671),
.Y(n_5800)
);

AOI22xp33_ASAP7_75t_L g5801 ( 
.A1(n_5359),
.A2(n_5338),
.B1(n_5475),
.B2(n_5625),
.Y(n_5801)
);

OAI21x1_ASAP7_75t_L g5802 ( 
.A1(n_5369),
.A2(n_5257),
.B(n_5248),
.Y(n_5802)
);

NOR2xp33_ASAP7_75t_SL g5803 ( 
.A(n_5673),
.B(n_5185),
.Y(n_5803)
);

OAI21xp33_ASAP7_75t_SL g5804 ( 
.A1(n_5414),
.A2(n_1386),
.B(n_1347),
.Y(n_5804)
);

NOR2x1_ASAP7_75t_SL g5805 ( 
.A(n_5506),
.B(n_5195),
.Y(n_5805)
);

OAI21x1_ASAP7_75t_L g5806 ( 
.A1(n_5375),
.A2(n_5257),
.B(n_4998),
.Y(n_5806)
);

AOI21xp5_ASAP7_75t_L g5807 ( 
.A1(n_5673),
.A2(n_3928),
.B(n_3923),
.Y(n_5807)
);

AOI21xp5_ASAP7_75t_L g5808 ( 
.A1(n_5351),
.A2(n_3928),
.B(n_3923),
.Y(n_5808)
);

AOI21xp5_ASAP7_75t_L g5809 ( 
.A1(n_5354),
.A2(n_3928),
.B(n_3923),
.Y(n_5809)
);

AOI21xp33_ASAP7_75t_L g5810 ( 
.A1(n_5594),
.A2(n_4984),
.B(n_4968),
.Y(n_5810)
);

OAI21xp5_ASAP7_75t_L g5811 ( 
.A1(n_5558),
.A2(n_1386),
.B(n_1347),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_5702),
.A2(n_3876),
.B(n_3873),
.Y(n_5812)
);

AOI21xp5_ASAP7_75t_L g5813 ( 
.A1(n_5458),
.A2(n_3928),
.B(n_3923),
.Y(n_5813)
);

O2A1O1Ixp5_ASAP7_75t_L g5814 ( 
.A1(n_5477),
.A2(n_1455),
.B(n_1386),
.C(n_1911),
.Y(n_5814)
);

CKINVDCx5p33_ASAP7_75t_R g5815 ( 
.A(n_5657),
.Y(n_5815)
);

INVx2_ASAP7_75t_L g5816 ( 
.A(n_5308),
.Y(n_5816)
);

AOI221x1_ASAP7_75t_L g5817 ( 
.A1(n_5601),
.A2(n_1455),
.B1(n_4984),
.B2(n_4968),
.C(n_1274),
.Y(n_5817)
);

INVx2_ASAP7_75t_L g5818 ( 
.A(n_5314),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5355),
.Y(n_5819)
);

INVxp67_ASAP7_75t_L g5820 ( 
.A(n_5313),
.Y(n_5820)
);

NAND2xp5_ASAP7_75t_L g5821 ( 
.A(n_5474),
.B(n_4984),
.Y(n_5821)
);

AOI21xp5_ASAP7_75t_L g5822 ( 
.A1(n_5417),
.A2(n_3680),
.B(n_3671),
.Y(n_5822)
);

INVx2_ASAP7_75t_SL g5823 ( 
.A(n_5310),
.Y(n_5823)
);

AOI21xp5_ASAP7_75t_L g5824 ( 
.A1(n_5426),
.A2(n_3680),
.B(n_3671),
.Y(n_5824)
);

AO31x2_ASAP7_75t_L g5825 ( 
.A1(n_5708),
.A2(n_3879),
.A3(n_3876),
.B(n_3804),
.Y(n_5825)
);

INVx1_ASAP7_75t_L g5826 ( 
.A(n_5381),
.Y(n_5826)
);

OAI21xp5_ASAP7_75t_L g5827 ( 
.A1(n_5558),
.A2(n_3315),
.B(n_3311),
.Y(n_5827)
);

A2O1A1Ixp33_ASAP7_75t_L g5828 ( 
.A1(n_5483),
.A2(n_1318),
.B(n_1320),
.C(n_1317),
.Y(n_5828)
);

AOI21x1_ASAP7_75t_L g5829 ( 
.A1(n_5678),
.A2(n_1931),
.B(n_1911),
.Y(n_5829)
);

OAI21x1_ASAP7_75t_L g5830 ( 
.A1(n_5704),
.A2(n_3879),
.B(n_3680),
.Y(n_5830)
);

OAI21x1_ASAP7_75t_SL g5831 ( 
.A1(n_5607),
.A2(n_2777),
.B(n_2775),
.Y(n_5831)
);

AND2x2_ASAP7_75t_L g5832 ( 
.A(n_5340),
.B(n_5216),
.Y(n_5832)
);

OAI21xp5_ASAP7_75t_L g5833 ( 
.A1(n_5724),
.A2(n_3316),
.B(n_3315),
.Y(n_5833)
);

AOI21xp5_ASAP7_75t_L g5834 ( 
.A1(n_5623),
.A2(n_3887),
.B(n_3680),
.Y(n_5834)
);

OAI22xp5_ASAP7_75t_L g5835 ( 
.A1(n_5338),
.A2(n_1201),
.B1(n_1274),
.B2(n_991),
.Y(n_5835)
);

AOI21x1_ASAP7_75t_L g5836 ( 
.A1(n_5621),
.A2(n_1975),
.B(n_1931),
.Y(n_5836)
);

OAI21x1_ASAP7_75t_L g5837 ( 
.A1(n_5400),
.A2(n_3707),
.B(n_3671),
.Y(n_5837)
);

NOR2x1_ASAP7_75t_L g5838 ( 
.A(n_5394),
.B(n_3529),
.Y(n_5838)
);

OAI21xp5_ASAP7_75t_L g5839 ( 
.A1(n_5468),
.A2(n_3318),
.B(n_3316),
.Y(n_5839)
);

AOI21xp5_ASAP7_75t_L g5840 ( 
.A1(n_5623),
.A2(n_3714),
.B(n_3707),
.Y(n_5840)
);

OAI22x1_ASAP7_75t_L g5841 ( 
.A1(n_5517),
.A2(n_1324),
.B1(n_1325),
.B2(n_1323),
.Y(n_5841)
);

NAND2xp5_ASAP7_75t_SL g5842 ( 
.A(n_5509),
.B(n_2913),
.Y(n_5842)
);

OAI21x1_ASAP7_75t_L g5843 ( 
.A1(n_5416),
.A2(n_3714),
.B(n_3707),
.Y(n_5843)
);

AOI21xp5_ASAP7_75t_L g5844 ( 
.A1(n_5409),
.A2(n_3714),
.B(n_3707),
.Y(n_5844)
);

NAND2xp5_ASAP7_75t_L g5845 ( 
.A(n_5598),
.B(n_5550),
.Y(n_5845)
);

BUFx2_ASAP7_75t_L g5846 ( 
.A(n_5537),
.Y(n_5846)
);

AOI21xp5_ASAP7_75t_L g5847 ( 
.A1(n_5473),
.A2(n_3742),
.B(n_3714),
.Y(n_5847)
);

OAI21x1_ASAP7_75t_L g5848 ( 
.A1(n_5513),
.A2(n_3777),
.B(n_3742),
.Y(n_5848)
);

AO31x2_ASAP7_75t_L g5849 ( 
.A1(n_5401),
.A2(n_3804),
.A3(n_3810),
.B(n_3802),
.Y(n_5849)
);

INVx2_ASAP7_75t_SL g5850 ( 
.A(n_5496),
.Y(n_5850)
);

NOR2xp33_ASAP7_75t_SL g5851 ( 
.A(n_5470),
.B(n_3511),
.Y(n_5851)
);

OAI21x1_ASAP7_75t_L g5852 ( 
.A1(n_5583),
.A2(n_3777),
.B(n_3742),
.Y(n_5852)
);

INVx2_ASAP7_75t_SL g5853 ( 
.A(n_5543),
.Y(n_5853)
);

AOI21x1_ASAP7_75t_L g5854 ( 
.A1(n_5639),
.A2(n_5538),
.B(n_5536),
.Y(n_5854)
);

INVx3_ASAP7_75t_L g5855 ( 
.A(n_5309),
.Y(n_5855)
);

OAI21xp5_ASAP7_75t_L g5856 ( 
.A1(n_5606),
.A2(n_3322),
.B(n_3318),
.Y(n_5856)
);

NOR2xp33_ASAP7_75t_L g5857 ( 
.A(n_5421),
.B(n_342),
.Y(n_5857)
);

OAI21xp33_ASAP7_75t_SL g5858 ( 
.A1(n_5656),
.A2(n_3777),
.B(n_3742),
.Y(n_5858)
);

O2A1O1Ixp5_ASAP7_75t_L g5859 ( 
.A1(n_5624),
.A2(n_1991),
.B(n_1975),
.C(n_3529),
.Y(n_5859)
);

NAND2xp5_ASAP7_75t_SL g5860 ( 
.A(n_5631),
.B(n_2914),
.Y(n_5860)
);

NAND2xp5_ASAP7_75t_L g5861 ( 
.A(n_5383),
.B(n_991),
.Y(n_5861)
);

AND2x2_ASAP7_75t_L g5862 ( 
.A(n_5371),
.B(n_1201),
.Y(n_5862)
);

OAI21x1_ASAP7_75t_L g5863 ( 
.A1(n_5649),
.A2(n_3887),
.B(n_3865),
.Y(n_5863)
);

AOI21xp5_ASAP7_75t_L g5864 ( 
.A1(n_5479),
.A2(n_3887),
.B(n_3865),
.Y(n_5864)
);

AOI21x1_ASAP7_75t_L g5865 ( 
.A1(n_5528),
.A2(n_5529),
.B(n_5642),
.Y(n_5865)
);

BUFx2_ASAP7_75t_L g5866 ( 
.A(n_5683),
.Y(n_5866)
);

OAI21x1_ASAP7_75t_L g5867 ( 
.A1(n_5670),
.A2(n_3887),
.B(n_3865),
.Y(n_5867)
);

NAND2xp5_ASAP7_75t_L g5868 ( 
.A(n_5425),
.B(n_5617),
.Y(n_5868)
);

OAI21x1_ASAP7_75t_L g5869 ( 
.A1(n_5382),
.A2(n_3865),
.B(n_3777),
.Y(n_5869)
);

AOI21xp33_ASAP7_75t_L g5870 ( 
.A1(n_5592),
.A2(n_1274),
.B(n_1201),
.Y(n_5870)
);

CKINVDCx11_ASAP7_75t_R g5871 ( 
.A(n_5697),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_5408),
.Y(n_5872)
);

AOI21xp5_ASAP7_75t_L g5873 ( 
.A1(n_5488),
.A2(n_3877),
.B(n_3558),
.Y(n_5873)
);

AOI21xp5_ASAP7_75t_L g5874 ( 
.A1(n_5591),
.A2(n_3877),
.B(n_3558),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5419),
.Y(n_5875)
);

AOI21x1_ASAP7_75t_SL g5876 ( 
.A1(n_5428),
.A2(n_5686),
.B(n_5682),
.Y(n_5876)
);

AND2x2_ASAP7_75t_L g5877 ( 
.A(n_5471),
.B(n_1201),
.Y(n_5877)
);

NAND2xp5_ASAP7_75t_L g5878 ( 
.A(n_5576),
.B(n_1201),
.Y(n_5878)
);

AOI21xp5_ASAP7_75t_L g5879 ( 
.A1(n_5435),
.A2(n_3877),
.B(n_3558),
.Y(n_5879)
);

AOI21xp5_ASAP7_75t_L g5880 ( 
.A1(n_5489),
.A2(n_3877),
.B(n_3569),
.Y(n_5880)
);

BUFx6f_ASAP7_75t_L g5881 ( 
.A(n_5336),
.Y(n_5881)
);

AOI21xp5_ASAP7_75t_L g5882 ( 
.A1(n_5503),
.A2(n_3569),
.B(n_3531),
.Y(n_5882)
);

INVx2_ASAP7_75t_L g5883 ( 
.A(n_5390),
.Y(n_5883)
);

BUFx2_ASAP7_75t_L g5884 ( 
.A(n_5759),
.Y(n_5884)
);

NAND2xp5_ASAP7_75t_L g5885 ( 
.A(n_5578),
.B(n_1201),
.Y(n_5885)
);

NAND2xp5_ASAP7_75t_L g5886 ( 
.A(n_5344),
.B(n_5352),
.Y(n_5886)
);

BUFx2_ASAP7_75t_L g5887 ( 
.A(n_5579),
.Y(n_5887)
);

INVx1_ASAP7_75t_L g5888 ( 
.A(n_5476),
.Y(n_5888)
);

INVx3_ASAP7_75t_L g5889 ( 
.A(n_5309),
.Y(n_5889)
);

AOI21xp5_ASAP7_75t_L g5890 ( 
.A1(n_5599),
.A2(n_3569),
.B(n_3531),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5486),
.Y(n_5891)
);

AOI21xp5_ASAP7_75t_L g5892 ( 
.A1(n_5493),
.A2(n_3569),
.B(n_3531),
.Y(n_5892)
);

A2O1A1Ixp33_ASAP7_75t_L g5893 ( 
.A1(n_5475),
.A2(n_1328),
.B(n_1329),
.C(n_1327),
.Y(n_5893)
);

AO31x2_ASAP7_75t_L g5894 ( 
.A1(n_5406),
.A2(n_3804),
.A3(n_3810),
.B(n_3802),
.Y(n_5894)
);

AOI221x1_ASAP7_75t_L g5895 ( 
.A1(n_5318),
.A2(n_1337),
.B1(n_1443),
.B2(n_1274),
.C(n_1201),
.Y(n_5895)
);

A2O1A1Ixp33_ASAP7_75t_L g5896 ( 
.A1(n_5461),
.A2(n_5437),
.B(n_5618),
.C(n_5530),
.Y(n_5896)
);

OAI21x1_ASAP7_75t_L g5897 ( 
.A1(n_5431),
.A2(n_3618),
.B(n_3584),
.Y(n_5897)
);

INVx2_ASAP7_75t_L g5898 ( 
.A(n_5396),
.Y(n_5898)
);

NAND2xp5_ASAP7_75t_SL g5899 ( 
.A(n_5429),
.B(n_5459),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5495),
.Y(n_5900)
);

OAI21x1_ASAP7_75t_L g5901 ( 
.A1(n_5699),
.A2(n_3618),
.B(n_3584),
.Y(n_5901)
);

INVx3_ASAP7_75t_L g5902 ( 
.A(n_5328),
.Y(n_5902)
);

AOI221xp5_ASAP7_75t_SL g5903 ( 
.A1(n_5337),
.A2(n_1443),
.B1(n_1337),
.B2(n_1274),
.C(n_7),
.Y(n_5903)
);

AO21x1_ASAP7_75t_L g5904 ( 
.A1(n_5553),
.A2(n_1739),
.B(n_1737),
.Y(n_5904)
);

AOI21xp5_ASAP7_75t_L g5905 ( 
.A1(n_5493),
.A2(n_3618),
.B(n_3584),
.Y(n_5905)
);

AOI21xp5_ASAP7_75t_L g5906 ( 
.A1(n_5575),
.A2(n_3618),
.B(n_3584),
.Y(n_5906)
);

NOR2xp67_ASAP7_75t_L g5907 ( 
.A(n_5534),
.B(n_3633),
.Y(n_5907)
);

BUFx6f_ASAP7_75t_L g5908 ( 
.A(n_5336),
.Y(n_5908)
);

INVx2_ASAP7_75t_L g5909 ( 
.A(n_5422),
.Y(n_5909)
);

INVxp67_ASAP7_75t_SL g5910 ( 
.A(n_5330),
.Y(n_5910)
);

OAI21x1_ASAP7_75t_L g5911 ( 
.A1(n_5718),
.A2(n_3633),
.B(n_3802),
.Y(n_5911)
);

OAI21xp5_ASAP7_75t_L g5912 ( 
.A1(n_5606),
.A2(n_3327),
.B(n_3322),
.Y(n_5912)
);

OAI21x1_ASAP7_75t_L g5913 ( 
.A1(n_5532),
.A2(n_3633),
.B(n_3810),
.Y(n_5913)
);

NAND2xp33_ASAP7_75t_L g5914 ( 
.A(n_5387),
.B(n_1274),
.Y(n_5914)
);

NOR2x1_ASAP7_75t_L g5915 ( 
.A(n_5325),
.B(n_3633),
.Y(n_5915)
);

INVxp67_ASAP7_75t_SL g5916 ( 
.A(n_5434),
.Y(n_5916)
);

NAND2xp5_ASAP7_75t_L g5917 ( 
.A(n_5397),
.B(n_1274),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5436),
.Y(n_5918)
);

NAND2xp5_ASAP7_75t_L g5919 ( 
.A(n_5403),
.B(n_1337),
.Y(n_5919)
);

AOI21xp5_ASAP7_75t_L g5920 ( 
.A1(n_5362),
.A2(n_3648),
.B(n_3646),
.Y(n_5920)
);

OAI21x1_ASAP7_75t_L g5921 ( 
.A1(n_5554),
.A2(n_3815),
.B(n_3814),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5438),
.Y(n_5922)
);

INVx4_ASAP7_75t_L g5923 ( 
.A(n_5470),
.Y(n_5923)
);

AOI21x1_ASAP7_75t_SL g5924 ( 
.A1(n_5698),
.A2(n_5),
.B(n_6),
.Y(n_5924)
);

BUFx5_ASAP7_75t_L g5925 ( 
.A(n_5418),
.Y(n_5925)
);

OAI21x1_ASAP7_75t_L g5926 ( 
.A1(n_5560),
.A2(n_3815),
.B(n_3814),
.Y(n_5926)
);

A2O1A1Ixp33_ASAP7_75t_L g5927 ( 
.A1(n_5437),
.A2(n_1334),
.B(n_1336),
.C(n_1330),
.Y(n_5927)
);

OAI21x1_ASAP7_75t_L g5928 ( 
.A1(n_5743),
.A2(n_3815),
.B(n_3814),
.Y(n_5928)
);

NAND2xp5_ASAP7_75t_L g5929 ( 
.A(n_5379),
.B(n_5384),
.Y(n_5929)
);

OAI21x1_ASAP7_75t_L g5930 ( 
.A1(n_5326),
.A2(n_3824),
.B(n_3819),
.Y(n_5930)
);

NAND3xp33_ASAP7_75t_SL g5931 ( 
.A(n_5339),
.B(n_1343),
.C(n_1335),
.Y(n_5931)
);

OAI21x1_ASAP7_75t_L g5932 ( 
.A1(n_5442),
.A2(n_3851),
.B(n_3850),
.Y(n_5932)
);

OAI22xp5_ASAP7_75t_L g5933 ( 
.A1(n_5730),
.A2(n_1443),
.B1(n_1337),
.B2(n_1349),
.Y(n_5933)
);

HB1xp67_ASAP7_75t_L g5934 ( 
.A(n_5316),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5526),
.Y(n_5935)
);

AOI21xp5_ASAP7_75t_L g5936 ( 
.A1(n_5362),
.A2(n_3648),
.B(n_3646),
.Y(n_5936)
);

AO31x2_ASAP7_75t_L g5937 ( 
.A1(n_5446),
.A2(n_5472),
.A3(n_5376),
.B(n_5721),
.Y(n_5937)
);

OAI21xp5_ASAP7_75t_L g5938 ( 
.A1(n_5608),
.A2(n_3329),
.B(n_3327),
.Y(n_5938)
);

AOI21xp5_ASAP7_75t_L g5939 ( 
.A1(n_5448),
.A2(n_3648),
.B(n_3646),
.Y(n_5939)
);

AOI21xp5_ASAP7_75t_L g5940 ( 
.A1(n_5464),
.A2(n_3648),
.B(n_3646),
.Y(n_5940)
);

NAND2xp5_ASAP7_75t_L g5941 ( 
.A(n_5324),
.B(n_5385),
.Y(n_5941)
);

INVx1_ASAP7_75t_L g5942 ( 
.A(n_5535),
.Y(n_5942)
);

NAND2xp5_ASAP7_75t_SL g5943 ( 
.A(n_5429),
.B(n_2914),
.Y(n_5943)
);

NAND2xp5_ASAP7_75t_L g5944 ( 
.A(n_5392),
.B(n_1337),
.Y(n_5944)
);

OAI21x1_ASAP7_75t_L g5945 ( 
.A1(n_5638),
.A2(n_3824),
.B(n_3819),
.Y(n_5945)
);

NAND2xp5_ASAP7_75t_L g5946 ( 
.A(n_5541),
.B(n_1337),
.Y(n_5946)
);

OAI22xp5_ASAP7_75t_L g5947 ( 
.A1(n_5730),
.A2(n_1443),
.B1(n_1337),
.B2(n_1353),
.Y(n_5947)
);

AND2x2_ASAP7_75t_L g5948 ( 
.A(n_5391),
.B(n_1443),
.Y(n_5948)
);

NAND2x1p5_ASAP7_75t_L g5949 ( 
.A(n_5534),
.B(n_3555),
.Y(n_5949)
);

OAI21xp5_ASAP7_75t_L g5950 ( 
.A1(n_5608),
.A2(n_5412),
.B(n_5592),
.Y(n_5950)
);

INVx2_ASAP7_75t_L g5951 ( 
.A(n_5445),
.Y(n_5951)
);

OAI21xp5_ASAP7_75t_L g5952 ( 
.A1(n_5615),
.A2(n_3331),
.B(n_3329),
.Y(n_5952)
);

BUFx6f_ASAP7_75t_L g5953 ( 
.A(n_5427),
.Y(n_5953)
);

NAND3xp33_ASAP7_75t_L g5954 ( 
.A(n_5343),
.B(n_1443),
.C(n_1366),
.Y(n_5954)
);

OAI21x1_ASAP7_75t_L g5955 ( 
.A1(n_5647),
.A2(n_3824),
.B(n_3819),
.Y(n_5955)
);

INVx2_ASAP7_75t_L g5956 ( 
.A(n_5457),
.Y(n_5956)
);

NAND2xp5_ASAP7_75t_L g5957 ( 
.A(n_5552),
.B(n_1443),
.Y(n_5957)
);

NAND2xp5_ASAP7_75t_L g5958 ( 
.A(n_5565),
.B(n_6),
.Y(n_5958)
);

INVx2_ASAP7_75t_L g5959 ( 
.A(n_5510),
.Y(n_5959)
);

OAI21xp33_ASAP7_75t_L g5960 ( 
.A1(n_5619),
.A2(n_1368),
.B(n_1345),
.Y(n_5960)
);

AOI21x1_ASAP7_75t_L g5961 ( 
.A1(n_5644),
.A2(n_1991),
.B(n_1640),
.Y(n_5961)
);

OAI21x1_ASAP7_75t_L g5962 ( 
.A1(n_5587),
.A2(n_5512),
.B(n_5641),
.Y(n_5962)
);

AOI21xp5_ASAP7_75t_L g5963 ( 
.A1(n_5492),
.A2(n_3657),
.B(n_3546),
.Y(n_5963)
);

OAI21x1_ASAP7_75t_L g5964 ( 
.A1(n_5320),
.A2(n_3850),
.B(n_3846),
.Y(n_5964)
);

HB1xp67_ASAP7_75t_L g5965 ( 
.A(n_5589),
.Y(n_5965)
);

NAND2x1_ASAP7_75t_L g5966 ( 
.A(n_5328),
.B(n_3324),
.Y(n_5966)
);

AOI22xp5_ASAP7_75t_L g5967 ( 
.A1(n_5530),
.A2(n_1373),
.B1(n_1375),
.B2(n_1369),
.Y(n_5967)
);

INVx1_ASAP7_75t_SL g5968 ( 
.A(n_5726),
.Y(n_5968)
);

A2O1A1Ixp33_ASAP7_75t_L g5969 ( 
.A1(n_5648),
.A2(n_1391),
.B(n_1392),
.C(n_1387),
.Y(n_5969)
);

INVx5_ASAP7_75t_L g5970 ( 
.A(n_5506),
.Y(n_5970)
);

AND2x2_ASAP7_75t_SL g5971 ( 
.A(n_5569),
.B(n_3363),
.Y(n_5971)
);

AOI21xp33_ASAP7_75t_L g5972 ( 
.A1(n_5521),
.A2(n_2778),
.B(n_3331),
.Y(n_5972)
);

NOR2x1_ASAP7_75t_L g5973 ( 
.A(n_5731),
.B(n_3555),
.Y(n_5973)
);

AOI21xp5_ASAP7_75t_L g5974 ( 
.A1(n_5519),
.A2(n_3657),
.B(n_3546),
.Y(n_5974)
);

INVx3_ASAP7_75t_L g5975 ( 
.A(n_5542),
.Y(n_5975)
);

OAI21x1_ASAP7_75t_L g5976 ( 
.A1(n_5322),
.A2(n_3846),
.B(n_3827),
.Y(n_5976)
);

AOI221x1_ASAP7_75t_L g5977 ( 
.A1(n_5715),
.A2(n_1750),
.B1(n_1752),
.B2(n_1748),
.C(n_1745),
.Y(n_5977)
);

OAI21x1_ASAP7_75t_L g5978 ( 
.A1(n_5612),
.A2(n_3846),
.B(n_3827),
.Y(n_5978)
);

OAI21x1_ASAP7_75t_L g5979 ( 
.A1(n_5755),
.A2(n_3850),
.B(n_3827),
.Y(n_5979)
);

AOI21xp5_ASAP7_75t_L g5980 ( 
.A1(n_5544),
.A2(n_3657),
.B(n_3354),
.Y(n_5980)
);

INVx1_ASAP7_75t_SL g5981 ( 
.A(n_5726),
.Y(n_5981)
);

INVx2_ASAP7_75t_L g5982 ( 
.A(n_5525),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_5597),
.B(n_7),
.Y(n_5983)
);

NAND2xp5_ASAP7_75t_L g5984 ( 
.A(n_5628),
.B(n_8),
.Y(n_5984)
);

OAI21x1_ASAP7_75t_L g5985 ( 
.A1(n_5341),
.A2(n_5660),
.B(n_5734),
.Y(n_5985)
);

NAND2xp5_ASAP7_75t_L g5986 ( 
.A(n_5645),
.B(n_8),
.Y(n_5986)
);

NAND2xp5_ASAP7_75t_L g5987 ( 
.A(n_5674),
.B(n_9),
.Y(n_5987)
);

AOI22xp33_ASAP7_75t_L g5988 ( 
.A1(n_5527),
.A2(n_5342),
.B1(n_5501),
.B2(n_5561),
.Y(n_5988)
);

NOR2xp67_ASAP7_75t_L g5989 ( 
.A(n_5542),
.B(n_3851),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_5689),
.B(n_9),
.Y(n_5990)
);

OAI21x1_ASAP7_75t_L g5991 ( 
.A1(n_5736),
.A2(n_3860),
.B(n_3851),
.Y(n_5991)
);

AOI21xp5_ASAP7_75t_L g5992 ( 
.A1(n_5348),
.A2(n_5456),
.B(n_5563),
.Y(n_5992)
);

O2A1O1Ixp5_ASAP7_75t_L g5993 ( 
.A1(n_5447),
.A2(n_1755),
.B(n_1756),
.C(n_1753),
.Y(n_5993)
);

INVx1_ASAP7_75t_L g5994 ( 
.A(n_5737),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5748),
.Y(n_5995)
);

INVx2_ASAP7_75t_SL g5996 ( 
.A(n_5627),
.Y(n_5996)
);

INVx5_ASAP7_75t_L g5997 ( 
.A(n_5506),
.Y(n_5997)
);

OAI22x1_ASAP7_75t_L g5998 ( 
.A1(n_5360),
.A2(n_1395),
.B1(n_1396),
.B2(n_1394),
.Y(n_5998)
);

NAND2xp5_ASAP7_75t_L g5999 ( 
.A(n_5444),
.B(n_10),
.Y(n_5999)
);

OAI21x1_ASAP7_75t_L g6000 ( 
.A1(n_5669),
.A2(n_3860),
.B(n_3364),
.Y(n_6000)
);

OAI21x1_ASAP7_75t_L g6001 ( 
.A1(n_5323),
.A2(n_3860),
.B(n_3364),
.Y(n_6001)
);

CKINVDCx5p33_ASAP7_75t_R g6002 ( 
.A(n_5420),
.Y(n_6002)
);

OAI21xp5_ASAP7_75t_L g6003 ( 
.A1(n_5687),
.A2(n_3354),
.B(n_3333),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_SL g6004 ( 
.A(n_5429),
.B(n_2914),
.Y(n_6004)
);

BUFx2_ASAP7_75t_L g6005 ( 
.A(n_5549),
.Y(n_6005)
);

NAND2xp5_ASAP7_75t_L g6006 ( 
.A(n_5449),
.B(n_10),
.Y(n_6006)
);

NAND2xp5_ASAP7_75t_L g6007 ( 
.A(n_5451),
.B(n_10),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5756),
.Y(n_6008)
);

OAI21xp5_ASAP7_75t_L g6009 ( 
.A1(n_5735),
.A2(n_3333),
.B(n_3317),
.Y(n_6009)
);

AOI21x1_ASAP7_75t_L g6010 ( 
.A1(n_5662),
.A2(n_5665),
.B(n_5664),
.Y(n_6010)
);

AOI21x1_ASAP7_75t_L g6011 ( 
.A1(n_5671),
.A2(n_1640),
.B(n_1638),
.Y(n_6011)
);

NOR2xp33_ASAP7_75t_L g6012 ( 
.A(n_5353),
.B(n_342),
.Y(n_6012)
);

NAND2xp33_ASAP7_75t_L g6013 ( 
.A(n_5427),
.B(n_1400),
.Y(n_6013)
);

NAND2xp5_ASAP7_75t_L g6014 ( 
.A(n_5455),
.B(n_11),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5593),
.Y(n_6015)
);

AND2x2_ASAP7_75t_L g6016 ( 
.A(n_5367),
.B(n_11),
.Y(n_6016)
);

OAI21x1_ASAP7_75t_L g6017 ( 
.A1(n_5323),
.A2(n_5335),
.B(n_5661),
.Y(n_6017)
);

OAI21x1_ASAP7_75t_L g6018 ( 
.A1(n_5335),
.A2(n_2948),
.B(n_2902),
.Y(n_6018)
);

NAND2xp5_ASAP7_75t_SL g6019 ( 
.A(n_5459),
.B(n_2914),
.Y(n_6019)
);

AOI21xp5_ASAP7_75t_L g6020 ( 
.A1(n_5456),
.A2(n_5566),
.B(n_5378),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5440),
.Y(n_6021)
);

AOI21xp5_ASAP7_75t_L g6022 ( 
.A1(n_5668),
.A2(n_3657),
.B(n_3101),
.Y(n_6022)
);

INVx2_ASAP7_75t_L g6023 ( 
.A(n_5540),
.Y(n_6023)
);

NAND3xp33_ASAP7_75t_L g6024 ( 
.A(n_5482),
.B(n_1405),
.C(n_1402),
.Y(n_6024)
);

OR2x2_ASAP7_75t_L g6025 ( 
.A(n_5374),
.B(n_1645),
.Y(n_6025)
);

NAND2xp5_ASAP7_75t_L g6026 ( 
.A(n_5466),
.B(n_5370),
.Y(n_6026)
);

AOI21xp33_ASAP7_75t_L g6027 ( 
.A1(n_5705),
.A2(n_3384),
.B(n_3379),
.Y(n_6027)
);

OAI21xp5_ASAP7_75t_L g6028 ( 
.A1(n_5568),
.A2(n_3317),
.B(n_3314),
.Y(n_6028)
);

OAI21x1_ASAP7_75t_SL g6029 ( 
.A1(n_5469),
.A2(n_3908),
.B(n_3892),
.Y(n_6029)
);

AOI21x1_ASAP7_75t_L g6030 ( 
.A1(n_5677),
.A2(n_1682),
.B(n_1645),
.Y(n_6030)
);

OAI21xp5_ASAP7_75t_L g6031 ( 
.A1(n_5568),
.A2(n_3323),
.B(n_3314),
.Y(n_6031)
);

CKINVDCx5p33_ASAP7_75t_R g6032 ( 
.A(n_5633),
.Y(n_6032)
);

OAI22xp5_ASAP7_75t_L g6033 ( 
.A1(n_5551),
.A2(n_1425),
.B1(n_1432),
.B2(n_1409),
.Y(n_6033)
);

INVx1_ASAP7_75t_L g6034 ( 
.A(n_5373),
.Y(n_6034)
);

AO21x1_ASAP7_75t_L g6035 ( 
.A1(n_5523),
.A2(n_5620),
.B(n_5531),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5411),
.Y(n_6036)
);

OAI21xp5_ASAP7_75t_L g6037 ( 
.A1(n_5706),
.A2(n_3336),
.B(n_3323),
.Y(n_6037)
);

AOI21xp5_ASAP7_75t_L g6038 ( 
.A1(n_5582),
.A2(n_3101),
.B(n_3072),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5368),
.B(n_11),
.Y(n_6039)
);

AO31x2_ASAP7_75t_L g6040 ( 
.A1(n_5654),
.A2(n_3379),
.A3(n_3386),
.B(n_3384),
.Y(n_6040)
);

OAI21xp33_ASAP7_75t_L g6041 ( 
.A1(n_5482),
.A2(n_1434),
.B(n_1433),
.Y(n_6041)
);

NAND2xp5_ASAP7_75t_SL g6042 ( 
.A(n_5459),
.B(n_2914),
.Y(n_6042)
);

AOI21xp5_ASAP7_75t_L g6043 ( 
.A1(n_5679),
.A2(n_3101),
.B(n_3072),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5415),
.Y(n_6044)
);

OAI21x1_ASAP7_75t_L g6045 ( 
.A1(n_5573),
.A2(n_2948),
.B(n_2902),
.Y(n_6045)
);

NAND2xp5_ASAP7_75t_L g6046 ( 
.A(n_5707),
.B(n_12),
.Y(n_6046)
);

OAI21x1_ASAP7_75t_L g6047 ( 
.A1(n_5680),
.A2(n_3012),
.B(n_2902),
.Y(n_6047)
);

CKINVDCx6p67_ASAP7_75t_R g6048 ( 
.A(n_5454),
.Y(n_6048)
);

AND2x2_ASAP7_75t_L g6049 ( 
.A(n_5399),
.B(n_12),
.Y(n_6049)
);

OAI21xp5_ASAP7_75t_L g6050 ( 
.A1(n_5706),
.A2(n_3338),
.B(n_3336),
.Y(n_6050)
);

AOI21xp5_ASAP7_75t_L g6051 ( 
.A1(n_5692),
.A2(n_3113),
.B(n_3101),
.Y(n_6051)
);

AOI22xp5_ASAP7_75t_L g6052 ( 
.A1(n_5557),
.A2(n_1448),
.B1(n_1447),
.B2(n_2722),
.Y(n_6052)
);

AOI21xp5_ASAP7_75t_SL g6053 ( 
.A1(n_5430),
.A2(n_3557),
.B(n_3555),
.Y(n_6053)
);

AOI21xp5_ASAP7_75t_L g6054 ( 
.A1(n_5511),
.A2(n_3113),
.B(n_3101),
.Y(n_6054)
);

OAI21x1_ASAP7_75t_L g6055 ( 
.A1(n_5504),
.A2(n_3012),
.B(n_3386),
.Y(n_6055)
);

INVx3_ASAP7_75t_L g6056 ( 
.A(n_5731),
.Y(n_6056)
);

OAI21xp5_ASAP7_75t_L g6057 ( 
.A1(n_5676),
.A2(n_5402),
.B(n_5494),
.Y(n_6057)
);

AOI21x1_ASAP7_75t_L g6058 ( 
.A1(n_5577),
.A2(n_1683),
.B(n_1682),
.Y(n_6058)
);

AOI21xp5_ASAP7_75t_L g6059 ( 
.A1(n_5695),
.A2(n_3115),
.B(n_3113),
.Y(n_6059)
);

BUFx6f_ASAP7_75t_L g6060 ( 
.A(n_5427),
.Y(n_6060)
);

NAND2xp5_ASAP7_75t_L g6061 ( 
.A(n_5604),
.B(n_12),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_L g6062 ( 
.A(n_5653),
.B(n_13),
.Y(n_6062)
);

NAND2xp5_ASAP7_75t_L g6063 ( 
.A(n_5508),
.B(n_14),
.Y(n_6063)
);

INVx3_ASAP7_75t_L g6064 ( 
.A(n_5611),
.Y(n_6064)
);

OAI21x1_ASAP7_75t_L g6065 ( 
.A1(n_5502),
.A2(n_5424),
.B(n_5650),
.Y(n_6065)
);

AOI21xp5_ASAP7_75t_L g6066 ( 
.A1(n_5729),
.A2(n_3115),
.B(n_3113),
.Y(n_6066)
);

INVx2_ASAP7_75t_SL g6067 ( 
.A(n_5634),
.Y(n_6067)
);

OAI21x1_ASAP7_75t_L g6068 ( 
.A1(n_5502),
.A2(n_3012),
.B(n_3391),
.Y(n_6068)
);

INVxp67_ASAP7_75t_SL g6069 ( 
.A(n_5571),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_5547),
.Y(n_6070)
);

INVx3_ASAP7_75t_SL g6071 ( 
.A(n_5358),
.Y(n_6071)
);

AOI21xp5_ASAP7_75t_L g6072 ( 
.A1(n_5729),
.A2(n_3115),
.B(n_3113),
.Y(n_6072)
);

O2A1O1Ixp5_ASAP7_75t_L g6073 ( 
.A1(n_5732),
.A2(n_1764),
.B(n_1769),
.C(n_1762),
.Y(n_6073)
);

INVx1_ASAP7_75t_SL g6074 ( 
.A(n_5462),
.Y(n_6074)
);

AND2x6_ASAP7_75t_L g6075 ( 
.A(n_5610),
.B(n_3557),
.Y(n_6075)
);

OAI21x1_ASAP7_75t_L g6076 ( 
.A1(n_5651),
.A2(n_3407),
.B(n_3391),
.Y(n_6076)
);

AOI21xp5_ASAP7_75t_L g6077 ( 
.A1(n_5614),
.A2(n_3129),
.B(n_3115),
.Y(n_6077)
);

BUFx6f_ASAP7_75t_L g6078 ( 
.A(n_5590),
.Y(n_6078)
);

OAI21x1_ASAP7_75t_L g6079 ( 
.A1(n_5658),
.A2(n_5659),
.B(n_5630),
.Y(n_6079)
);

AOI21x1_ASAP7_75t_L g6080 ( 
.A1(n_5580),
.A2(n_1690),
.B(n_1683),
.Y(n_6080)
);

AOI21xp5_ASAP7_75t_L g6081 ( 
.A1(n_5364),
.A2(n_3129),
.B(n_3115),
.Y(n_6081)
);

INVx3_ASAP7_75t_L g6082 ( 
.A(n_5611),
.Y(n_6082)
);

AOI21xp5_ASAP7_75t_L g6083 ( 
.A1(n_5365),
.A2(n_3140),
.B(n_3129),
.Y(n_6083)
);

NAND2x1p5_ASAP7_75t_L g6084 ( 
.A(n_5610),
.B(n_3557),
.Y(n_6084)
);

BUFx2_ASAP7_75t_R g6085 ( 
.A(n_5605),
.Y(n_6085)
);

OAI21x1_ASAP7_75t_L g6086 ( 
.A1(n_5637),
.A2(n_3408),
.B(n_3407),
.Y(n_6086)
);

OAI21x1_ASAP7_75t_L g6087 ( 
.A1(n_5643),
.A2(n_3414),
.B(n_3408),
.Y(n_6087)
);

INVx2_ASAP7_75t_SL g6088 ( 
.A(n_5590),
.Y(n_6088)
);

OAI21x1_ASAP7_75t_SL g6089 ( 
.A1(n_5480),
.A2(n_3913),
.B(n_3908),
.Y(n_6089)
);

AND2x2_ASAP7_75t_SL g6090 ( 
.A(n_5524),
.B(n_1690),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_5562),
.Y(n_6091)
);

OAI21x1_ASAP7_75t_L g6092 ( 
.A1(n_5643),
.A2(n_3418),
.B(n_3414),
.Y(n_6092)
);

NAND2xp5_ASAP7_75t_L g6093 ( 
.A(n_5548),
.B(n_15),
.Y(n_6093)
);

A2O1A1Ixp33_ASAP7_75t_L g6094 ( 
.A1(n_5405),
.A2(n_2560),
.B(n_2609),
.C(n_2551),
.Y(n_6094)
);

OAI21xp5_ASAP7_75t_L g6095 ( 
.A1(n_5676),
.A2(n_5494),
.B(n_5386),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_L g6096 ( 
.A(n_5564),
.B(n_15),
.Y(n_6096)
);

NOR2x1_ASAP7_75t_L g6097 ( 
.A(n_5584),
.B(n_5588),
.Y(n_6097)
);

AOI21xp33_ASAP7_75t_L g6098 ( 
.A1(n_5380),
.A2(n_3421),
.B(n_3418),
.Y(n_6098)
);

OAI21x1_ASAP7_75t_L g6099 ( 
.A1(n_5514),
.A2(n_3428),
.B(n_3421),
.Y(n_6099)
);

AOI21xp5_ASAP7_75t_L g6100 ( 
.A1(n_5487),
.A2(n_3140),
.B(n_3129),
.Y(n_6100)
);

NOR2xp67_ASAP7_75t_L g6101 ( 
.A(n_5709),
.B(n_343),
.Y(n_6101)
);

AO31x2_ASAP7_75t_L g6102 ( 
.A1(n_5581),
.A2(n_3428),
.A3(n_3434),
.B(n_3431),
.Y(n_6102)
);

CKINVDCx20_ASAP7_75t_R g6103 ( 
.A(n_5723),
.Y(n_6103)
);

NAND2xp5_ASAP7_75t_L g6104 ( 
.A(n_5567),
.B(n_5484),
.Y(n_6104)
);

OAI21xp33_ASAP7_75t_L g6105 ( 
.A1(n_5404),
.A2(n_15),
.B(n_16),
.Y(n_6105)
);

NOR2xp33_ASAP7_75t_L g6106 ( 
.A(n_5388),
.B(n_5745),
.Y(n_6106)
);

BUFx8_ASAP7_75t_L g6107 ( 
.A(n_5590),
.Y(n_6107)
);

INVx2_ASAP7_75t_L g6108 ( 
.A(n_5609),
.Y(n_6108)
);

INVx3_ASAP7_75t_L g6109 ( 
.A(n_5611),
.Y(n_6109)
);

OR2x2_ASAP7_75t_L g6110 ( 
.A(n_5520),
.B(n_1701),
.Y(n_6110)
);

NAND2xp5_ASAP7_75t_L g6111 ( 
.A(n_5490),
.B(n_17),
.Y(n_6111)
);

AOI21xp5_ASAP7_75t_L g6112 ( 
.A1(n_5467),
.A2(n_3140),
.B(n_3129),
.Y(n_6112)
);

AND2x2_ASAP7_75t_L g6113 ( 
.A(n_5586),
.B(n_17),
.Y(n_6113)
);

AOI21xp5_ASAP7_75t_L g6114 ( 
.A1(n_5684),
.A2(n_3144),
.B(n_3140),
.Y(n_6114)
);

OAI21x1_ASAP7_75t_L g6115 ( 
.A1(n_5717),
.A2(n_3434),
.B(n_3431),
.Y(n_6115)
);

AOI21x1_ASAP7_75t_SL g6116 ( 
.A1(n_5720),
.A2(n_18),
.B(n_19),
.Y(n_6116)
);

BUFx8_ASAP7_75t_L g6117 ( 
.A(n_5758),
.Y(n_6117)
);

AO221x1_ASAP7_75t_L g6118 ( 
.A1(n_5622),
.A2(n_1572),
.B1(n_1582),
.B2(n_1481),
.C(n_1477),
.Y(n_6118)
);

AOI21x1_ASAP7_75t_L g6119 ( 
.A1(n_5596),
.A2(n_1717),
.B(n_1701),
.Y(n_6119)
);

OAI21x1_ASAP7_75t_L g6120 ( 
.A1(n_5710),
.A2(n_3443),
.B(n_3435),
.Y(n_6120)
);

A2O1A1Ixp33_ASAP7_75t_L g6121 ( 
.A1(n_5603),
.A2(n_2560),
.B(n_2609),
.C(n_2551),
.Y(n_6121)
);

AOI21xp5_ASAP7_75t_L g6122 ( 
.A1(n_5684),
.A2(n_3144),
.B(n_3140),
.Y(n_6122)
);

NAND2xp5_ASAP7_75t_L g6123 ( 
.A(n_5491),
.B(n_18),
.Y(n_6123)
);

NAND2x1p5_ASAP7_75t_L g6124 ( 
.A(n_5632),
.B(n_2924),
.Y(n_6124)
);

NAND2x1p5_ASAP7_75t_L g6125 ( 
.A(n_5632),
.B(n_2924),
.Y(n_6125)
);

AOI21x1_ASAP7_75t_L g6126 ( 
.A1(n_5545),
.A2(n_1727),
.B(n_1717),
.Y(n_6126)
);

NAND2x1_ASAP7_75t_L g6127 ( 
.A(n_5418),
.B(n_3326),
.Y(n_6127)
);

NAND2xp5_ASAP7_75t_L g6128 ( 
.A(n_5574),
.B(n_19),
.Y(n_6128)
);

OAI21x1_ASAP7_75t_L g6129 ( 
.A1(n_5713),
.A2(n_3443),
.B(n_3435),
.Y(n_6129)
);

AOI21x1_ASAP7_75t_L g6130 ( 
.A1(n_5546),
.A2(n_1759),
.B(n_1727),
.Y(n_6130)
);

NAND2xp5_ASAP7_75t_SL g6131 ( 
.A(n_5622),
.B(n_2924),
.Y(n_6131)
);

OAI21x1_ASAP7_75t_L g6132 ( 
.A1(n_5688),
.A2(n_3451),
.B(n_3446),
.Y(n_6132)
);

A2O1A1Ixp33_ASAP7_75t_L g6133 ( 
.A1(n_5350),
.A2(n_2684),
.B(n_2773),
.C(n_2722),
.Y(n_6133)
);

NAND2xp5_ASAP7_75t_L g6134 ( 
.A(n_5681),
.B(n_19),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_5693),
.B(n_20),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_5696),
.B(n_20),
.Y(n_6136)
);

AO31x2_ASAP7_75t_L g6137 ( 
.A1(n_5613),
.A2(n_3446),
.A3(n_3459),
.B(n_3451),
.Y(n_6137)
);

AOI21xp5_ASAP7_75t_L g6138 ( 
.A1(n_5684),
.A2(n_5333),
.B(n_5714),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_L g6139 ( 
.A(n_5500),
.B(n_20),
.Y(n_6139)
);

AND2x2_ASAP7_75t_L g6140 ( 
.A(n_5357),
.B(n_5622),
.Y(n_6140)
);

OAI21xp5_ASAP7_75t_L g6141 ( 
.A1(n_5432),
.A2(n_3340),
.B(n_3338),
.Y(n_6141)
);

OAI21x1_ASAP7_75t_L g6142 ( 
.A1(n_5377),
.A2(n_3464),
.B(n_3459),
.Y(n_6142)
);

OAI21xp5_ASAP7_75t_L g6143 ( 
.A1(n_5722),
.A2(n_3341),
.B(n_3340),
.Y(n_6143)
);

OAI21x1_ASAP7_75t_L g6144 ( 
.A1(n_5363),
.A2(n_3464),
.B(n_3377),
.Y(n_6144)
);

AO31x2_ASAP7_75t_L g6145 ( 
.A1(n_5636),
.A2(n_3523),
.A3(n_3524),
.B(n_3377),
.Y(n_6145)
);

OAI21x1_ASAP7_75t_L g6146 ( 
.A1(n_5629),
.A2(n_3523),
.B(n_3377),
.Y(n_6146)
);

OAI21x1_ASAP7_75t_L g6147 ( 
.A1(n_5744),
.A2(n_3524),
.B(n_3523),
.Y(n_6147)
);

AOI21xp5_ASAP7_75t_L g6148 ( 
.A1(n_5719),
.A2(n_3156),
.B(n_3144),
.Y(n_6148)
);

AOI21x1_ASAP7_75t_L g6149 ( 
.A1(n_5507),
.A2(n_1773),
.B(n_1759),
.Y(n_6149)
);

INVx5_ASAP7_75t_SL g6150 ( 
.A(n_5666),
.Y(n_6150)
);

NAND2xp5_ASAP7_75t_L g6151 ( 
.A(n_5515),
.B(n_21),
.Y(n_6151)
);

OAI21x1_ASAP7_75t_L g6152 ( 
.A1(n_5733),
.A2(n_3528),
.B(n_3524),
.Y(n_6152)
);

OAI21x1_ASAP7_75t_L g6153 ( 
.A1(n_5733),
.A2(n_3532),
.B(n_3528),
.Y(n_6153)
);

OAI21xp33_ASAP7_75t_L g6154 ( 
.A1(n_5754),
.A2(n_21),
.B(n_22),
.Y(n_6154)
);

OAI21xp5_ASAP7_75t_L g6155 ( 
.A1(n_5551),
.A2(n_3344),
.B(n_3341),
.Y(n_6155)
);

OAI21x1_ASAP7_75t_L g6156 ( 
.A1(n_5750),
.A2(n_3532),
.B(n_3528),
.Y(n_6156)
);

AOI21x1_ASAP7_75t_L g6157 ( 
.A1(n_5516),
.A2(n_5522),
.B(n_5518),
.Y(n_6157)
);

OAI21x1_ASAP7_75t_SL g6158 ( 
.A1(n_5498),
.A2(n_3919),
.B(n_3913),
.Y(n_6158)
);

OAI21x1_ASAP7_75t_L g6159 ( 
.A1(n_5753),
.A2(n_3535),
.B(n_3532),
.Y(n_6159)
);

AOI21xp5_ASAP7_75t_L g6160 ( 
.A1(n_5725),
.A2(n_3156),
.B(n_3144),
.Y(n_6160)
);

OAI21x1_ASAP7_75t_SL g6161 ( 
.A1(n_5652),
.A2(n_5728),
.B(n_5727),
.Y(n_6161)
);

INVx4_ASAP7_75t_L g6162 ( 
.A(n_5666),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_L g6163 ( 
.A(n_5443),
.B(n_23),
.Y(n_6163)
);

AO31x2_ASAP7_75t_L g6164 ( 
.A1(n_5663),
.A2(n_3539),
.A3(n_3540),
.B(n_3535),
.Y(n_6164)
);

INVxp67_ASAP7_75t_SL g6165 ( 
.A(n_5571),
.Y(n_6165)
);

NAND2xp5_ASAP7_75t_L g6166 ( 
.A(n_5700),
.B(n_24),
.Y(n_6166)
);

AND2x2_ASAP7_75t_L g6167 ( 
.A(n_5666),
.B(n_24),
.Y(n_6167)
);

OAI21x1_ASAP7_75t_L g6168 ( 
.A1(n_5452),
.A2(n_3539),
.B(n_3535),
.Y(n_6168)
);

NOR2xp33_ASAP7_75t_L g6169 ( 
.A(n_5439),
.B(n_5559),
.Y(n_6169)
);

AND2x6_ASAP7_75t_L g6170 ( 
.A(n_5600),
.B(n_5602),
.Y(n_6170)
);

OAI21xp33_ASAP7_75t_L g6171 ( 
.A1(n_5555),
.A2(n_24),
.B(n_25),
.Y(n_6171)
);

OAI21xp5_ASAP7_75t_L g6172 ( 
.A1(n_5395),
.A2(n_3348),
.B(n_3344),
.Y(n_6172)
);

OAI21x1_ASAP7_75t_L g6173 ( 
.A1(n_5675),
.A2(n_3540),
.B(n_3539),
.Y(n_6173)
);

OA21x2_ASAP7_75t_L g6174 ( 
.A1(n_5556),
.A2(n_1776),
.B(n_1773),
.Y(n_6174)
);

AOI21x1_ASAP7_75t_L g6175 ( 
.A1(n_5738),
.A2(n_1776),
.B(n_1772),
.Y(n_6175)
);

OAI21xp5_ASAP7_75t_L g6176 ( 
.A1(n_5465),
.A2(n_3352),
.B(n_3348),
.Y(n_6176)
);

NAND2xp5_ASAP7_75t_L g6177 ( 
.A(n_5570),
.B(n_25),
.Y(n_6177)
);

OAI21x1_ASAP7_75t_L g6178 ( 
.A1(n_5739),
.A2(n_3548),
.B(n_3540),
.Y(n_6178)
);

AND2x2_ASAP7_75t_L g6179 ( 
.A(n_5716),
.B(n_25),
.Y(n_6179)
);

BUFx12f_ASAP7_75t_L g6180 ( 
.A(n_5716),
.Y(n_6180)
);

INVx5_ASAP7_75t_L g6181 ( 
.A(n_5539),
.Y(n_6181)
);

OAI21xp5_ASAP7_75t_L g6182 ( 
.A1(n_5752),
.A2(n_3359),
.B(n_3352),
.Y(n_6182)
);

AND2x2_ASAP7_75t_L g6183 ( 
.A(n_5716),
.B(n_26),
.Y(n_6183)
);

OAI21x1_ASAP7_75t_L g6184 ( 
.A1(n_5740),
.A2(n_3559),
.B(n_3548),
.Y(n_6184)
);

INVx1_ASAP7_75t_SL g6185 ( 
.A(n_5757),
.Y(n_6185)
);

NAND2xp5_ASAP7_75t_L g6186 ( 
.A(n_5570),
.B(n_26),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_5741),
.B(n_5757),
.Y(n_6187)
);

AO21x1_ASAP7_75t_L g6188 ( 
.A1(n_5635),
.A2(n_5646),
.B(n_5640),
.Y(n_6188)
);

NAND2x1p5_ASAP7_75t_L g6189 ( 
.A(n_5757),
.B(n_5600),
.Y(n_6189)
);

INVx1_ASAP7_75t_L g6190 ( 
.A(n_5667),
.Y(n_6190)
);

OAI21xp5_ASAP7_75t_L g6191 ( 
.A1(n_5626),
.A2(n_3359),
.B(n_3919),
.Y(n_6191)
);

OR2x2_ASAP7_75t_L g6192 ( 
.A(n_5703),
.B(n_1770),
.Y(n_6192)
);

AND3x2_ASAP7_75t_L g6193 ( 
.A(n_5685),
.B(n_1775),
.C(n_1774),
.Y(n_6193)
);

OAI21x1_ASAP7_75t_L g6194 ( 
.A1(n_5742),
.A2(n_3559),
.B(n_3548),
.Y(n_6194)
);

OAI21x1_ASAP7_75t_SL g6195 ( 
.A1(n_5317),
.A2(n_3933),
.B(n_3932),
.Y(n_6195)
);

AND2x2_ASAP7_75t_L g6196 ( 
.A(n_5768),
.B(n_5524),
.Y(n_6196)
);

AOI221x1_ASAP7_75t_L g6197 ( 
.A1(n_6105),
.A2(n_5505),
.B1(n_5460),
.B2(n_5711),
.C(n_5690),
.Y(n_6197)
);

OAI21x1_ASAP7_75t_L g6198 ( 
.A1(n_5985),
.A2(n_5749),
.B(n_5616),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_5965),
.Y(n_6199)
);

NAND3x1_ASAP7_75t_L g6200 ( 
.A(n_5789),
.B(n_5655),
.C(n_5712),
.Y(n_6200)
);

OAI21x1_ASAP7_75t_L g6201 ( 
.A1(n_6079),
.A2(n_5585),
.B(n_5334),
.Y(n_6201)
);

NAND2x1p5_ASAP7_75t_L g6202 ( 
.A(n_5971),
.B(n_5602),
.Y(n_6202)
);

AOI22xp33_ASAP7_75t_L g6203 ( 
.A1(n_5801),
.A2(n_5539),
.B1(n_5418),
.B2(n_3477),
.Y(n_6203)
);

AO22x2_ASAP7_75t_L g6204 ( 
.A1(n_5910),
.A2(n_5423),
.B1(n_5672),
.B2(n_5539),
.Y(n_6204)
);

OR2x6_ASAP7_75t_L g6205 ( 
.A(n_5799),
.B(n_5418),
.Y(n_6205)
);

AOI221x1_ASAP7_75t_L g6206 ( 
.A1(n_6105),
.A2(n_5595),
.B1(n_5747),
.B2(n_1572),
.C(n_1582),
.Y(n_6206)
);

INVxp67_ASAP7_75t_SL g6207 ( 
.A(n_5821),
.Y(n_6207)
);

INVxp67_ASAP7_75t_SL g6208 ( 
.A(n_5885),
.Y(n_6208)
);

OAI21x1_ASAP7_75t_L g6209 ( 
.A1(n_5790),
.A2(n_5423),
.B(n_5672),
.Y(n_6209)
);

AOI21xp5_ASAP7_75t_L g6210 ( 
.A1(n_5992),
.A2(n_5499),
.B(n_5485),
.Y(n_6210)
);

INVx4_ASAP7_75t_L g6211 ( 
.A(n_6180),
.Y(n_6211)
);

NAND2xp5_ASAP7_75t_L g6212 ( 
.A(n_5929),
.B(n_344),
.Y(n_6212)
);

INVx5_ASAP7_75t_L g6213 ( 
.A(n_6075),
.Y(n_6213)
);

NAND2x1p5_ASAP7_75t_L g6214 ( 
.A(n_6127),
.B(n_2924),
.Y(n_6214)
);

A2O1A1Ixp33_ASAP7_75t_L g6215 ( 
.A1(n_6171),
.A2(n_5423),
.B(n_2684),
.C(n_28),
.Y(n_6215)
);

NOR2x1_ASAP7_75t_R g6216 ( 
.A(n_5871),
.B(n_2433),
.Y(n_6216)
);

OAI21x1_ASAP7_75t_L g6217 ( 
.A1(n_5767),
.A2(n_5672),
.B(n_3575),
.Y(n_6217)
);

OAI22x1_ASAP7_75t_L g6218 ( 
.A1(n_5820),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_6218)
);

OAI21xp5_ASAP7_75t_L g6219 ( 
.A1(n_5893),
.A2(n_3326),
.B(n_3932),
.Y(n_6219)
);

OA21x2_ASAP7_75t_L g6220 ( 
.A1(n_6138),
.A2(n_3575),
.B(n_3559),
.Y(n_6220)
);

CKINVDCx16_ASAP7_75t_R g6221 ( 
.A(n_6103),
.Y(n_6221)
);

OAI21x1_ASAP7_75t_L g6222 ( 
.A1(n_6017),
.A2(n_3589),
.B(n_3575),
.Y(n_6222)
);

AOI21x1_ASAP7_75t_L g6223 ( 
.A1(n_5865),
.A2(n_6010),
.B(n_5854),
.Y(n_6223)
);

AND2x4_ASAP7_75t_L g6224 ( 
.A(n_5855),
.B(n_27),
.Y(n_6224)
);

AO31x2_ASAP7_75t_L g6225 ( 
.A1(n_6008),
.A2(n_5805),
.A3(n_6035),
.B(n_5835),
.Y(n_6225)
);

OAI21xp5_ASAP7_75t_L g6226 ( 
.A1(n_5903),
.A2(n_3326),
.B(n_3933),
.Y(n_6226)
);

OR2x6_ASAP7_75t_L g6227 ( 
.A(n_5799),
.B(n_3441),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_6026),
.B(n_346),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_5934),
.Y(n_6229)
);

AOI21x1_ASAP7_75t_L g6230 ( 
.A1(n_5878),
.A2(n_3590),
.B(n_3589),
.Y(n_6230)
);

O2A1O1Ixp5_ASAP7_75t_L g6231 ( 
.A1(n_5933),
.A2(n_3940),
.B(n_3941),
.C(n_3938),
.Y(n_6231)
);

AOI22x1_ASAP7_75t_SL g6232 ( 
.A1(n_6032),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_6232)
);

AOI21xp5_ASAP7_75t_L g6233 ( 
.A1(n_5803),
.A2(n_5842),
.B(n_6066),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_5760),
.Y(n_6234)
);

OAI21x1_ASAP7_75t_L g6235 ( 
.A1(n_6065),
.A2(n_3590),
.B(n_3589),
.Y(n_6235)
);

INVx1_ASAP7_75t_L g6236 ( 
.A(n_5775),
.Y(n_6236)
);

A2O1A1Ixp33_ASAP7_75t_L g6237 ( 
.A1(n_6171),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_6237)
);

NAND2xp5_ASAP7_75t_L g6238 ( 
.A(n_5886),
.B(n_346),
.Y(n_6238)
);

INVx5_ASAP7_75t_L g6239 ( 
.A(n_6075),
.Y(n_6239)
);

CKINVDCx20_ASAP7_75t_R g6240 ( 
.A(n_5815),
.Y(n_6240)
);

INVx1_ASAP7_75t_L g6241 ( 
.A(n_5791),
.Y(n_6241)
);

AO31x2_ASAP7_75t_L g6242 ( 
.A1(n_5835),
.A2(n_3600),
.A3(n_3605),
.B(n_3590),
.Y(n_6242)
);

AOI21xp5_ASAP7_75t_L g6243 ( 
.A1(n_5803),
.A2(n_6072),
.B(n_6020),
.Y(n_6243)
);

OAI21xp5_ASAP7_75t_L g6244 ( 
.A1(n_5903),
.A2(n_3940),
.B(n_3938),
.Y(n_6244)
);

AOI21x1_ASAP7_75t_L g6245 ( 
.A1(n_6157),
.A2(n_3605),
.B(n_3600),
.Y(n_6245)
);

AO21x1_ASAP7_75t_L g6246 ( 
.A1(n_5933),
.A2(n_30),
.B(n_32),
.Y(n_6246)
);

NOR2xp33_ASAP7_75t_L g6247 ( 
.A(n_6071),
.B(n_347),
.Y(n_6247)
);

INVx3_ASAP7_75t_L g6248 ( 
.A(n_5855),
.Y(n_6248)
);

AO32x2_ASAP7_75t_L g6249 ( 
.A1(n_6067),
.A2(n_3534),
.A3(n_3527),
.B1(n_3448),
.B2(n_34),
.Y(n_6249)
);

INVxp67_ASAP7_75t_L g6250 ( 
.A(n_5884),
.Y(n_6250)
);

OAI21x1_ASAP7_75t_L g6251 ( 
.A1(n_5771),
.A2(n_3605),
.B(n_3600),
.Y(n_6251)
);

OAI21x1_ASAP7_75t_L g6252 ( 
.A1(n_5776),
.A2(n_3615),
.B(n_3607),
.Y(n_6252)
);

OAI21x1_ASAP7_75t_L g6253 ( 
.A1(n_5779),
.A2(n_3615),
.B(n_3607),
.Y(n_6253)
);

NAND2xp5_ASAP7_75t_L g6254 ( 
.A(n_5868),
.B(n_347),
.Y(n_6254)
);

INVx2_ASAP7_75t_SL g6255 ( 
.A(n_5823),
.Y(n_6255)
);

O2A1O1Ixp5_ASAP7_75t_L g6256 ( 
.A1(n_5947),
.A2(n_3943),
.B(n_3941),
.C(n_35),
.Y(n_6256)
);

NAND2xp5_ASAP7_75t_L g6257 ( 
.A(n_5761),
.B(n_348),
.Y(n_6257)
);

AOI211x1_ASAP7_75t_L g6258 ( 
.A1(n_6188),
.A2(n_36),
.B(n_32),
.C(n_33),
.Y(n_6258)
);

NAND2xp5_ASAP7_75t_L g6259 ( 
.A(n_6034),
.B(n_6036),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_6044),
.B(n_348),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_5795),
.B(n_349),
.Y(n_6261)
);

AND2x2_ASAP7_75t_L g6262 ( 
.A(n_5866),
.B(n_36),
.Y(n_6262)
);

OAI21xp5_ASAP7_75t_L g6263 ( 
.A1(n_5947),
.A2(n_3943),
.B(n_3527),
.Y(n_6263)
);

AOI21xp5_ASAP7_75t_SL g6264 ( 
.A1(n_6101),
.A2(n_2943),
.B(n_2924),
.Y(n_6264)
);

AND2x4_ASAP7_75t_L g6265 ( 
.A(n_5889),
.B(n_37),
.Y(n_6265)
);

INVx1_ASAP7_75t_L g6266 ( 
.A(n_5826),
.Y(n_6266)
);

BUFx12f_ASAP7_75t_L g6267 ( 
.A(n_5770),
.Y(n_6267)
);

AOI211x1_ASAP7_75t_L g6268 ( 
.A1(n_5777),
.A2(n_40),
.B(n_37),
.C(n_38),
.Y(n_6268)
);

NAND2xp5_ASAP7_75t_L g6269 ( 
.A(n_5845),
.B(n_351),
.Y(n_6269)
);

AO31x2_ASAP7_75t_L g6270 ( 
.A1(n_5817),
.A2(n_3615),
.A3(n_3616),
.B(n_3607),
.Y(n_6270)
);

HB1xp67_ASAP7_75t_L g6271 ( 
.A(n_5766),
.Y(n_6271)
);

NAND2xp5_ASAP7_75t_SL g6272 ( 
.A(n_5925),
.B(n_2943),
.Y(n_6272)
);

AOI21xp5_ASAP7_75t_L g6273 ( 
.A1(n_5950),
.A2(n_3534),
.B(n_3448),
.Y(n_6273)
);

OAI22xp5_ASAP7_75t_L g6274 ( 
.A1(n_5896),
.A2(n_2773),
.B1(n_2774),
.B2(n_2722),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5872),
.Y(n_6275)
);

CKINVDCx5p33_ASAP7_75t_R g6276 ( 
.A(n_6002),
.Y(n_6276)
);

AOI21xp5_ASAP7_75t_L g6277 ( 
.A1(n_5950),
.A2(n_2964),
.B(n_2943),
.Y(n_6277)
);

AOI21xp5_ASAP7_75t_L g6278 ( 
.A1(n_5858),
.A2(n_2964),
.B(n_2943),
.Y(n_6278)
);

OAI21x1_ASAP7_75t_L g6279 ( 
.A1(n_5806),
.A2(n_3622),
.B(n_3616),
.Y(n_6279)
);

OA21x2_ASAP7_75t_L g6280 ( 
.A1(n_5777),
.A2(n_3622),
.B(n_3616),
.Y(n_6280)
);

NAND2xp5_ASAP7_75t_L g6281 ( 
.A(n_5941),
.B(n_351),
.Y(n_6281)
);

AOI21xp5_ASAP7_75t_L g6282 ( 
.A1(n_5858),
.A2(n_2964),
.B(n_2943),
.Y(n_6282)
);

NOR2xp33_ASAP7_75t_L g6283 ( 
.A(n_6048),
.B(n_352),
.Y(n_6283)
);

OAI21xp5_ASAP7_75t_L g6284 ( 
.A1(n_5798),
.A2(n_3045),
.B(n_3037),
.Y(n_6284)
);

AOI221x1_ASAP7_75t_L g6285 ( 
.A1(n_5841),
.A2(n_1572),
.B1(n_1582),
.B2(n_1481),
.C(n_1477),
.Y(n_6285)
);

AOI221xp5_ASAP7_75t_SL g6286 ( 
.A1(n_5857),
.A2(n_41),
.B1(n_37),
.B2(n_40),
.C(n_42),
.Y(n_6286)
);

AO32x2_ASAP7_75t_L g6287 ( 
.A1(n_5850),
.A2(n_42),
.A3(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_6287)
);

NOR2xp33_ASAP7_75t_L g6288 ( 
.A(n_5762),
.B(n_353),
.Y(n_6288)
);

OAI21xp33_ASAP7_75t_L g6289 ( 
.A1(n_6177),
.A2(n_1481),
.B(n_1477),
.Y(n_6289)
);

AND2x4_ASAP7_75t_L g6290 ( 
.A(n_5889),
.B(n_43),
.Y(n_6290)
);

OAI21x1_ASAP7_75t_L g6291 ( 
.A1(n_6114),
.A2(n_3732),
.B(n_3622),
.Y(n_6291)
);

OAI21x1_ASAP7_75t_L g6292 ( 
.A1(n_6122),
.A2(n_3736),
.B(n_3732),
.Y(n_6292)
);

NAND2xp5_ASAP7_75t_L g6293 ( 
.A(n_6104),
.B(n_354),
.Y(n_6293)
);

A2O1A1Ixp33_ASAP7_75t_L g6294 ( 
.A1(n_6154),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_6294)
);

AOI21xp5_ASAP7_75t_L g6295 ( 
.A1(n_6095),
.A2(n_6112),
.B(n_6051),
.Y(n_6295)
);

NAND2xp5_ASAP7_75t_L g6296 ( 
.A(n_5916),
.B(n_354),
.Y(n_6296)
);

NAND2xp5_ASAP7_75t_L g6297 ( 
.A(n_5763),
.B(n_355),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_5887),
.B(n_5846),
.Y(n_6298)
);

NAND2xp5_ASAP7_75t_L g6299 ( 
.A(n_5968),
.B(n_357),
.Y(n_6299)
);

OAI21xp5_ASAP7_75t_L g6300 ( 
.A1(n_5914),
.A2(n_3052),
.B(n_3045),
.Y(n_6300)
);

NAND2xp5_ASAP7_75t_L g6301 ( 
.A(n_5968),
.B(n_358),
.Y(n_6301)
);

OAI21x1_ASAP7_75t_L g6302 ( 
.A1(n_6043),
.A2(n_3736),
.B(n_3732),
.Y(n_6302)
);

NAND2xp5_ASAP7_75t_L g6303 ( 
.A(n_5981),
.B(n_359),
.Y(n_6303)
);

AO21x2_ASAP7_75t_L g6304 ( 
.A1(n_5946),
.A2(n_3736),
.B(n_3679),
.Y(n_6304)
);

AO22x2_ASAP7_75t_L g6305 ( 
.A1(n_6021),
.A2(n_3477),
.B1(n_3478),
.B2(n_3473),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_5875),
.Y(n_6306)
);

INVxp67_ASAP7_75t_L g6307 ( 
.A(n_6005),
.Y(n_6307)
);

BUFx6f_ASAP7_75t_L g6308 ( 
.A(n_6078),
.Y(n_6308)
);

AND2x2_ASAP7_75t_L g6309 ( 
.A(n_5981),
.B(n_44),
.Y(n_6309)
);

AO32x2_ASAP7_75t_L g6310 ( 
.A1(n_6088),
.A2(n_47),
.A3(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_5781),
.Y(n_6311)
);

AOI211x1_ASAP7_75t_L g6312 ( 
.A1(n_6061),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_6312)
);

NAND2xp33_ASAP7_75t_R g6313 ( 
.A(n_5784),
.B(n_47),
.Y(n_6313)
);

AND2x2_ASAP7_75t_L g6314 ( 
.A(n_5902),
.B(n_49),
.Y(n_6314)
);

NAND2xp5_ASAP7_75t_L g6315 ( 
.A(n_6015),
.B(n_359),
.Y(n_6315)
);

OAI21xp5_ASAP7_75t_L g6316 ( 
.A1(n_6024),
.A2(n_3053),
.B(n_3052),
.Y(n_6316)
);

OAI21x1_ASAP7_75t_L g6317 ( 
.A1(n_5788),
.A2(n_3087),
.B(n_3084),
.Y(n_6317)
);

OR2x2_ASAP7_75t_L g6318 ( 
.A(n_5764),
.B(n_49),
.Y(n_6318)
);

OAI21x1_ASAP7_75t_L g6319 ( 
.A1(n_6059),
.A2(n_3094),
.B(n_3473),
.Y(n_6319)
);

NAND2xp5_ASAP7_75t_L g6320 ( 
.A(n_6074),
.B(n_360),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5888),
.Y(n_6321)
);

NAND2xp5_ASAP7_75t_L g6322 ( 
.A(n_6074),
.B(n_360),
.Y(n_6322)
);

INVx1_ASAP7_75t_SL g6323 ( 
.A(n_6085),
.Y(n_6323)
);

NOR2xp33_ASAP7_75t_L g6324 ( 
.A(n_6169),
.B(n_361),
.Y(n_6324)
);

NAND2xp5_ASAP7_75t_L g6325 ( 
.A(n_5780),
.B(n_361),
.Y(n_6325)
);

INVx2_ASAP7_75t_L g6326 ( 
.A(n_5816),
.Y(n_6326)
);

NAND2xp5_ASAP7_75t_L g6327 ( 
.A(n_5995),
.B(n_362),
.Y(n_6327)
);

OAI21x1_ASAP7_75t_L g6328 ( 
.A1(n_6100),
.A2(n_3094),
.B(n_3478),
.Y(n_6328)
);

OAI21x1_ASAP7_75t_L g6329 ( 
.A1(n_5962),
.A2(n_3483),
.B(n_3482),
.Y(n_6329)
);

AOI21xp5_ASAP7_75t_L g6330 ( 
.A1(n_6095),
.A2(n_2970),
.B(n_2964),
.Y(n_6330)
);

O2A1O1Ixp5_ASAP7_75t_SL g6331 ( 
.A1(n_5958),
.A2(n_2480),
.B(n_2467),
.C(n_3290),
.Y(n_6331)
);

NAND3xp33_ASAP7_75t_L g6332 ( 
.A(n_5773),
.B(n_1572),
.C(n_1481),
.Y(n_6332)
);

OAI22xp33_ASAP7_75t_L g6333 ( 
.A1(n_6057),
.A2(n_2773),
.B1(n_2774),
.B2(n_2722),
.Y(n_6333)
);

CKINVDCx20_ASAP7_75t_R g6334 ( 
.A(n_6117),
.Y(n_6334)
);

INVx3_ASAP7_75t_L g6335 ( 
.A(n_5902),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_5891),
.B(n_5900),
.Y(n_6336)
);

OAI22xp33_ASAP7_75t_L g6337 ( 
.A1(n_6057),
.A2(n_2773),
.B1(n_2774),
.B2(n_2722),
.Y(n_6337)
);

NAND3xp33_ASAP7_75t_L g6338 ( 
.A(n_5773),
.B(n_6006),
.C(n_5999),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_5935),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_5942),
.Y(n_6340)
);

OAI21x1_ASAP7_75t_L g6341 ( 
.A1(n_5802),
.A2(n_3483),
.B(n_3482),
.Y(n_6341)
);

INVx5_ASAP7_75t_L g6342 ( 
.A(n_6075),
.Y(n_6342)
);

AOI21xp5_ASAP7_75t_L g6343 ( 
.A1(n_5834),
.A2(n_2970),
.B(n_2964),
.Y(n_6343)
);

INVx2_ASAP7_75t_L g6344 ( 
.A(n_5818),
.Y(n_6344)
);

AOI21x1_ASAP7_75t_L g6345 ( 
.A1(n_5917),
.A2(n_5919),
.B(n_5861),
.Y(n_6345)
);

BUFx3_ASAP7_75t_L g6346 ( 
.A(n_5996),
.Y(n_6346)
);

OAI21x1_ASAP7_75t_L g6347 ( 
.A1(n_5836),
.A2(n_5869),
.B(n_5961),
.Y(n_6347)
);

OAI21xp33_ASAP7_75t_L g6348 ( 
.A1(n_6186),
.A2(n_1572),
.B(n_1481),
.Y(n_6348)
);

AOI221xp5_ASAP7_75t_SL g6349 ( 
.A1(n_6012),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.C(n_53),
.Y(n_6349)
);

A2O1A1Ixp33_ASAP7_75t_L g6350 ( 
.A1(n_6154),
.A2(n_6041),
.B(n_6024),
.C(n_6101),
.Y(n_6350)
);

AND2x2_ASAP7_75t_L g6351 ( 
.A(n_5975),
.B(n_51),
.Y(n_6351)
);

INVx4_ASAP7_75t_L g6352 ( 
.A(n_6078),
.Y(n_6352)
);

INVx5_ASAP7_75t_L g6353 ( 
.A(n_6075),
.Y(n_6353)
);

INVx1_ASAP7_75t_L g6354 ( 
.A(n_5994),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_5769),
.Y(n_6355)
);

OAI21x1_ASAP7_75t_L g6356 ( 
.A1(n_6011),
.A2(n_6030),
.B(n_5897),
.Y(n_6356)
);

OAI21x1_ASAP7_75t_L g6357 ( 
.A1(n_6058),
.A2(n_3491),
.B(n_3490),
.Y(n_6357)
);

NAND2xp33_ASAP7_75t_L g6358 ( 
.A(n_5925),
.B(n_2970),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_SL g6359 ( 
.A(n_5925),
.B(n_2970),
.Y(n_6359)
);

OAI21x1_ASAP7_75t_L g6360 ( 
.A1(n_6080),
.A2(n_3491),
.B(n_3490),
.Y(n_6360)
);

BUFx2_ASAP7_75t_R g6361 ( 
.A(n_6063),
.Y(n_6361)
);

AOI21xp5_ASAP7_75t_L g6362 ( 
.A1(n_5840),
.A2(n_2970),
.B(n_3117),
.Y(n_6362)
);

BUFx6f_ASAP7_75t_L g6363 ( 
.A(n_6078),
.Y(n_6363)
);

AOI21x1_ASAP7_75t_L g6364 ( 
.A1(n_5944),
.A2(n_3053),
.B(n_3496),
.Y(n_6364)
);

OAI21x1_ASAP7_75t_L g6365 ( 
.A1(n_6149),
.A2(n_3501),
.B(n_3496),
.Y(n_6365)
);

A2O1A1Ixp33_ASAP7_75t_L g6366 ( 
.A1(n_6041),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_6366)
);

OAI21x1_ASAP7_75t_L g6367 ( 
.A1(n_6126),
.A2(n_3505),
.B(n_3501),
.Y(n_6367)
);

AOI21xp5_ASAP7_75t_L g6368 ( 
.A1(n_5785),
.A2(n_3120),
.B(n_3117),
.Y(n_6368)
);

AOI21xp5_ASAP7_75t_L g6369 ( 
.A1(n_5827),
.A2(n_3121),
.B(n_3120),
.Y(n_6369)
);

NAND2xp5_ASAP7_75t_L g6370 ( 
.A(n_5862),
.B(n_363),
.Y(n_6370)
);

NOR3xp33_ASAP7_75t_SL g6371 ( 
.A(n_5931),
.B(n_52),
.C(n_53),
.Y(n_6371)
);

BUFx6f_ASAP7_75t_L g6372 ( 
.A(n_5796),
.Y(n_6372)
);

INVx2_ASAP7_75t_L g6373 ( 
.A(n_5819),
.Y(n_6373)
);

NAND2xp5_ASAP7_75t_L g6374 ( 
.A(n_5877),
.B(n_364),
.Y(n_6374)
);

OAI21x1_ASAP7_75t_L g6375 ( 
.A1(n_6130),
.A2(n_3508),
.B(n_3505),
.Y(n_6375)
);

OAI21x1_ASAP7_75t_L g6376 ( 
.A1(n_5830),
.A2(n_3513),
.B(n_3508),
.Y(n_6376)
);

NOR4xp25_ASAP7_75t_L g6377 ( 
.A(n_6007),
.B(n_56),
.C(n_54),
.D(n_55),
.Y(n_6377)
);

NAND2xp5_ASAP7_75t_L g6378 ( 
.A(n_6016),
.B(n_364),
.Y(n_6378)
);

INVx2_ASAP7_75t_L g6379 ( 
.A(n_5883),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_5898),
.Y(n_6380)
);

NAND3xp33_ASAP7_75t_L g6381 ( 
.A(n_6014),
.B(n_1636),
.C(n_1582),
.Y(n_6381)
);

AOI21xp5_ASAP7_75t_L g6382 ( 
.A1(n_5827),
.A2(n_5772),
.B(n_5980),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6070),
.Y(n_6383)
);

BUFx4_ASAP7_75t_SL g6384 ( 
.A(n_5799),
.Y(n_6384)
);

INVx3_ASAP7_75t_L g6385 ( 
.A(n_5975),
.Y(n_6385)
);

O2A1O1Ixp33_ASAP7_75t_SL g6386 ( 
.A1(n_5853),
.A2(n_57),
.B(n_54),
.C(n_55),
.Y(n_6386)
);

AOI21xp5_ASAP7_75t_L g6387 ( 
.A1(n_5772),
.A2(n_3122),
.B(n_3121),
.Y(n_6387)
);

AO31x2_ASAP7_75t_L g6388 ( 
.A1(n_6133),
.A2(n_5957),
.A3(n_6190),
.B(n_5895),
.Y(n_6388)
);

OAI21x1_ASAP7_75t_L g6389 ( 
.A1(n_6119),
.A2(n_5848),
.B(n_6184),
.Y(n_6389)
);

A2O1A1Ixp33_ASAP7_75t_L g6390 ( 
.A1(n_5960),
.A2(n_59),
.B(n_57),
.C(n_58),
.Y(n_6390)
);

AND2x2_ASAP7_75t_L g6391 ( 
.A(n_6140),
.B(n_58),
.Y(n_6391)
);

BUFx3_ASAP7_75t_L g6392 ( 
.A(n_6117),
.Y(n_6392)
);

AOI21xp5_ASAP7_75t_L g6393 ( 
.A1(n_5920),
.A2(n_3124),
.B(n_3122),
.Y(n_6393)
);

AND2x4_ASAP7_75t_L g6394 ( 
.A(n_5970),
.B(n_59),
.Y(n_6394)
);

AOI21xp5_ASAP7_75t_L g6395 ( 
.A1(n_5936),
.A2(n_3135),
.B(n_3124),
.Y(n_6395)
);

AO31x2_ASAP7_75t_L g6396 ( 
.A1(n_5909),
.A2(n_3516),
.A3(n_3563),
.B(n_3513),
.Y(n_6396)
);

NOR2xp67_ASAP7_75t_L g6397 ( 
.A(n_5970),
.B(n_59),
.Y(n_6397)
);

AND2x2_ASAP7_75t_L g6398 ( 
.A(n_5832),
.B(n_6056),
.Y(n_6398)
);

AO31x2_ASAP7_75t_L g6399 ( 
.A1(n_5918),
.A2(n_3563),
.A3(n_3571),
.B(n_3516),
.Y(n_6399)
);

OAI21x1_ASAP7_75t_L g6400 ( 
.A1(n_6178),
.A2(n_3573),
.B(n_3571),
.Y(n_6400)
);

AND2x2_ASAP7_75t_L g6401 ( 
.A(n_6056),
.B(n_60),
.Y(n_6401)
);

OAI21x1_ASAP7_75t_L g6402 ( 
.A1(n_5837),
.A2(n_3627),
.B(n_3573),
.Y(n_6402)
);

OAI21x1_ASAP7_75t_L g6403 ( 
.A1(n_5843),
.A2(n_3634),
.B(n_3627),
.Y(n_6403)
);

O2A1O1Ixp33_ASAP7_75t_L g6404 ( 
.A1(n_5828),
.A2(n_64),
.B(n_61),
.C(n_62),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_L g6405 ( 
.A(n_6097),
.B(n_365),
.Y(n_6405)
);

O2A1O1Ixp5_ASAP7_75t_SL g6406 ( 
.A1(n_5983),
.A2(n_2480),
.B(n_2467),
.C(n_3290),
.Y(n_6406)
);

AO31x2_ASAP7_75t_L g6407 ( 
.A1(n_5922),
.A2(n_3636),
.A3(n_3643),
.B(n_3634),
.Y(n_6407)
);

AOI21x1_ASAP7_75t_L g6408 ( 
.A1(n_5984),
.A2(n_5987),
.B(n_5986),
.Y(n_6408)
);

AOI21xp5_ASAP7_75t_L g6409 ( 
.A1(n_5851),
.A2(n_3150),
.B(n_3135),
.Y(n_6409)
);

INVx5_ASAP7_75t_L g6410 ( 
.A(n_5796),
.Y(n_6410)
);

OAI22x1_ASAP7_75t_L g6411 ( 
.A1(n_5970),
.A2(n_5997),
.B1(n_6039),
.B2(n_6106),
.Y(n_6411)
);

NAND2xp5_ASAP7_75t_L g6412 ( 
.A(n_5948),
.B(n_365),
.Y(n_6412)
);

OAI21x1_ASAP7_75t_L g6413 ( 
.A1(n_6175),
.A2(n_3643),
.B(n_3636),
.Y(n_6413)
);

NAND2xp5_ASAP7_75t_L g6414 ( 
.A(n_6111),
.B(n_366),
.Y(n_6414)
);

NOR2x1_ASAP7_75t_SL g6415 ( 
.A(n_5923),
.B(n_1582),
.Y(n_6415)
);

NAND2xp5_ASAP7_75t_L g6416 ( 
.A(n_6123),
.B(n_366),
.Y(n_6416)
);

AOI21xp5_ASAP7_75t_L g6417 ( 
.A1(n_5851),
.A2(n_3159),
.B(n_3150),
.Y(n_6417)
);

NAND2xp5_ASAP7_75t_L g6418 ( 
.A(n_6163),
.B(n_368),
.Y(n_6418)
);

NAND2xp5_ASAP7_75t_L g6419 ( 
.A(n_5838),
.B(n_369),
.Y(n_6419)
);

INVx4_ASAP7_75t_L g6420 ( 
.A(n_5796),
.Y(n_6420)
);

OA21x2_ASAP7_75t_L g6421 ( 
.A1(n_6069),
.A2(n_6165),
.B(n_5990),
.Y(n_6421)
);

AND2x2_ASAP7_75t_L g6422 ( 
.A(n_6185),
.B(n_61),
.Y(n_6422)
);

AND2x2_ASAP7_75t_L g6423 ( 
.A(n_6185),
.B(n_61),
.Y(n_6423)
);

NAND2xp5_ASAP7_75t_L g6424 ( 
.A(n_5915),
.B(n_371),
.Y(n_6424)
);

INVxp67_ASAP7_75t_SL g6425 ( 
.A(n_6025),
.Y(n_6425)
);

INVx2_ASAP7_75t_L g6426 ( 
.A(n_5951),
.Y(n_6426)
);

INVx1_ASAP7_75t_L g6427 ( 
.A(n_5956),
.Y(n_6427)
);

AO31x2_ASAP7_75t_L g6428 ( 
.A1(n_5959),
.A2(n_6023),
.A3(n_6091),
.B(n_5982),
.Y(n_6428)
);

INVx3_ASAP7_75t_L g6429 ( 
.A(n_6162),
.Y(n_6429)
);

CKINVDCx5p33_ASAP7_75t_R g6430 ( 
.A(n_6107),
.Y(n_6430)
);

O2A1O1Ixp5_ASAP7_75t_SL g6431 ( 
.A1(n_5860),
.A2(n_2480),
.B(n_3293),
.C(n_3290),
.Y(n_6431)
);

OAI21x1_ASAP7_75t_L g6432 ( 
.A1(n_5973),
.A2(n_5913),
.B(n_5812),
.Y(n_6432)
);

BUFx3_ASAP7_75t_L g6433 ( 
.A(n_6107),
.Y(n_6433)
);

BUFx12f_ASAP7_75t_L g6434 ( 
.A(n_6113),
.Y(n_6434)
);

A2O1A1Ixp33_ASAP7_75t_L g6435 ( 
.A1(n_5960),
.A2(n_65),
.B(n_62),
.C(n_64),
.Y(n_6435)
);

OAI21xp5_ASAP7_75t_L g6436 ( 
.A1(n_5782),
.A2(n_64),
.B(n_65),
.Y(n_6436)
);

OAI21xp5_ASAP7_75t_L g6437 ( 
.A1(n_5794),
.A2(n_66),
.B(n_67),
.Y(n_6437)
);

NAND2xp5_ASAP7_75t_L g6438 ( 
.A(n_6187),
.B(n_371),
.Y(n_6438)
);

OAI21xp5_ASAP7_75t_L g6439 ( 
.A1(n_5954),
.A2(n_66),
.B(n_67),
.Y(n_6439)
);

NAND2xp5_ASAP7_75t_SL g6440 ( 
.A(n_5925),
.B(n_5881),
.Y(n_6440)
);

AND2x2_ASAP7_75t_L g6441 ( 
.A(n_6049),
.B(n_66),
.Y(n_6441)
);

NAND2xp5_ASAP7_75t_L g6442 ( 
.A(n_6128),
.B(n_372),
.Y(n_6442)
);

AOI21xp5_ASAP7_75t_L g6443 ( 
.A1(n_5774),
.A2(n_3166),
.B(n_3159),
.Y(n_6443)
);

OAI21x1_ASAP7_75t_L g6444 ( 
.A1(n_5793),
.A2(n_3665),
.B(n_3659),
.Y(n_6444)
);

AO31x2_ASAP7_75t_L g6445 ( 
.A1(n_6108),
.A2(n_3665),
.A3(n_3666),
.B(n_3659),
.Y(n_6445)
);

NAND2xp5_ASAP7_75t_L g6446 ( 
.A(n_6139),
.B(n_373),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_5792),
.Y(n_6447)
);

AOI21x1_ASAP7_75t_L g6448 ( 
.A1(n_5899),
.A2(n_3677),
.B(n_3666),
.Y(n_6448)
);

INVxp67_ASAP7_75t_SL g6449 ( 
.A(n_5989),
.Y(n_6449)
);

O2A1O1Ixp33_ASAP7_75t_L g6450 ( 
.A1(n_5927),
.A2(n_5969),
.B(n_6033),
.C(n_6161),
.Y(n_6450)
);

NAND2xp5_ASAP7_75t_L g6451 ( 
.A(n_6151),
.B(n_374),
.Y(n_6451)
);

OAI21x1_ASAP7_75t_L g6452 ( 
.A1(n_5793),
.A2(n_3678),
.B(n_3677),
.Y(n_6452)
);

OAI22xp5_ASAP7_75t_L g6453 ( 
.A1(n_5988),
.A2(n_2774),
.B1(n_2773),
.B2(n_3293),
.Y(n_6453)
);

BUFx12f_ASAP7_75t_L g6454 ( 
.A(n_5881),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_5792),
.Y(n_6455)
);

NAND2xp5_ASAP7_75t_L g6456 ( 
.A(n_6134),
.B(n_374),
.Y(n_6456)
);

OAI22x1_ASAP7_75t_L g6457 ( 
.A1(n_5997),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_6457)
);

NAND2xp5_ASAP7_75t_L g6458 ( 
.A(n_6046),
.B(n_375),
.Y(n_6458)
);

OAI21x1_ASAP7_75t_L g6459 ( 
.A1(n_6054),
.A2(n_6089),
.B(n_6029),
.Y(n_6459)
);

NAND2xp5_ASAP7_75t_L g6460 ( 
.A(n_6166),
.B(n_375),
.Y(n_6460)
);

AOI21xp5_ASAP7_75t_L g6461 ( 
.A1(n_5800),
.A2(n_3167),
.B(n_3166),
.Y(n_6461)
);

INVx2_ASAP7_75t_L g6462 ( 
.A(n_5792),
.Y(n_6462)
);

INVx1_ASAP7_75t_L g6463 ( 
.A(n_6110),
.Y(n_6463)
);

A2O1A1Ixp33_ASAP7_75t_L g6464 ( 
.A1(n_5967),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_6192),
.Y(n_6465)
);

A2O1A1Ixp33_ASAP7_75t_L g6466 ( 
.A1(n_5967),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_6466)
);

AOI21xp5_ASAP7_75t_L g6467 ( 
.A1(n_5870),
.A2(n_3172),
.B(n_3167),
.Y(n_6467)
);

OAI22xp5_ASAP7_75t_L g6468 ( 
.A1(n_5833),
.A2(n_2774),
.B1(n_3302),
.B2(n_3293),
.Y(n_6468)
);

OAI21x1_ASAP7_75t_L g6469 ( 
.A1(n_5852),
.A2(n_3679),
.B(n_3678),
.Y(n_6469)
);

AND2x2_ASAP7_75t_L g6470 ( 
.A(n_6162),
.B(n_71),
.Y(n_6470)
);

AOI21xp5_ASAP7_75t_L g6471 ( 
.A1(n_5870),
.A2(n_3173),
.B(n_3172),
.Y(n_6471)
);

O2A1O1Ixp5_ASAP7_75t_L g6472 ( 
.A1(n_6136),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_6472)
);

HB1xp67_ASAP7_75t_L g6473 ( 
.A(n_6064),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_L g6474 ( 
.A(n_6064),
.B(n_376),
.Y(n_6474)
);

NAND2xp5_ASAP7_75t_L g6475 ( 
.A(n_6082),
.B(n_377),
.Y(n_6475)
);

A2O1A1Ixp33_ASAP7_75t_L g6476 ( 
.A1(n_5833),
.A2(n_74),
.B(n_72),
.C(n_73),
.Y(n_6476)
);

AOI21xp5_ASAP7_75t_L g6477 ( 
.A1(n_5778),
.A2(n_5783),
.B(n_5786),
.Y(n_6477)
);

OAI21xp5_ASAP7_75t_L g6478 ( 
.A1(n_5954),
.A2(n_73),
.B(n_75),
.Y(n_6478)
);

INVx5_ASAP7_75t_L g6479 ( 
.A(n_5881),
.Y(n_6479)
);

BUFx6f_ASAP7_75t_L g6480 ( 
.A(n_5908),
.Y(n_6480)
);

NAND2xp5_ASAP7_75t_SL g6481 ( 
.A(n_5925),
.B(n_2583),
.Y(n_6481)
);

AOI21x1_ASAP7_75t_SL g6482 ( 
.A1(n_6062),
.A2(n_75),
.B(n_76),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6189),
.B(n_76),
.Y(n_6483)
);

INVx4_ASAP7_75t_L g6484 ( 
.A(n_5908),
.Y(n_6484)
);

INVx2_ASAP7_75t_L g6485 ( 
.A(n_6145),
.Y(n_6485)
);

NAND2xp5_ASAP7_75t_L g6486 ( 
.A(n_6082),
.B(n_377),
.Y(n_6486)
);

AOI21xp5_ASAP7_75t_L g6487 ( 
.A1(n_5844),
.A2(n_5808),
.B(n_5874),
.Y(n_6487)
);

BUFx2_ASAP7_75t_L g6488 ( 
.A(n_6109),
.Y(n_6488)
);

OAI21x1_ASAP7_75t_L g6489 ( 
.A1(n_5863),
.A2(n_3686),
.B(n_3685),
.Y(n_6489)
);

AO31x2_ASAP7_75t_L g6490 ( 
.A1(n_5977),
.A2(n_3686),
.A3(n_3693),
.B(n_3685),
.Y(n_6490)
);

AOI221x1_ASAP7_75t_L g6491 ( 
.A1(n_5998),
.A2(n_6096),
.B1(n_6093),
.B2(n_5810),
.C(n_6167),
.Y(n_6491)
);

OAI21xp5_ASAP7_75t_L g6492 ( 
.A1(n_5804),
.A2(n_77),
.B(n_78),
.Y(n_6492)
);

NOR2xp33_ASAP7_75t_L g6493 ( 
.A(n_5908),
.B(n_378),
.Y(n_6493)
);

NOR4xp25_ASAP7_75t_L g6494 ( 
.A(n_6135),
.B(n_80),
.C(n_77),
.D(n_79),
.Y(n_6494)
);

NAND3xp33_ASAP7_75t_L g6495 ( 
.A(n_5804),
.B(n_1677),
.C(n_1636),
.Y(n_6495)
);

OAI22xp5_ASAP7_75t_L g6496 ( 
.A1(n_6033),
.A2(n_3302),
.B1(n_3083),
.B2(n_2601),
.Y(n_6496)
);

AOI21xp5_ASAP7_75t_L g6497 ( 
.A1(n_6053),
.A2(n_3179),
.B(n_3173),
.Y(n_6497)
);

AO21x2_ASAP7_75t_L g6498 ( 
.A1(n_6118),
.A2(n_3704),
.B(n_3693),
.Y(n_6498)
);

AOI21xp5_ASAP7_75t_L g6499 ( 
.A1(n_5797),
.A2(n_5813),
.B(n_5807),
.Y(n_6499)
);

OAI21x1_ASAP7_75t_L g6500 ( 
.A1(n_5867),
.A2(n_3710),
.B(n_3704),
.Y(n_6500)
);

AOI21xp5_ASAP7_75t_L g6501 ( 
.A1(n_5822),
.A2(n_5824),
.B(n_5892),
.Y(n_6501)
);

INVx2_ASAP7_75t_SL g6502 ( 
.A(n_5953),
.Y(n_6502)
);

INVx3_ASAP7_75t_L g6503 ( 
.A(n_6109),
.Y(n_6503)
);

OAI21xp5_ASAP7_75t_L g6504 ( 
.A1(n_6052),
.A2(n_77),
.B(n_79),
.Y(n_6504)
);

BUFx6f_ASAP7_75t_L g6505 ( 
.A(n_5953),
.Y(n_6505)
);

AOI21xp5_ASAP7_75t_L g6506 ( 
.A1(n_5905),
.A2(n_3188),
.B(n_3179),
.Y(n_6506)
);

NOR4xp25_ASAP7_75t_L g6507 ( 
.A(n_5765),
.B(n_81),
.C(n_79),
.D(n_80),
.Y(n_6507)
);

OAI21x1_ASAP7_75t_L g6508 ( 
.A1(n_6168),
.A2(n_3716),
.B(n_3710),
.Y(n_6508)
);

NAND2xp5_ASAP7_75t_L g6509 ( 
.A(n_6179),
.B(n_379),
.Y(n_6509)
);

OA21x2_ASAP7_75t_L g6510 ( 
.A1(n_6038),
.A2(n_3722),
.B(n_3716),
.Y(n_6510)
);

OAI22xp5_ASAP7_75t_L g6511 ( 
.A1(n_6052),
.A2(n_5952),
.B1(n_6003),
.B2(n_5765),
.Y(n_6511)
);

INVx2_ASAP7_75t_L g6512 ( 
.A(n_6145),
.Y(n_6512)
);

NAND2xp5_ASAP7_75t_L g6513 ( 
.A(n_6183),
.B(n_382),
.Y(n_6513)
);

A2O1A1Ixp33_ASAP7_75t_L g6514 ( 
.A1(n_6013),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_6514)
);

INVx3_ASAP7_75t_L g6515 ( 
.A(n_5923),
.Y(n_6515)
);

OAI21x1_ASAP7_75t_L g6516 ( 
.A1(n_5901),
.A2(n_3724),
.B(n_3722),
.Y(n_6516)
);

OAI22xp33_ASAP7_75t_L g6517 ( 
.A1(n_5811),
.A2(n_3728),
.B1(n_3724),
.B2(n_2628),
.Y(n_6517)
);

CKINVDCx5p33_ASAP7_75t_R g6518 ( 
.A(n_5953),
.Y(n_6518)
);

AOI21xp5_ASAP7_75t_SL g6519 ( 
.A1(n_5949),
.A2(n_2628),
.B(n_2601),
.Y(n_6519)
);

OAI21x1_ASAP7_75t_L g6520 ( 
.A1(n_6099),
.A2(n_3728),
.B(n_3044),
.Y(n_6520)
);

OAI21x1_ASAP7_75t_L g6521 ( 
.A1(n_6115),
.A2(n_3044),
.B(n_3043),
.Y(n_6521)
);

NOR2xp33_ASAP7_75t_L g6522 ( 
.A(n_6060),
.B(n_382),
.Y(n_6522)
);

OA21x2_ASAP7_75t_L g6523 ( 
.A1(n_6068),
.A2(n_3048),
.B(n_3043),
.Y(n_6523)
);

AOI21xp5_ASAP7_75t_L g6524 ( 
.A1(n_5847),
.A2(n_3191),
.B(n_3188),
.Y(n_6524)
);

NAND2xp5_ASAP7_75t_L g6525 ( 
.A(n_6170),
.B(n_384),
.Y(n_6525)
);

OAI22xp5_ASAP7_75t_L g6526 ( 
.A1(n_5952),
.A2(n_6003),
.B1(n_6094),
.B2(n_6009),
.Y(n_6526)
);

AND2x2_ASAP7_75t_L g6527 ( 
.A(n_6189),
.B(n_81),
.Y(n_6527)
);

INVx1_ASAP7_75t_L g6528 ( 
.A(n_6145),
.Y(n_6528)
);

OR2x2_ASAP7_75t_L g6529 ( 
.A(n_5937),
.B(n_83),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_6170),
.B(n_384),
.Y(n_6530)
);

AND2x4_ASAP7_75t_L g6531 ( 
.A(n_5997),
.B(n_83),
.Y(n_6531)
);

NAND2xp5_ASAP7_75t_L g6532 ( 
.A(n_6170),
.B(n_385),
.Y(n_6532)
);

INVx1_ASAP7_75t_L g6533 ( 
.A(n_6164),
.Y(n_6533)
);

NOR2x1_ASAP7_75t_SL g6534 ( 
.A(n_6181),
.B(n_1636),
.Y(n_6534)
);

AO22x2_ASAP7_75t_L g6535 ( 
.A1(n_5831),
.A2(n_3048),
.B1(n_3083),
.B2(n_3191),
.Y(n_6535)
);

BUFx4f_ASAP7_75t_L g6536 ( 
.A(n_6060),
.Y(n_6536)
);

INVx1_ASAP7_75t_L g6537 ( 
.A(n_6164),
.Y(n_6537)
);

AND2x4_ASAP7_75t_L g6538 ( 
.A(n_6181),
.B(n_84),
.Y(n_6538)
);

BUFx4_ASAP7_75t_SL g6539 ( 
.A(n_5876),
.Y(n_6539)
);

OAI22xp5_ASAP7_75t_L g6540 ( 
.A1(n_6009),
.A2(n_3302),
.B1(n_2601),
.B2(n_2634),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6164),
.Y(n_6541)
);

OAI21x1_ASAP7_75t_L g6542 ( 
.A1(n_6132),
.A2(n_3090),
.B(n_3193),
.Y(n_6542)
);

NOR2xp33_ASAP7_75t_L g6543 ( 
.A(n_6060),
.B(n_386),
.Y(n_6543)
);

AOI21xp5_ASAP7_75t_L g6544 ( 
.A1(n_5864),
.A2(n_3194),
.B(n_3193),
.Y(n_6544)
);

OAI21x1_ASAP7_75t_L g6545 ( 
.A1(n_5945),
.A2(n_3090),
.B(n_3194),
.Y(n_6545)
);

BUFx12f_ASAP7_75t_L g6546 ( 
.A(n_6090),
.Y(n_6546)
);

OAI22xp5_ASAP7_75t_L g6547 ( 
.A1(n_5811),
.A2(n_2628),
.B1(n_2634),
.B2(n_2690),
.Y(n_6547)
);

O2A1O1Ixp33_ASAP7_75t_SL g6548 ( 
.A1(n_5966),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_6548)
);

CKINVDCx20_ASAP7_75t_R g6549 ( 
.A(n_6150),
.Y(n_6549)
);

O2A1O1Ixp5_ASAP7_75t_SL g6550 ( 
.A1(n_5943),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_6550)
);

INVx1_ASAP7_75t_L g6551 ( 
.A(n_6102),
.Y(n_6551)
);

OAI22xp33_ASAP7_75t_L g6552 ( 
.A1(n_6181),
.A2(n_2634),
.B1(n_2690),
.B2(n_3195),
.Y(n_6552)
);

AOI21xp5_ASAP7_75t_L g6553 ( 
.A1(n_5873),
.A2(n_3196),
.B(n_3195),
.Y(n_6553)
);

INVx1_ASAP7_75t_L g6554 ( 
.A(n_6102),
.Y(n_6554)
);

AOI21xp5_ASAP7_75t_L g6555 ( 
.A1(n_6022),
.A2(n_3197),
.B(n_3196),
.Y(n_6555)
);

AOI21xp33_ASAP7_75t_L g6556 ( 
.A1(n_6195),
.A2(n_87),
.B(n_88),
.Y(n_6556)
);

NAND2xp5_ASAP7_75t_L g6557 ( 
.A(n_6170),
.B(n_386),
.Y(n_6557)
);

A2O1A1Ixp33_ASAP7_75t_L g6558 ( 
.A1(n_5787),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_6558)
);

AO31x2_ASAP7_75t_L g6559 ( 
.A1(n_5904),
.A2(n_3205),
.A3(n_3207),
.B(n_3197),
.Y(n_6559)
);

O2A1O1Ixp33_ASAP7_75t_SL g6560 ( 
.A1(n_6121),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_6560)
);

INVx2_ASAP7_75t_L g6561 ( 
.A(n_6102),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_6137),
.Y(n_6562)
);

AOI21xp5_ASAP7_75t_L g6563 ( 
.A1(n_5880),
.A2(n_5882),
.B(n_6077),
.Y(n_6563)
);

OA22x2_ASAP7_75t_L g6564 ( 
.A1(n_6158),
.A2(n_3207),
.B1(n_3211),
.B2(n_3205),
.Y(n_6564)
);

AND2x4_ASAP7_75t_L g6565 ( 
.A(n_5989),
.B(n_90),
.Y(n_6565)
);

BUFx2_ASAP7_75t_L g6566 ( 
.A(n_6473),
.Y(n_6566)
);

OAI21x1_ASAP7_75t_L g6567 ( 
.A1(n_6223),
.A2(n_6116),
.B(n_5924),
.Y(n_6567)
);

AO21x2_ASAP7_75t_L g6568 ( 
.A1(n_6447),
.A2(n_6455),
.B(n_6382),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6199),
.Y(n_6569)
);

OA21x2_ASAP7_75t_L g6570 ( 
.A1(n_6209),
.A2(n_6000),
.B(n_6055),
.Y(n_6570)
);

BUFx2_ASAP7_75t_SL g6571 ( 
.A(n_6334),
.Y(n_6571)
);

AOI22xp5_ASAP7_75t_L g6572 ( 
.A1(n_6511),
.A2(n_5856),
.B1(n_5938),
.B2(n_5912),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6336),
.Y(n_6573)
);

OAI21x1_ASAP7_75t_L g6574 ( 
.A1(n_6243),
.A2(n_5955),
.B(n_5926),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_6234),
.Y(n_6575)
);

OAI21x1_ASAP7_75t_L g6576 ( 
.A1(n_6295),
.A2(n_5921),
.B(n_5911),
.Y(n_6576)
);

AOI21xp5_ASAP7_75t_L g6577 ( 
.A1(n_6487),
.A2(n_5912),
.B(n_5856),
.Y(n_6577)
);

BUFx3_ASAP7_75t_L g6578 ( 
.A(n_6267),
.Y(n_6578)
);

AO21x1_ASAP7_75t_L g6579 ( 
.A1(n_6529),
.A2(n_6526),
.B(n_6296),
.Y(n_6579)
);

INVx2_ASAP7_75t_L g6580 ( 
.A(n_6428),
.Y(n_6580)
);

INVx6_ASAP7_75t_L g6581 ( 
.A(n_6221),
.Y(n_6581)
);

HB1xp67_ASAP7_75t_L g6582 ( 
.A(n_6421),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6236),
.Y(n_6583)
);

OAI21x1_ASAP7_75t_L g6584 ( 
.A1(n_6233),
.A2(n_5978),
.B(n_5928),
.Y(n_6584)
);

INVx1_ASAP7_75t_L g6585 ( 
.A(n_6241),
.Y(n_6585)
);

OAI21x1_ASAP7_75t_L g6586 ( 
.A1(n_6499),
.A2(n_5991),
.B(n_6144),
.Y(n_6586)
);

OA21x2_ASAP7_75t_L g6587 ( 
.A1(n_6462),
.A2(n_6045),
.B(n_6001),
.Y(n_6587)
);

CKINVDCx5p33_ASAP7_75t_R g6588 ( 
.A(n_6240),
.Y(n_6588)
);

INVx6_ASAP7_75t_L g6589 ( 
.A(n_6211),
.Y(n_6589)
);

INVx4_ASAP7_75t_L g6590 ( 
.A(n_6430),
.Y(n_6590)
);

AO21x2_ASAP7_75t_L g6591 ( 
.A1(n_6528),
.A2(n_6155),
.B(n_6027),
.Y(n_6591)
);

OAI21x1_ASAP7_75t_L g6592 ( 
.A1(n_6330),
.A2(n_5859),
.B(n_6081),
.Y(n_6592)
);

INVx1_ASAP7_75t_L g6593 ( 
.A(n_6266),
.Y(n_6593)
);

OAI21x1_ASAP7_75t_L g6594 ( 
.A1(n_6459),
.A2(n_6083),
.B(n_6047),
.Y(n_6594)
);

AOI221xp5_ASAP7_75t_L g6595 ( 
.A1(n_6377),
.A2(n_5938),
.B1(n_5972),
.B2(n_6176),
.C(n_6172),
.Y(n_6595)
);

OAI21x1_ASAP7_75t_L g6596 ( 
.A1(n_6501),
.A2(n_5949),
.B(n_6076),
.Y(n_6596)
);

OAI21x1_ASAP7_75t_L g6597 ( 
.A1(n_6477),
.A2(n_6432),
.B(n_6563),
.Y(n_6597)
);

INVx1_ASAP7_75t_SL g6598 ( 
.A(n_6539),
.Y(n_6598)
);

OAI21x1_ASAP7_75t_L g6599 ( 
.A1(n_6421),
.A2(n_5976),
.B(n_5964),
.Y(n_6599)
);

AO31x2_ASAP7_75t_L g6600 ( 
.A1(n_6411),
.A2(n_5906),
.A3(n_5890),
.B(n_5879),
.Y(n_6600)
);

OAI21x1_ASAP7_75t_L g6601 ( 
.A1(n_6345),
.A2(n_5930),
.B(n_6084),
.Y(n_6601)
);

OA21x2_ASAP7_75t_L g6602 ( 
.A1(n_6207),
.A2(n_6491),
.B(n_6533),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_6428),
.Y(n_6603)
);

AO21x2_ASAP7_75t_L g6604 ( 
.A1(n_6537),
.A2(n_6155),
.B(n_6050),
.Y(n_6604)
);

AND2x4_ASAP7_75t_L g6605 ( 
.A(n_6298),
.B(n_5937),
.Y(n_6605)
);

AOI21xp5_ASAP7_75t_L g6606 ( 
.A1(n_6278),
.A2(n_6019),
.B(n_6004),
.Y(n_6606)
);

NAND2xp5_ASAP7_75t_L g6607 ( 
.A(n_6355),
.B(n_5849),
.Y(n_6607)
);

BUFx2_ASAP7_75t_R g6608 ( 
.A(n_6392),
.Y(n_6608)
);

OAI21x1_ASAP7_75t_SL g6609 ( 
.A1(n_6255),
.A2(n_5839),
.B(n_6028),
.Y(n_6609)
);

OAI21x1_ASAP7_75t_L g6610 ( 
.A1(n_6210),
.A2(n_6084),
.B(n_6174),
.Y(n_6610)
);

OAI21xp5_ASAP7_75t_L g6611 ( 
.A1(n_6197),
.A2(n_5814),
.B(n_6172),
.Y(n_6611)
);

NAND2xp5_ASAP7_75t_L g6612 ( 
.A(n_6208),
.B(n_5849),
.Y(n_6612)
);

BUFx3_ASAP7_75t_L g6613 ( 
.A(n_6276),
.Y(n_6613)
);

OAI21x1_ASAP7_75t_L g6614 ( 
.A1(n_6198),
.A2(n_6174),
.B(n_6018),
.Y(n_6614)
);

OAI21x1_ASAP7_75t_L g6615 ( 
.A1(n_6245),
.A2(n_5979),
.B(n_6120),
.Y(n_6615)
);

OAI21x1_ASAP7_75t_L g6616 ( 
.A1(n_6291),
.A2(n_6129),
.B(n_6125),
.Y(n_6616)
);

OA21x2_ASAP7_75t_L g6617 ( 
.A1(n_6541),
.A2(n_6194),
.B(n_6147),
.Y(n_6617)
);

HB1xp67_ASAP7_75t_L g6618 ( 
.A(n_6271),
.Y(n_6618)
);

HB1xp67_ASAP7_75t_L g6619 ( 
.A(n_6229),
.Y(n_6619)
);

BUFx2_ASAP7_75t_L g6620 ( 
.A(n_6248),
.Y(n_6620)
);

NAND2x1p5_ASAP7_75t_L g6621 ( 
.A(n_6213),
.B(n_5907),
.Y(n_6621)
);

BUFx2_ASAP7_75t_L g6622 ( 
.A(n_6248),
.Y(n_6622)
);

INVx3_ASAP7_75t_L g6623 ( 
.A(n_6335),
.Y(n_6623)
);

OAI21x1_ASAP7_75t_L g6624 ( 
.A1(n_6292),
.A2(n_6125),
.B(n_6124),
.Y(n_6624)
);

AND2x4_ASAP7_75t_L g6625 ( 
.A(n_6398),
.B(n_5937),
.Y(n_6625)
);

AND2x2_ASAP7_75t_L g6626 ( 
.A(n_6307),
.B(n_6150),
.Y(n_6626)
);

AO21x2_ASAP7_75t_L g6627 ( 
.A1(n_6405),
.A2(n_6050),
.B(n_6037),
.Y(n_6627)
);

AND2x4_ASAP7_75t_L g6628 ( 
.A(n_6250),
.B(n_5907),
.Y(n_6628)
);

AND3x2_ASAP7_75t_L g6629 ( 
.A(n_6538),
.B(n_6031),
.C(n_6028),
.Y(n_6629)
);

OAI21x1_ASAP7_75t_L g6630 ( 
.A1(n_6408),
.A2(n_6124),
.B(n_6086),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_L g6631 ( 
.A(n_6275),
.B(n_5849),
.Y(n_6631)
);

OAI21x1_ASAP7_75t_L g6632 ( 
.A1(n_6235),
.A2(n_6159),
.B(n_6156),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6306),
.Y(n_6633)
);

AO21x2_ASAP7_75t_L g6634 ( 
.A1(n_6551),
.A2(n_6037),
.B(n_5839),
.Y(n_6634)
);

BUFx2_ASAP7_75t_SL g6635 ( 
.A(n_6549),
.Y(n_6635)
);

BUFx12f_ASAP7_75t_L g6636 ( 
.A(n_6211),
.Y(n_6636)
);

INVx1_ASAP7_75t_L g6637 ( 
.A(n_6321),
.Y(n_6637)
);

AO21x2_ASAP7_75t_L g6638 ( 
.A1(n_6554),
.A2(n_6031),
.B(n_6098),
.Y(n_6638)
);

AND2x4_ASAP7_75t_L g6639 ( 
.A(n_6335),
.B(n_5894),
.Y(n_6639)
);

OAI21x1_ASAP7_75t_L g6640 ( 
.A1(n_6217),
.A2(n_6142),
.B(n_5829),
.Y(n_6640)
);

BUFx2_ASAP7_75t_L g6641 ( 
.A(n_6385),
.Y(n_6641)
);

OA21x2_ASAP7_75t_L g6642 ( 
.A1(n_6562),
.A2(n_6146),
.B(n_6092),
.Y(n_6642)
);

BUFx2_ASAP7_75t_SL g6643 ( 
.A(n_6323),
.Y(n_6643)
);

NAND2x1p5_ASAP7_75t_L g6644 ( 
.A(n_6213),
.B(n_6042),
.Y(n_6644)
);

INVx1_ASAP7_75t_L g6645 ( 
.A(n_6339),
.Y(n_6645)
);

OAI21x1_ASAP7_75t_L g6646 ( 
.A1(n_6282),
.A2(n_6087),
.B(n_6143),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6340),
.Y(n_6647)
);

CKINVDCx20_ASAP7_75t_R g6648 ( 
.A(n_6433),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6354),
.Y(n_6649)
);

NAND2xp5_ASAP7_75t_L g6650 ( 
.A(n_6259),
.B(n_5894),
.Y(n_6650)
);

AND2x4_ASAP7_75t_L g6651 ( 
.A(n_6385),
.B(n_5894),
.Y(n_6651)
);

BUFx3_ASAP7_75t_L g6652 ( 
.A(n_6346),
.Y(n_6652)
);

NAND2x1p5_ASAP7_75t_L g6653 ( 
.A(n_6213),
.B(n_6131),
.Y(n_6653)
);

AO21x2_ASAP7_75t_L g6654 ( 
.A1(n_6387),
.A2(n_6141),
.B(n_6191),
.Y(n_6654)
);

BUFx3_ASAP7_75t_L g6655 ( 
.A(n_6434),
.Y(n_6655)
);

INVx1_ASAP7_75t_L g6656 ( 
.A(n_6311),
.Y(n_6656)
);

BUFx2_ASAP7_75t_L g6657 ( 
.A(n_6488),
.Y(n_6657)
);

OR3x4_ASAP7_75t_SL g6658 ( 
.A(n_6232),
.B(n_90),
.C(n_91),
.Y(n_6658)
);

AND2x4_ASAP7_75t_L g6659 ( 
.A(n_6394),
.B(n_6040),
.Y(n_6659)
);

OA21x2_ASAP7_75t_L g6660 ( 
.A1(n_6485),
.A2(n_6153),
.B(n_6152),
.Y(n_6660)
);

NAND2x1p5_ASAP7_75t_L g6661 ( 
.A(n_6239),
.B(n_6173),
.Y(n_6661)
);

AND2x4_ASAP7_75t_L g6662 ( 
.A(n_6394),
.B(n_6040),
.Y(n_6662)
);

OAI21x1_ASAP7_75t_L g6663 ( 
.A1(n_6389),
.A2(n_6143),
.B(n_6148),
.Y(n_6663)
);

AOI21xp5_ASAP7_75t_L g6664 ( 
.A1(n_6277),
.A2(n_5939),
.B(n_6160),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_6383),
.Y(n_6665)
);

BUFx2_ASAP7_75t_L g6666 ( 
.A(n_6518),
.Y(n_6666)
);

CKINVDCx11_ASAP7_75t_R g6667 ( 
.A(n_6454),
.Y(n_6667)
);

NAND2xp5_ASAP7_75t_L g6668 ( 
.A(n_6220),
.B(n_5825),
.Y(n_6668)
);

OR2x6_ASAP7_75t_L g6669 ( 
.A(n_6205),
.B(n_6176),
.Y(n_6669)
);

OAI21x1_ASAP7_75t_L g6670 ( 
.A1(n_6429),
.A2(n_5932),
.B(n_6141),
.Y(n_6670)
);

OAI21xp33_ASAP7_75t_SL g6671 ( 
.A1(n_6440),
.A2(n_5974),
.B(n_5963),
.Y(n_6671)
);

OA21x2_ASAP7_75t_L g6672 ( 
.A1(n_6512),
.A2(n_6182),
.B(n_6073),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6463),
.Y(n_6673)
);

OAI21x1_ASAP7_75t_SL g6674 ( 
.A1(n_6299),
.A2(n_5940),
.B(n_5809),
.Y(n_6674)
);

INVx2_ASAP7_75t_L g6675 ( 
.A(n_6428),
.Y(n_6675)
);

NAND2xp5_ASAP7_75t_L g6676 ( 
.A(n_6220),
.B(n_5825),
.Y(n_6676)
);

OAI21x1_ASAP7_75t_L g6677 ( 
.A1(n_6429),
.A2(n_6182),
.B(n_5993),
.Y(n_6677)
);

BUFx3_ASAP7_75t_L g6678 ( 
.A(n_6196),
.Y(n_6678)
);

OAI21x1_ASAP7_75t_L g6679 ( 
.A1(n_6230),
.A2(n_6191),
.B(n_5825),
.Y(n_6679)
);

BUFx6f_ASAP7_75t_L g6680 ( 
.A(n_6372),
.Y(n_6680)
);

AOI21xp5_ASAP7_75t_L g6681 ( 
.A1(n_6358),
.A2(n_6215),
.B(n_6264),
.Y(n_6681)
);

BUFx12f_ASAP7_75t_L g6682 ( 
.A(n_6262),
.Y(n_6682)
);

CKINVDCx6p67_ASAP7_75t_R g6683 ( 
.A(n_6309),
.Y(n_6683)
);

BUFx6f_ASAP7_75t_L g6684 ( 
.A(n_6372),
.Y(n_6684)
);

NOR2xp33_ASAP7_75t_L g6685 ( 
.A(n_6324),
.B(n_387),
.Y(n_6685)
);

AO21x2_ASAP7_75t_L g6686 ( 
.A1(n_6397),
.A2(n_6040),
.B(n_6137),
.Y(n_6686)
);

INVx2_ASAP7_75t_L g6687 ( 
.A(n_6326),
.Y(n_6687)
);

INVx6_ASAP7_75t_SL g6688 ( 
.A(n_6538),
.Y(n_6688)
);

OA21x2_ASAP7_75t_L g6689 ( 
.A1(n_6561),
.A2(n_6137),
.B(n_3215),
.Y(n_6689)
);

OAI21x1_ASAP7_75t_L g6690 ( 
.A1(n_6564),
.A2(n_3090),
.B(n_3211),
.Y(n_6690)
);

HB1xp67_ASAP7_75t_L g6691 ( 
.A(n_6318),
.Y(n_6691)
);

AO21x1_ASAP7_75t_L g6692 ( 
.A1(n_6313),
.A2(n_91),
.B(n_92),
.Y(n_6692)
);

CKINVDCx5p33_ASAP7_75t_R g6693 ( 
.A(n_6384),
.Y(n_6693)
);

OR2x2_ASAP7_75t_L g6694 ( 
.A(n_6425),
.B(n_6465),
.Y(n_6694)
);

INVx1_ASAP7_75t_L g6695 ( 
.A(n_6427),
.Y(n_6695)
);

AOI21x1_ASAP7_75t_SL g6696 ( 
.A1(n_6301),
.A2(n_93),
.B(n_94),
.Y(n_6696)
);

NAND2x1p5_ASAP7_75t_L g6697 ( 
.A(n_6239),
.B(n_3292),
.Y(n_6697)
);

BUFx2_ASAP7_75t_L g6698 ( 
.A(n_6503),
.Y(n_6698)
);

NAND2x1p5_ASAP7_75t_L g6699 ( 
.A(n_6239),
.B(n_3292),
.Y(n_6699)
);

AND2x4_ASAP7_75t_L g6700 ( 
.A(n_6531),
.B(n_93),
.Y(n_6700)
);

NAND2x1p5_ASAP7_75t_L g6701 ( 
.A(n_6342),
.B(n_3292),
.Y(n_6701)
);

AO21x2_ASAP7_75t_L g6702 ( 
.A1(n_6325),
.A2(n_6327),
.B(n_6315),
.Y(n_6702)
);

AO21x1_ASAP7_75t_L g6703 ( 
.A1(n_6224),
.A2(n_94),
.B(n_95),
.Y(n_6703)
);

NAND2xp5_ASAP7_75t_L g6704 ( 
.A(n_6204),
.B(n_95),
.Y(n_6704)
);

AO21x2_ASAP7_75t_L g6705 ( 
.A1(n_6347),
.A2(n_3219),
.B(n_3215),
.Y(n_6705)
);

INVxp67_ASAP7_75t_SL g6706 ( 
.A(n_6204),
.Y(n_6706)
);

NAND2xp5_ASAP7_75t_L g6707 ( 
.A(n_6281),
.B(n_96),
.Y(n_6707)
);

OAI22x1_ASAP7_75t_L g6708 ( 
.A1(n_6531),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_6708)
);

CKINVDCx5p33_ASAP7_75t_R g6709 ( 
.A(n_6361),
.Y(n_6709)
);

INVx1_ASAP7_75t_L g6710 ( 
.A(n_6344),
.Y(n_6710)
);

OAI21x1_ASAP7_75t_L g6711 ( 
.A1(n_6515),
.A2(n_3231),
.B(n_3230),
.Y(n_6711)
);

OAI21x1_ASAP7_75t_L g6712 ( 
.A1(n_6515),
.A2(n_3231),
.B(n_3230),
.Y(n_6712)
);

INVx3_ASAP7_75t_L g6713 ( 
.A(n_6503),
.Y(n_6713)
);

AOI21xp5_ASAP7_75t_L g6714 ( 
.A1(n_6274),
.A2(n_3221),
.B(n_3219),
.Y(n_6714)
);

AOI22x1_ASAP7_75t_L g6715 ( 
.A1(n_6218),
.A2(n_99),
.B1(n_96),
.B2(n_98),
.Y(n_6715)
);

BUFx3_ASAP7_75t_L g6716 ( 
.A(n_6391),
.Y(n_6716)
);

OR2x2_ASAP7_75t_L g6717 ( 
.A(n_6257),
.B(n_98),
.Y(n_6717)
);

NOR2xp33_ASAP7_75t_L g6718 ( 
.A(n_6269),
.B(n_387),
.Y(n_6718)
);

OAI21x1_ASAP7_75t_L g6719 ( 
.A1(n_6222),
.A2(n_3223),
.B(n_3221),
.Y(n_6719)
);

OAI21x1_ASAP7_75t_L g6720 ( 
.A1(n_6364),
.A2(n_3226),
.B(n_3223),
.Y(n_6720)
);

AOI21xp5_ASAP7_75t_L g6721 ( 
.A1(n_6343),
.A2(n_3226),
.B(n_3156),
.Y(n_6721)
);

NAND3xp33_ASAP7_75t_L g6722 ( 
.A(n_6349),
.B(n_6193),
.C(n_1677),
.Y(n_6722)
);

BUFx2_ASAP7_75t_L g6723 ( 
.A(n_6224),
.Y(n_6723)
);

OA21x2_ASAP7_75t_L g6724 ( 
.A1(n_6303),
.A2(n_99),
.B(n_100),
.Y(n_6724)
);

OAI21x1_ASAP7_75t_L g6725 ( 
.A1(n_6279),
.A2(n_2546),
.B(n_2477),
.Y(n_6725)
);

OA21x2_ASAP7_75t_L g6726 ( 
.A1(n_6449),
.A2(n_100),
.B(n_101),
.Y(n_6726)
);

BUFx2_ASAP7_75t_L g6727 ( 
.A(n_6265),
.Y(n_6727)
);

NAND2x1p5_ASAP7_75t_L g6728 ( 
.A(n_6342),
.B(n_3292),
.Y(n_6728)
);

OAI21x1_ASAP7_75t_L g6729 ( 
.A1(n_6356),
.A2(n_6341),
.B(n_6329),
.Y(n_6729)
);

AO31x2_ASAP7_75t_L g6730 ( 
.A1(n_6457),
.A2(n_102),
.A3(n_100),
.B(n_101),
.Y(n_6730)
);

AOI22xp33_ASAP7_75t_L g6731 ( 
.A1(n_6246),
.A2(n_2634),
.B1(n_2690),
.B2(n_2895),
.Y(n_6731)
);

CKINVDCx5p33_ASAP7_75t_R g6732 ( 
.A(n_6283),
.Y(n_6732)
);

INVx1_ASAP7_75t_L g6733 ( 
.A(n_6373),
.Y(n_6733)
);

OAI21xp5_ASAP7_75t_L g6734 ( 
.A1(n_6350),
.A2(n_102),
.B(n_103),
.Y(n_6734)
);

HB1xp67_ASAP7_75t_L g6735 ( 
.A(n_6320),
.Y(n_6735)
);

INVx8_ASAP7_75t_L g6736 ( 
.A(n_6227),
.Y(n_6736)
);

INVx1_ASAP7_75t_L g6737 ( 
.A(n_6379),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6380),
.Y(n_6738)
);

OAI21x1_ASAP7_75t_L g6739 ( 
.A1(n_6328),
.A2(n_2674),
.B(n_2558),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6426),
.Y(n_6740)
);

OA21x2_ASAP7_75t_L g6741 ( 
.A1(n_6261),
.A2(n_102),
.B(n_103),
.Y(n_6741)
);

INVx3_ASAP7_75t_SL g6742 ( 
.A(n_6265),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6502),
.B(n_103),
.Y(n_6743)
);

NOR2xp33_ASAP7_75t_L g6744 ( 
.A(n_6254),
.B(n_388),
.Y(n_6744)
);

HB1xp67_ASAP7_75t_L g6745 ( 
.A(n_6225),
.Y(n_6745)
);

OAI21x1_ASAP7_75t_L g6746 ( 
.A1(n_6319),
.A2(n_2989),
.B(n_2963),
.Y(n_6746)
);

OR2x6_ASAP7_75t_L g6747 ( 
.A(n_6205),
.B(n_3292),
.Y(n_6747)
);

INVx2_ASAP7_75t_L g6748 ( 
.A(n_6305),
.Y(n_6748)
);

OAI21x1_ASAP7_75t_L g6749 ( 
.A1(n_6525),
.A2(n_2989),
.B(n_2963),
.Y(n_6749)
);

INVx1_ASAP7_75t_L g6750 ( 
.A(n_6260),
.Y(n_6750)
);

CKINVDCx8_ASAP7_75t_R g6751 ( 
.A(n_6290),
.Y(n_6751)
);

AO31x2_ASAP7_75t_L g6752 ( 
.A1(n_6237),
.A2(n_106),
.A3(n_104),
.B(n_105),
.Y(n_6752)
);

OAI21x1_ASAP7_75t_L g6753 ( 
.A1(n_6530),
.A2(n_6557),
.B(n_6532),
.Y(n_6753)
);

BUFx3_ASAP7_75t_L g6754 ( 
.A(n_6288),
.Y(n_6754)
);

AOI21xp5_ASAP7_75t_L g6755 ( 
.A1(n_6333),
.A2(n_3156),
.B(n_3144),
.Y(n_6755)
);

OAI21x1_ASAP7_75t_L g6756 ( 
.A1(n_6317),
.A2(n_2989),
.B(n_2963),
.Y(n_6756)
);

AO21x2_ASAP7_75t_L g6757 ( 
.A1(n_6322),
.A2(n_3861),
.B(n_104),
.Y(n_6757)
);

NAND2x1_ASAP7_75t_L g6758 ( 
.A(n_6290),
.B(n_1636),
.Y(n_6758)
);

OAI21xp5_ASAP7_75t_L g6759 ( 
.A1(n_6200),
.A2(n_105),
.B(n_106),
.Y(n_6759)
);

OAI21x1_ASAP7_75t_L g6760 ( 
.A1(n_6280),
.A2(n_3051),
.B(n_3020),
.Y(n_6760)
);

OAI21x1_ASAP7_75t_L g6761 ( 
.A1(n_6280),
.A2(n_3051),
.B(n_3020),
.Y(n_6761)
);

OAI21x1_ASAP7_75t_L g6762 ( 
.A1(n_6469),
.A2(n_3051),
.B(n_3020),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_6305),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_6314),
.Y(n_6764)
);

INVx4_ASAP7_75t_L g6765 ( 
.A(n_6372),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6351),
.Y(n_6766)
);

OAI21x1_ASAP7_75t_L g6767 ( 
.A1(n_6489),
.A2(n_3100),
.B(n_3071),
.Y(n_6767)
);

INVx2_ASAP7_75t_L g6768 ( 
.A(n_6225),
.Y(n_6768)
);

BUFx2_ASAP7_75t_SL g6769 ( 
.A(n_6342),
.Y(n_6769)
);

AND2x4_ASAP7_75t_L g6770 ( 
.A(n_6353),
.B(n_107),
.Y(n_6770)
);

AND2x2_ASAP7_75t_L g6771 ( 
.A(n_6352),
.B(n_107),
.Y(n_6771)
);

INVxp67_ASAP7_75t_L g6772 ( 
.A(n_6228),
.Y(n_6772)
);

AND2x4_ASAP7_75t_L g6773 ( 
.A(n_6353),
.B(n_108),
.Y(n_6773)
);

BUFx3_ASAP7_75t_L g6774 ( 
.A(n_6441),
.Y(n_6774)
);

NAND2xp5_ASAP7_75t_L g6775 ( 
.A(n_6225),
.B(n_108),
.Y(n_6775)
);

AO21x2_ASAP7_75t_L g6776 ( 
.A1(n_6419),
.A2(n_3861),
.B(n_108),
.Y(n_6776)
);

BUFx3_ASAP7_75t_L g6777 ( 
.A(n_6470),
.Y(n_6777)
);

BUFx3_ASAP7_75t_L g6778 ( 
.A(n_6422),
.Y(n_6778)
);

OAI21x1_ASAP7_75t_L g6779 ( 
.A1(n_6500),
.A2(n_3149),
.B(n_3100),
.Y(n_6779)
);

AO31x2_ASAP7_75t_L g6780 ( 
.A1(n_6453),
.A2(n_111),
.A3(n_109),
.B(n_110),
.Y(n_6780)
);

OAI21x1_ASAP7_75t_L g6781 ( 
.A1(n_6272),
.A2(n_3149),
.B(n_3100),
.Y(n_6781)
);

INVx6_ASAP7_75t_L g6782 ( 
.A(n_6546),
.Y(n_6782)
);

BUFx2_ASAP7_75t_L g6783 ( 
.A(n_6420),
.Y(n_6783)
);

AO21x2_ASAP7_75t_L g6784 ( 
.A1(n_6424),
.A2(n_3861),
.B(n_109),
.Y(n_6784)
);

NOR2xp33_ASAP7_75t_L g6785 ( 
.A(n_6212),
.B(n_388),
.Y(n_6785)
);

OAI21x1_ASAP7_75t_L g6786 ( 
.A1(n_6359),
.A2(n_3149),
.B(n_3071),
.Y(n_6786)
);

AO21x2_ASAP7_75t_L g6787 ( 
.A1(n_6438),
.A2(n_109),
.B(n_110),
.Y(n_6787)
);

OAI21x1_ASAP7_75t_L g6788 ( 
.A1(n_6448),
.A2(n_3071),
.B(n_110),
.Y(n_6788)
);

BUFx12f_ASAP7_75t_L g6789 ( 
.A(n_6423),
.Y(n_6789)
);

OAI21x1_ASAP7_75t_L g6790 ( 
.A1(n_6331),
.A2(n_111),
.B(n_112),
.Y(n_6790)
);

OA21x2_ASAP7_75t_L g6791 ( 
.A1(n_6297),
.A2(n_111),
.B(n_112),
.Y(n_6791)
);

BUFx2_ASAP7_75t_SL g6792 ( 
.A(n_6353),
.Y(n_6792)
);

OAI22xp5_ASAP7_75t_L g6793 ( 
.A1(n_6476),
.A2(n_6258),
.B1(n_6294),
.B2(n_6268),
.Y(n_6793)
);

INVx2_ASAP7_75t_L g6794 ( 
.A(n_6396),
.Y(n_6794)
);

INVx2_ASAP7_75t_L g6795 ( 
.A(n_6396),
.Y(n_6795)
);

OAI21x1_ASAP7_75t_L g6796 ( 
.A1(n_6406),
.A2(n_112),
.B(n_113),
.Y(n_6796)
);

HB1xp67_ASAP7_75t_L g6797 ( 
.A(n_6401),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_L g6798 ( 
.A(n_6238),
.B(n_6293),
.Y(n_6798)
);

OAI21x1_ASAP7_75t_L g6799 ( 
.A1(n_6520),
.A2(n_6521),
.B(n_6253),
.Y(n_6799)
);

OAI21x1_ASAP7_75t_L g6800 ( 
.A1(n_6400),
.A2(n_115),
.B(n_116),
.Y(n_6800)
);

NAND2xp5_ASAP7_75t_SL g6801 ( 
.A(n_6480),
.B(n_1636),
.Y(n_6801)
);

INVx8_ASAP7_75t_L g6802 ( 
.A(n_6227),
.Y(n_6802)
);

AND2x4_ASAP7_75t_L g6803 ( 
.A(n_6565),
.B(n_115),
.Y(n_6803)
);

OAI21x1_ASAP7_75t_L g6804 ( 
.A1(n_6201),
.A2(n_6302),
.B(n_6231),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_L g6805 ( 
.A(n_6338),
.B(n_115),
.Y(n_6805)
);

INVx1_ASAP7_75t_SL g6806 ( 
.A(n_6483),
.Y(n_6806)
);

OA21x2_ASAP7_75t_L g6807 ( 
.A1(n_6381),
.A2(n_116),
.B(n_117),
.Y(n_6807)
);

OAI21x1_ASAP7_75t_L g6808 ( 
.A1(n_6252),
.A2(n_116),
.B(n_117),
.Y(n_6808)
);

INVx2_ASAP7_75t_L g6809 ( 
.A(n_6396),
.Y(n_6809)
);

OAI21x1_ASAP7_75t_L g6810 ( 
.A1(n_6510),
.A2(n_117),
.B(n_118),
.Y(n_6810)
);

INVx2_ASAP7_75t_L g6811 ( 
.A(n_6399),
.Y(n_6811)
);

INVx2_ASAP7_75t_SL g6812 ( 
.A(n_6527),
.Y(n_6812)
);

CKINVDCx20_ASAP7_75t_R g6813 ( 
.A(n_6509),
.Y(n_6813)
);

CKINVDCx6p67_ASAP7_75t_R g6814 ( 
.A(n_6378),
.Y(n_6814)
);

INVx2_ASAP7_75t_L g6815 ( 
.A(n_6399),
.Y(n_6815)
);

OA21x2_ASAP7_75t_L g6816 ( 
.A1(n_6474),
.A2(n_118),
.B(n_119),
.Y(n_6816)
);

OAI21xp5_ASAP7_75t_L g6817 ( 
.A1(n_6507),
.A2(n_118),
.B(n_119),
.Y(n_6817)
);

INVx2_ASAP7_75t_L g6818 ( 
.A(n_6399),
.Y(n_6818)
);

INVx2_ASAP7_75t_L g6819 ( 
.A(n_6407),
.Y(n_6819)
);

INVx1_ASAP7_75t_L g6820 ( 
.A(n_6304),
.Y(n_6820)
);

NAND3xp33_ASAP7_75t_L g6821 ( 
.A(n_6286),
.B(n_1678),
.C(n_1677),
.Y(n_6821)
);

OR2x6_ASAP7_75t_L g6822 ( 
.A(n_6202),
.B(n_3335),
.Y(n_6822)
);

AND2x2_ASAP7_75t_L g6823 ( 
.A(n_6352),
.B(n_119),
.Y(n_6823)
);

OAI21x1_ASAP7_75t_L g6824 ( 
.A1(n_6510),
.A2(n_120),
.B(n_121),
.Y(n_6824)
);

AO21x2_ASAP7_75t_L g6825 ( 
.A1(n_6556),
.A2(n_120),
.B(n_121),
.Y(n_6825)
);

INVx2_ASAP7_75t_L g6826 ( 
.A(n_6407),
.Y(n_6826)
);

AO21x1_ASAP7_75t_L g6827 ( 
.A1(n_6414),
.A2(n_6416),
.B(n_6247),
.Y(n_6827)
);

BUFx4f_ASAP7_75t_SL g6828 ( 
.A(n_6480),
.Y(n_6828)
);

NAND2x1p5_ASAP7_75t_L g6829 ( 
.A(n_6410),
.B(n_6479),
.Y(n_6829)
);

INVx2_ASAP7_75t_SL g6830 ( 
.A(n_6410),
.Y(n_6830)
);

BUFx3_ASAP7_75t_L g6831 ( 
.A(n_6513),
.Y(n_6831)
);

AND2x4_ASAP7_75t_L g6832 ( 
.A(n_6565),
.B(n_120),
.Y(n_6832)
);

INVx2_ASAP7_75t_L g6833 ( 
.A(n_6407),
.Y(n_6833)
);

NOR2xp33_ASAP7_75t_L g6834 ( 
.A(n_6418),
.B(n_389),
.Y(n_6834)
);

OAI21x1_ASAP7_75t_L g6835 ( 
.A1(n_6542),
.A2(n_121),
.B(n_122),
.Y(n_6835)
);

AOI21x1_ASAP7_75t_L g6836 ( 
.A1(n_6475),
.A2(n_122),
.B(n_123),
.Y(n_6836)
);

BUFx12f_ASAP7_75t_L g6837 ( 
.A(n_6480),
.Y(n_6837)
);

NOR2xp33_ASAP7_75t_L g6838 ( 
.A(n_6442),
.B(n_389),
.Y(n_6838)
);

OAI21xp5_ASAP7_75t_L g6839 ( 
.A1(n_6494),
.A2(n_123),
.B(n_124),
.Y(n_6839)
);

AOI22xp33_ASAP7_75t_L g6840 ( 
.A1(n_6504),
.A2(n_2690),
.B1(n_2959),
.B2(n_2895),
.Y(n_6840)
);

CKINVDCx5p33_ASAP7_75t_R g6841 ( 
.A(n_6505),
.Y(n_6841)
);

HB1xp67_ASAP7_75t_L g6842 ( 
.A(n_6308),
.Y(n_6842)
);

OAI21xp5_ASAP7_75t_L g6843 ( 
.A1(n_6472),
.A2(n_124),
.B(n_125),
.Y(n_6843)
);

OA21x2_ASAP7_75t_L g6844 ( 
.A1(n_6486),
.A2(n_125),
.B(n_126),
.Y(n_6844)
);

AOI21xp5_ASAP7_75t_L g6845 ( 
.A1(n_6337),
.A2(n_3198),
.B(n_3156),
.Y(n_6845)
);

AOI21xp5_ASAP7_75t_L g6846 ( 
.A1(n_6540),
.A2(n_3203),
.B(n_3198),
.Y(n_6846)
);

OAI21xp5_ASAP7_75t_L g6847 ( 
.A1(n_6256),
.A2(n_125),
.B(n_126),
.Y(n_6847)
);

AO21x2_ASAP7_75t_L g6848 ( 
.A1(n_6460),
.A2(n_127),
.B(n_128),
.Y(n_6848)
);

INVx3_ASAP7_75t_L g6849 ( 
.A(n_6420),
.Y(n_6849)
);

OA21x2_ASAP7_75t_L g6850 ( 
.A1(n_6289),
.A2(n_6348),
.B(n_6367),
.Y(n_6850)
);

AO21x2_ASAP7_75t_L g6851 ( 
.A1(n_6456),
.A2(n_127),
.B(n_128),
.Y(n_6851)
);

INVx1_ASAP7_75t_L g6852 ( 
.A(n_6249),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6249),
.Y(n_6853)
);

BUFx2_ASAP7_75t_R g6854 ( 
.A(n_6446),
.Y(n_6854)
);

AO21x2_ASAP7_75t_L g6855 ( 
.A1(n_6451),
.A2(n_127),
.B(n_129),
.Y(n_6855)
);

NAND2xp5_ASAP7_75t_L g6856 ( 
.A(n_6535),
.B(n_6312),
.Y(n_6856)
);

OR2x2_ASAP7_75t_L g6857 ( 
.A(n_6412),
.B(n_129),
.Y(n_6857)
);

INVx2_ASAP7_75t_L g6858 ( 
.A(n_6445),
.Y(n_6858)
);

INVx2_ASAP7_75t_SL g6859 ( 
.A(n_6410),
.Y(n_6859)
);

OAI21x1_ASAP7_75t_L g6860 ( 
.A1(n_6481),
.A2(n_130),
.B(n_131),
.Y(n_6860)
);

OAI21x1_ASAP7_75t_L g6861 ( 
.A1(n_6251),
.A2(n_130),
.B(n_131),
.Y(n_6861)
);

OAI21x1_ASAP7_75t_L g6862 ( 
.A1(n_6214),
.A2(n_130),
.B(n_131),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6249),
.Y(n_6863)
);

NOR2xp67_ASAP7_75t_L g6864 ( 
.A(n_6479),
.B(n_132),
.Y(n_6864)
);

INVx2_ASAP7_75t_L g6865 ( 
.A(n_6753),
.Y(n_6865)
);

OAI21x1_ASAP7_75t_L g6866 ( 
.A1(n_6768),
.A2(n_6582),
.B(n_6597),
.Y(n_6866)
);

BUFx2_ASAP7_75t_L g6867 ( 
.A(n_6581),
.Y(n_6867)
);

INVx1_ASAP7_75t_L g6868 ( 
.A(n_6631),
.Y(n_6868)
);

CKINVDCx8_ASAP7_75t_R g6869 ( 
.A(n_6635),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6631),
.Y(n_6870)
);

AO31x2_ASAP7_75t_L g6871 ( 
.A1(n_6579),
.A2(n_6775),
.A3(n_6704),
.B(n_6827),
.Y(n_6871)
);

INVx1_ASAP7_75t_L g6872 ( 
.A(n_6619),
.Y(n_6872)
);

NAND2xp5_ASAP7_75t_L g6873 ( 
.A(n_6772),
.B(n_6458),
.Y(n_6873)
);

CKINVDCx20_ASAP7_75t_R g6874 ( 
.A(n_6588),
.Y(n_6874)
);

INVx2_ASAP7_75t_L g6875 ( 
.A(n_6687),
.Y(n_6875)
);

OAI21x1_ASAP7_75t_L g6876 ( 
.A1(n_6582),
.A2(n_6482),
.B(n_6362),
.Y(n_6876)
);

OAI21x1_ASAP7_75t_L g6877 ( 
.A1(n_6704),
.A2(n_6431),
.B(n_6508),
.Y(n_6877)
);

OAI21x1_ASAP7_75t_L g6878 ( 
.A1(n_6607),
.A2(n_6523),
.B(n_6545),
.Y(n_6878)
);

AO21x2_ASAP7_75t_L g6879 ( 
.A1(n_6775),
.A2(n_6706),
.B(n_6745),
.Y(n_6879)
);

AO21x2_ASAP7_75t_L g6880 ( 
.A1(n_6706),
.A2(n_6374),
.B(n_6370),
.Y(n_6880)
);

AOI21xp5_ASAP7_75t_L g6881 ( 
.A1(n_6681),
.A2(n_6450),
.B(n_6386),
.Y(n_6881)
);

OA21x2_ASAP7_75t_L g6882 ( 
.A1(n_6745),
.A2(n_6285),
.B(n_6203),
.Y(n_6882)
);

AND2x4_ASAP7_75t_L g6883 ( 
.A(n_6625),
.B(n_6484),
.Y(n_6883)
);

AOI22x1_ASAP7_75t_L g6884 ( 
.A1(n_6598),
.A2(n_6693),
.B1(n_6839),
.B2(n_6571),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6797),
.B(n_6484),
.Y(n_6885)
);

OA21x2_ASAP7_75t_L g6886 ( 
.A1(n_6580),
.A2(n_6413),
.B(n_6375),
.Y(n_6886)
);

OAI21x1_ASAP7_75t_L g6887 ( 
.A1(n_6607),
.A2(n_6523),
.B(n_6452),
.Y(n_6887)
);

BUFx2_ASAP7_75t_SL g6888 ( 
.A(n_6648),
.Y(n_6888)
);

HB1xp67_ASAP7_75t_L g6889 ( 
.A(n_6618),
.Y(n_6889)
);

INVx2_ASAP7_75t_L g6890 ( 
.A(n_6603),
.Y(n_6890)
);

AO21x2_ASAP7_75t_L g6891 ( 
.A1(n_6759),
.A2(n_6478),
.B(n_6439),
.Y(n_6891)
);

AO21x2_ASAP7_75t_L g6892 ( 
.A1(n_6759),
.A2(n_6552),
.B(n_6534),
.Y(n_6892)
);

NAND3xp33_ASAP7_75t_L g6893 ( 
.A(n_6734),
.B(n_6685),
.C(n_6671),
.Y(n_6893)
);

AND2x4_ASAP7_75t_L g6894 ( 
.A(n_6625),
.B(n_6797),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_6619),
.Y(n_6895)
);

OAI21x1_ASAP7_75t_L g6896 ( 
.A1(n_6650),
.A2(n_6444),
.B(n_6360),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6575),
.Y(n_6897)
);

INVx2_ASAP7_75t_L g6898 ( 
.A(n_6675),
.Y(n_6898)
);

AOI21x1_ASAP7_75t_L g6899 ( 
.A1(n_6798),
.A2(n_6535),
.B(n_6468),
.Y(n_6899)
);

OAI21x1_ASAP7_75t_L g6900 ( 
.A1(n_6650),
.A2(n_6365),
.B(n_6357),
.Y(n_6900)
);

INVx2_ASAP7_75t_L g6901 ( 
.A(n_6694),
.Y(n_6901)
);

INVx2_ASAP7_75t_L g6902 ( 
.A(n_6602),
.Y(n_6902)
);

AND2x4_ASAP7_75t_L g6903 ( 
.A(n_6723),
.B(n_6727),
.Y(n_6903)
);

INVx1_ASAP7_75t_L g6904 ( 
.A(n_6583),
.Y(n_6904)
);

OAI21xp5_ASAP7_75t_L g6905 ( 
.A1(n_6734),
.A2(n_6435),
.B(n_6390),
.Y(n_6905)
);

OA21x2_ASAP7_75t_L g6906 ( 
.A1(n_6612),
.A2(n_6206),
.B(n_6492),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6602),
.Y(n_6907)
);

HB1xp67_ASAP7_75t_L g6908 ( 
.A(n_6726),
.Y(n_6908)
);

NAND2x1p5_ASAP7_75t_L g6909 ( 
.A(n_6770),
.B(n_6479),
.Y(n_6909)
);

OAI21x1_ASAP7_75t_L g6910 ( 
.A1(n_6612),
.A2(n_6376),
.B(n_6519),
.Y(n_6910)
);

NAND2xp5_ASAP7_75t_L g6911 ( 
.A(n_6772),
.B(n_6493),
.Y(n_6911)
);

AND2x2_ASAP7_75t_L g6912 ( 
.A(n_6657),
.B(n_6308),
.Y(n_6912)
);

AND2x2_ASAP7_75t_L g6913 ( 
.A(n_6678),
.B(n_6308),
.Y(n_6913)
);

OAI21x1_ASAP7_75t_L g6914 ( 
.A1(n_6713),
.A2(n_6300),
.B(n_6402),
.Y(n_6914)
);

OAI21x1_ASAP7_75t_L g6915 ( 
.A1(n_6713),
.A2(n_6623),
.B(n_6849),
.Y(n_6915)
);

OAI21x1_ASAP7_75t_L g6916 ( 
.A1(n_6623),
.A2(n_6403),
.B(n_6550),
.Y(n_6916)
);

NAND2x1p5_ASAP7_75t_L g6917 ( 
.A(n_6770),
.B(n_6536),
.Y(n_6917)
);

AO21x2_ASAP7_75t_L g6918 ( 
.A1(n_6805),
.A2(n_6436),
.B(n_6366),
.Y(n_6918)
);

AND2x4_ASAP7_75t_L g6919 ( 
.A(n_6605),
.B(n_6777),
.Y(n_6919)
);

NAND2xp5_ASAP7_75t_L g6920 ( 
.A(n_6573),
.B(n_6522),
.Y(n_6920)
);

AO21x2_ASAP7_75t_L g6921 ( 
.A1(n_6805),
.A2(n_6568),
.B(n_6820),
.Y(n_6921)
);

OAI21x1_ASAP7_75t_L g6922 ( 
.A1(n_6849),
.A2(n_6273),
.B(n_6516),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6585),
.Y(n_6923)
);

AOI21x1_ASAP7_75t_L g6924 ( 
.A1(n_6798),
.A2(n_6497),
.B(n_6368),
.Y(n_6924)
);

OAI21x1_ASAP7_75t_L g6925 ( 
.A1(n_6599),
.A2(n_6417),
.B(n_6409),
.Y(n_6925)
);

INVxp67_ASAP7_75t_L g6926 ( 
.A(n_6854),
.Y(n_6926)
);

BUFx12f_ASAP7_75t_L g6927 ( 
.A(n_6667),
.Y(n_6927)
);

OAI21xp5_ASAP7_75t_L g6928 ( 
.A1(n_6681),
.A2(n_6466),
.B(n_6464),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_L g6929 ( 
.A(n_6702),
.B(n_6543),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6593),
.Y(n_6930)
);

NAND2x1p5_ASAP7_75t_L g6931 ( 
.A(n_6773),
.B(n_6505),
.Y(n_6931)
);

INVx2_ASAP7_75t_L g6932 ( 
.A(n_6568),
.Y(n_6932)
);

AOI21xp33_ASAP7_75t_SL g6933 ( 
.A1(n_6742),
.A2(n_6404),
.B(n_6514),
.Y(n_6933)
);

OAI21xp5_ASAP7_75t_L g6934 ( 
.A1(n_6821),
.A2(n_6437),
.B(n_6558),
.Y(n_6934)
);

OR2x6_ASAP7_75t_L g6935 ( 
.A(n_6643),
.B(n_6505),
.Y(n_6935)
);

BUFx3_ASAP7_75t_L g6936 ( 
.A(n_6581),
.Y(n_6936)
);

OAI21x1_ASAP7_75t_L g6937 ( 
.A1(n_6630),
.A2(n_6670),
.B(n_6829),
.Y(n_6937)
);

AO21x2_ASAP7_75t_L g6938 ( 
.A1(n_6609),
.A2(n_6495),
.B(n_6443),
.Y(n_6938)
);

OAI21x1_ASAP7_75t_L g6939 ( 
.A1(n_6829),
.A2(n_6555),
.B(n_6461),
.Y(n_6939)
);

OAI21x1_ASAP7_75t_SL g6940 ( 
.A1(n_6703),
.A2(n_6415),
.B(n_6287),
.Y(n_6940)
);

INVxp33_ASAP7_75t_L g6941 ( 
.A(n_6666),
.Y(n_6941)
);

CKINVDCx11_ASAP7_75t_R g6942 ( 
.A(n_6636),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6633),
.Y(n_6943)
);

AO21x2_ASAP7_75t_L g6944 ( 
.A1(n_6692),
.A2(n_6506),
.B(n_6395),
.Y(n_6944)
);

AO21x2_ASAP7_75t_L g6945 ( 
.A1(n_6707),
.A2(n_6393),
.B(n_6498),
.Y(n_6945)
);

OAI21x1_ASAP7_75t_L g6946 ( 
.A1(n_6594),
.A2(n_6544),
.B(n_6524),
.Y(n_6946)
);

AO31x2_ASAP7_75t_L g6947 ( 
.A1(n_6852),
.A2(n_6496),
.A3(n_6547),
.B(n_6287),
.Y(n_6947)
);

AND2x4_ASAP7_75t_L g6948 ( 
.A(n_6605),
.B(n_6363),
.Y(n_6948)
);

INVx1_ASAP7_75t_L g6949 ( 
.A(n_6637),
.Y(n_6949)
);

NAND2xp5_ASAP7_75t_L g6950 ( 
.A(n_6702),
.B(n_6388),
.Y(n_6950)
);

BUFx2_ASAP7_75t_L g6951 ( 
.A(n_6682),
.Y(n_6951)
);

OA21x2_ASAP7_75t_L g6952 ( 
.A1(n_6620),
.A2(n_6332),
.B(n_6244),
.Y(n_6952)
);

AND2x4_ASAP7_75t_L g6953 ( 
.A(n_6778),
.B(n_6363),
.Y(n_6953)
);

NOR2xp33_ASAP7_75t_L g6954 ( 
.A(n_6590),
.B(n_6216),
.Y(n_6954)
);

OAI21xp5_ASAP7_75t_L g6955 ( 
.A1(n_6821),
.A2(n_6560),
.B(n_6371),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6645),
.Y(n_6956)
);

INVx2_ASAP7_75t_L g6957 ( 
.A(n_6726),
.Y(n_6957)
);

INVx1_ASAP7_75t_L g6958 ( 
.A(n_6647),
.Y(n_6958)
);

OR2x6_ASAP7_75t_L g6959 ( 
.A(n_6782),
.B(n_6363),
.Y(n_6959)
);

OAI21x1_ASAP7_75t_L g6960 ( 
.A1(n_6584),
.A2(n_6553),
.B(n_6471),
.Y(n_6960)
);

OAI21x1_ASAP7_75t_L g6961 ( 
.A1(n_6661),
.A2(n_6467),
.B(n_6369),
.Y(n_6961)
);

AOI21x1_ASAP7_75t_L g6962 ( 
.A1(n_6735),
.A2(n_6287),
.B(n_6310),
.Y(n_6962)
);

OAI21x1_ASAP7_75t_L g6963 ( 
.A1(n_6661),
.A2(n_6226),
.B(n_6263),
.Y(n_6963)
);

AOI22xp5_ASAP7_75t_L g6964 ( 
.A1(n_6793),
.A2(n_6548),
.B1(n_6310),
.B2(n_6219),
.Y(n_6964)
);

OAI21x1_ASAP7_75t_L g6965 ( 
.A1(n_6601),
.A2(n_6316),
.B(n_6284),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6649),
.Y(n_6966)
);

OA21x2_ASAP7_75t_L g6967 ( 
.A1(n_6622),
.A2(n_6310),
.B(n_6388),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6665),
.Y(n_6968)
);

BUFx3_ASAP7_75t_L g6969 ( 
.A(n_6613),
.Y(n_6969)
);

AO21x2_ASAP7_75t_L g6970 ( 
.A1(n_6707),
.A2(n_6517),
.B(n_6559),
.Y(n_6970)
);

OA21x2_ASAP7_75t_L g6971 ( 
.A1(n_6641),
.A2(n_6388),
.B(n_6559),
.Y(n_6971)
);

OAI21x1_ASAP7_75t_L g6972 ( 
.A1(n_6574),
.A2(n_6242),
.B(n_6559),
.Y(n_6972)
);

OAI21xp5_ASAP7_75t_L g6973 ( 
.A1(n_6577),
.A2(n_6270),
.B(n_133),
.Y(n_6973)
);

INVx2_ASAP7_75t_L g6974 ( 
.A(n_6639),
.Y(n_6974)
);

OAI21xp5_ASAP7_75t_L g6975 ( 
.A1(n_6577),
.A2(n_6270),
.B(n_133),
.Y(n_6975)
);

OAI21x1_ASAP7_75t_L g6976 ( 
.A1(n_6576),
.A2(n_6242),
.B(n_6270),
.Y(n_6976)
);

NOR2x1_ASAP7_75t_SL g6977 ( 
.A(n_6769),
.B(n_6242),
.Y(n_6977)
);

OAI21x1_ASAP7_75t_L g6978 ( 
.A1(n_6668),
.A2(n_6445),
.B(n_6490),
.Y(n_6978)
);

OAI21x1_ASAP7_75t_L g6979 ( 
.A1(n_6668),
.A2(n_6445),
.B(n_6490),
.Y(n_6979)
);

NOR2xp33_ASAP7_75t_L g6980 ( 
.A(n_6590),
.B(n_390),
.Y(n_6980)
);

OAI21x1_ASAP7_75t_L g6981 ( 
.A1(n_6676),
.A2(n_6490),
.B(n_133),
.Y(n_6981)
);

OA21x2_ASAP7_75t_L g6982 ( 
.A1(n_6698),
.A2(n_134),
.B(n_135),
.Y(n_6982)
);

OAI21x1_ASAP7_75t_L g6983 ( 
.A1(n_6676),
.A2(n_134),
.B(n_135),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6639),
.Y(n_6984)
);

OA21x2_ASAP7_75t_L g6985 ( 
.A1(n_6748),
.A2(n_135),
.B(n_136),
.Y(n_6985)
);

OAI21x1_ASAP7_75t_L g6986 ( 
.A1(n_6596),
.A2(n_136),
.B(n_137),
.Y(n_6986)
);

OA21x2_ASAP7_75t_L g6987 ( 
.A1(n_6763),
.A2(n_136),
.B(n_138),
.Y(n_6987)
);

AO22x2_ASAP7_75t_L g6988 ( 
.A1(n_6806),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_6988)
);

NOR2x1_ASAP7_75t_SL g6989 ( 
.A(n_6792),
.B(n_1677),
.Y(n_6989)
);

INVx1_ASAP7_75t_L g6990 ( 
.A(n_6695),
.Y(n_6990)
);

AND2x2_ASAP7_75t_L g6991 ( 
.A(n_6566),
.B(n_140),
.Y(n_6991)
);

AND2x4_ASAP7_75t_L g6992 ( 
.A(n_6812),
.B(n_141),
.Y(n_6992)
);

OAI21x1_ASAP7_75t_L g6993 ( 
.A1(n_6610),
.A2(n_141),
.B(n_142),
.Y(n_6993)
);

OAI21x1_ASAP7_75t_L g6994 ( 
.A1(n_6614),
.A2(n_141),
.B(n_142),
.Y(n_6994)
);

OAI21x1_ASAP7_75t_L g6995 ( 
.A1(n_6729),
.A2(n_6674),
.B(n_6621),
.Y(n_6995)
);

NOR2xp33_ASAP7_75t_L g6996 ( 
.A(n_6608),
.B(n_390),
.Y(n_6996)
);

OAI21x1_ASAP7_75t_L g6997 ( 
.A1(n_6621),
.A2(n_6863),
.B(n_6853),
.Y(n_6997)
);

OA21x2_ASAP7_75t_L g6998 ( 
.A1(n_6651),
.A2(n_6804),
.B(n_6656),
.Y(n_6998)
);

OAI21x1_ASAP7_75t_L g6999 ( 
.A1(n_6664),
.A2(n_142),
.B(n_143),
.Y(n_6999)
);

BUFx2_ASAP7_75t_L g7000 ( 
.A(n_6688),
.Y(n_7000)
);

OA21x2_ASAP7_75t_L g7001 ( 
.A1(n_6651),
.A2(n_6569),
.B(n_6856),
.Y(n_7001)
);

OAI21xp5_ASAP7_75t_L g7002 ( 
.A1(n_6718),
.A2(n_143),
.B(n_144),
.Y(n_7002)
);

OAI21xp5_ASAP7_75t_L g7003 ( 
.A1(n_6744),
.A2(n_145),
.B(n_146),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6673),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6691),
.Y(n_7005)
);

O2A1O1Ixp33_ASAP7_75t_L g7006 ( 
.A1(n_6839),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_7006)
);

OAI21x1_ASAP7_75t_L g7007 ( 
.A1(n_6664),
.A2(n_145),
.B(n_146),
.Y(n_7007)
);

OAI21x1_ASAP7_75t_L g7008 ( 
.A1(n_6663),
.A2(n_147),
.B(n_148),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6776),
.Y(n_7009)
);

INVx1_ASAP7_75t_L g7010 ( 
.A(n_6776),
.Y(n_7010)
);

NAND3xp33_ASAP7_75t_L g7011 ( 
.A(n_6671),
.B(n_6817),
.C(n_6816),
.Y(n_7011)
);

AO21x1_ASAP7_75t_L g7012 ( 
.A1(n_6856),
.A2(n_148),
.B(n_149),
.Y(n_7012)
);

INVx6_ASAP7_75t_L g7013 ( 
.A(n_6782),
.Y(n_7013)
);

OAI21x1_ASAP7_75t_L g7014 ( 
.A1(n_6586),
.A2(n_6679),
.B(n_6653),
.Y(n_7014)
);

OR2x2_ASAP7_75t_L g7015 ( 
.A(n_6750),
.B(n_148),
.Y(n_7015)
);

NAND2x1p5_ASAP7_75t_L g7016 ( 
.A(n_6773),
.B(n_1677),
.Y(n_7016)
);

BUFx8_ASAP7_75t_L g7017 ( 
.A(n_6578),
.Y(n_7017)
);

INVx1_ASAP7_75t_L g7018 ( 
.A(n_6784),
.Y(n_7018)
);

OAI21x1_ASAP7_75t_SL g7019 ( 
.A1(n_6817),
.A2(n_149),
.B(n_150),
.Y(n_7019)
);

NOR2x1_ASAP7_75t_SL g7020 ( 
.A(n_6747),
.B(n_6669),
.Y(n_7020)
);

INVx1_ASAP7_75t_L g7021 ( 
.A(n_6784),
.Y(n_7021)
);

OAI21x1_ASAP7_75t_SL g7022 ( 
.A1(n_6830),
.A2(n_149),
.B(n_150),
.Y(n_7022)
);

OA21x2_ASAP7_75t_L g7023 ( 
.A1(n_6710),
.A2(n_151),
.B(n_152),
.Y(n_7023)
);

BUFx2_ASAP7_75t_L g7024 ( 
.A(n_6688),
.Y(n_7024)
);

OAI21x1_ASAP7_75t_L g7025 ( 
.A1(n_6644),
.A2(n_151),
.B(n_152),
.Y(n_7025)
);

INVx2_ASAP7_75t_L g7026 ( 
.A(n_6733),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6757),
.Y(n_7027)
);

NOR2xp33_ASAP7_75t_L g7028 ( 
.A(n_6608),
.B(n_391),
.Y(n_7028)
);

INVx3_ASAP7_75t_L g7029 ( 
.A(n_6751),
.Y(n_7029)
);

OAI21x1_ASAP7_75t_L g7030 ( 
.A1(n_6644),
.A2(n_6653),
.B(n_6616),
.Y(n_7030)
);

NAND2x1p5_ASAP7_75t_L g7031 ( 
.A(n_6864),
.B(n_1678),
.Y(n_7031)
);

BUFx6f_ASAP7_75t_L g7032 ( 
.A(n_6758),
.Y(n_7032)
);

OAI21x1_ASAP7_75t_L g7033 ( 
.A1(n_6749),
.A2(n_151),
.B(n_152),
.Y(n_7033)
);

OR2x6_ASAP7_75t_L g7034 ( 
.A(n_6736),
.B(n_1678),
.Y(n_7034)
);

AND2x4_ASAP7_75t_L g7035 ( 
.A(n_6716),
.B(n_153),
.Y(n_7035)
);

INVx3_ASAP7_75t_L g7036 ( 
.A(n_6628),
.Y(n_7036)
);

OAI21x1_ASAP7_75t_SL g7037 ( 
.A1(n_6859),
.A2(n_153),
.B(n_154),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6757),
.Y(n_7038)
);

INVxp67_ASAP7_75t_L g7039 ( 
.A(n_6854),
.Y(n_7039)
);

OAI21x1_ASAP7_75t_L g7040 ( 
.A1(n_6646),
.A2(n_154),
.B(n_155),
.Y(n_7040)
);

OA21x2_ASAP7_75t_L g7041 ( 
.A1(n_6737),
.A2(n_155),
.B(n_156),
.Y(n_7041)
);

NAND2xp5_ASAP7_75t_L g7042 ( 
.A(n_6816),
.B(n_391),
.Y(n_7042)
);

BUFx3_ASAP7_75t_L g7043 ( 
.A(n_6652),
.Y(n_7043)
);

OAI21x1_ASAP7_75t_L g7044 ( 
.A1(n_6760),
.A2(n_157),
.B(n_158),
.Y(n_7044)
);

OA21x2_ASAP7_75t_L g7045 ( 
.A1(n_6738),
.A2(n_157),
.B(n_158),
.Y(n_7045)
);

CKINVDCx20_ASAP7_75t_R g7046 ( 
.A(n_6709),
.Y(n_7046)
);

AO21x2_ASAP7_75t_L g7047 ( 
.A1(n_6864),
.A2(n_6855),
.B(n_6787),
.Y(n_7047)
);

INVx2_ASAP7_75t_L g7048 ( 
.A(n_6740),
.Y(n_7048)
);

NOR2xp67_ASAP7_75t_L g7049 ( 
.A(n_6842),
.B(n_158),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_6810),
.Y(n_7050)
);

NAND2xp5_ASAP7_75t_L g7051 ( 
.A(n_6844),
.B(n_392),
.Y(n_7051)
);

OR2x2_ASAP7_75t_L g7052 ( 
.A(n_6764),
.B(n_159),
.Y(n_7052)
);

INVx1_ASAP7_75t_L g7053 ( 
.A(n_6824),
.Y(n_7053)
);

OAI21x1_ASAP7_75t_L g7054 ( 
.A1(n_6761),
.A2(n_160),
.B(n_161),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_6844),
.Y(n_7055)
);

AOI22xp33_ASAP7_75t_L g7056 ( 
.A1(n_6722),
.A2(n_2690),
.B1(n_1751),
.B2(n_1766),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6724),
.Y(n_7057)
);

BUFx3_ASAP7_75t_L g7058 ( 
.A(n_6655),
.Y(n_7058)
);

OR2x2_ASAP7_75t_L g7059 ( 
.A(n_6766),
.B(n_160),
.Y(n_7059)
);

OAI21x1_ASAP7_75t_L g7060 ( 
.A1(n_6799),
.A2(n_161),
.B(n_162),
.Y(n_7060)
);

NOR2xp67_ASAP7_75t_L g7061 ( 
.A(n_6842),
.B(n_161),
.Y(n_7061)
);

BUFx2_ASAP7_75t_L g7062 ( 
.A(n_6789),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_L g7063 ( 
.A(n_6791),
.B(n_392),
.Y(n_7063)
);

CKINVDCx14_ASAP7_75t_R g7064 ( 
.A(n_6683),
.Y(n_7064)
);

INVx2_ASAP7_75t_SL g7065 ( 
.A(n_6589),
.Y(n_7065)
);

INVx3_ASAP7_75t_L g7066 ( 
.A(n_6628),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6724),
.Y(n_7067)
);

OAI21x1_ASAP7_75t_L g7068 ( 
.A1(n_6624),
.A2(n_162),
.B(n_163),
.Y(n_7068)
);

INVxp67_ASAP7_75t_L g7069 ( 
.A(n_6848),
.Y(n_7069)
);

OA21x2_ASAP7_75t_L g7070 ( 
.A1(n_6783),
.A2(n_6795),
.B(n_6794),
.Y(n_7070)
);

INVx3_ASAP7_75t_L g7071 ( 
.A(n_6736),
.Y(n_7071)
);

CKINVDCx16_ASAP7_75t_R g7072 ( 
.A(n_6658),
.Y(n_7072)
);

INVx2_ASAP7_75t_L g7073 ( 
.A(n_6659),
.Y(n_7073)
);

BUFx2_ASAP7_75t_R g7074 ( 
.A(n_6732),
.Y(n_7074)
);

NAND2xp5_ASAP7_75t_L g7075 ( 
.A(n_6791),
.B(n_393),
.Y(n_7075)
);

NOR2xp33_ASAP7_75t_L g7076 ( 
.A(n_6598),
.B(n_394),
.Y(n_7076)
);

AND2x2_ASAP7_75t_L g7077 ( 
.A(n_6626),
.B(n_163),
.Y(n_7077)
);

OA21x2_ASAP7_75t_L g7078 ( 
.A1(n_6809),
.A2(n_164),
.B(n_165),
.Y(n_7078)
);

AOI22xp33_ASAP7_75t_L g7079 ( 
.A1(n_6722),
.A2(n_1751),
.B1(n_1766),
.B2(n_1678),
.Y(n_7079)
);

AOI22x1_ASAP7_75t_L g7080 ( 
.A1(n_6708),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_7080)
);

NAND2x1p5_ASAP7_75t_L g7081 ( 
.A(n_6700),
.B(n_1678),
.Y(n_7081)
);

OAI21x1_ASAP7_75t_L g7082 ( 
.A1(n_6640),
.A2(n_165),
.B(n_168),
.Y(n_7082)
);

OAI22xp5_ASAP7_75t_L g7083 ( 
.A1(n_6572),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_7083)
);

INVx2_ASAP7_75t_L g7084 ( 
.A(n_6659),
.Y(n_7084)
);

NAND2xp5_ASAP7_75t_L g7085 ( 
.A(n_6741),
.B(n_395),
.Y(n_7085)
);

INVx3_ASAP7_75t_L g7086 ( 
.A(n_6736),
.Y(n_7086)
);

OAI21x1_ASAP7_75t_L g7087 ( 
.A1(n_6615),
.A2(n_169),
.B(n_170),
.Y(n_7087)
);

CKINVDCx5p33_ASAP7_75t_R g7088 ( 
.A(n_6589),
.Y(n_7088)
);

OAI21x1_ASAP7_75t_L g7089 ( 
.A1(n_6632),
.A2(n_171),
.B(n_172),
.Y(n_7089)
);

INVx2_ASAP7_75t_L g7090 ( 
.A(n_6662),
.Y(n_7090)
);

OAI21x1_ASAP7_75t_L g7091 ( 
.A1(n_6606),
.A2(n_171),
.B(n_173),
.Y(n_7091)
);

INVx2_ASAP7_75t_L g7092 ( 
.A(n_6662),
.Y(n_7092)
);

INVx6_ASAP7_75t_L g7093 ( 
.A(n_6700),
.Y(n_7093)
);

INVx2_ASAP7_75t_L g7094 ( 
.A(n_6806),
.Y(n_7094)
);

OAI21x1_ASAP7_75t_L g7095 ( 
.A1(n_6606),
.A2(n_173),
.B(n_174),
.Y(n_7095)
);

OAI21x1_ASAP7_75t_L g7096 ( 
.A1(n_6721),
.A2(n_173),
.B(n_174),
.Y(n_7096)
);

OAI21xp5_ASAP7_75t_L g7097 ( 
.A1(n_6785),
.A2(n_175),
.B(n_176),
.Y(n_7097)
);

OAI21xp5_ASAP7_75t_L g7098 ( 
.A1(n_6834),
.A2(n_175),
.B(n_176),
.Y(n_7098)
);

AO31x2_ASAP7_75t_L g7099 ( 
.A1(n_6793),
.A2(n_177),
.A3(n_175),
.B(n_176),
.Y(n_7099)
);

NAND2xp5_ASAP7_75t_L g7100 ( 
.A(n_6741),
.B(n_395),
.Y(n_7100)
);

AO21x2_ASAP7_75t_L g7101 ( 
.A1(n_6855),
.A2(n_6787),
.B(n_6848),
.Y(n_7101)
);

CKINVDCx11_ASAP7_75t_R g7102 ( 
.A(n_6813),
.Y(n_7102)
);

OAI21x1_ASAP7_75t_L g7103 ( 
.A1(n_6721),
.A2(n_177),
.B(n_178),
.Y(n_7103)
);

OAI21x1_ASAP7_75t_L g7104 ( 
.A1(n_6697),
.A2(n_177),
.B(n_178),
.Y(n_7104)
);

OA21x2_ASAP7_75t_L g7105 ( 
.A1(n_6811),
.A2(n_178),
.B(n_179),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6851),
.Y(n_7106)
);

NOR2xp33_ASAP7_75t_L g7107 ( 
.A(n_6814),
.B(n_396),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6851),
.Y(n_7108)
);

OA21x2_ASAP7_75t_L g7109 ( 
.A1(n_6815),
.A2(n_6819),
.B(n_6818),
.Y(n_7109)
);

OAI21xp5_ASAP7_75t_L g7110 ( 
.A1(n_6838),
.A2(n_179),
.B(n_180),
.Y(n_7110)
);

NAND2xp5_ASAP7_75t_L g7111 ( 
.A(n_6627),
.B(n_396),
.Y(n_7111)
);

OAI21x1_ASAP7_75t_L g7112 ( 
.A1(n_6697),
.A2(n_180),
.B(n_181),
.Y(n_7112)
);

AND2x4_ASAP7_75t_L g7113 ( 
.A(n_6747),
.B(n_181),
.Y(n_7113)
);

NOR2xp33_ASAP7_75t_L g7114 ( 
.A(n_6754),
.B(n_397),
.Y(n_7114)
);

OA21x2_ASAP7_75t_L g7115 ( 
.A1(n_6826),
.A2(n_182),
.B(n_183),
.Y(n_7115)
);

INVx1_ASAP7_75t_L g7116 ( 
.A(n_6627),
.Y(n_7116)
);

OAI21x1_ASAP7_75t_L g7117 ( 
.A1(n_6699),
.A2(n_182),
.B(n_183),
.Y(n_7117)
);

INVx1_ASAP7_75t_SL g7118 ( 
.A(n_6831),
.Y(n_7118)
);

HB1xp67_ASAP7_75t_L g7119 ( 
.A(n_6836),
.Y(n_7119)
);

NAND2x1p5_ASAP7_75t_L g7120 ( 
.A(n_6803),
.B(n_6832),
.Y(n_7120)
);

OAI21x1_ASAP7_75t_L g7121 ( 
.A1(n_6699),
.A2(n_182),
.B(n_183),
.Y(n_7121)
);

OA21x2_ASAP7_75t_L g7122 ( 
.A1(n_6833),
.A2(n_185),
.B(n_187),
.Y(n_7122)
);

INVx4_ASAP7_75t_SL g7123 ( 
.A(n_6730),
.Y(n_7123)
);

NOR2x1_ASAP7_75t_SL g7124 ( 
.A(n_6747),
.B(n_1751),
.Y(n_7124)
);

INVx2_ASAP7_75t_L g7125 ( 
.A(n_6774),
.Y(n_7125)
);

OAI21x1_ASAP7_75t_L g7126 ( 
.A1(n_6701),
.A2(n_6728),
.B(n_6846),
.Y(n_7126)
);

INVx1_ASAP7_75t_L g7127 ( 
.A(n_6634),
.Y(n_7127)
);

INVx6_ASAP7_75t_L g7128 ( 
.A(n_6803),
.Y(n_7128)
);

AO31x2_ASAP7_75t_L g7129 ( 
.A1(n_6858),
.A2(n_188),
.A3(n_185),
.B(n_187),
.Y(n_7129)
);

OR2x2_ASAP7_75t_L g7130 ( 
.A(n_7005),
.B(n_6857),
.Y(n_7130)
);

OAI22xp5_ASAP7_75t_L g7131 ( 
.A1(n_6893),
.A2(n_6572),
.B1(n_6669),
.B2(n_6828),
.Y(n_7131)
);

BUFx12f_ASAP7_75t_L g7132 ( 
.A(n_6942),
.Y(n_7132)
);

OA21x2_ASAP7_75t_L g7133 ( 
.A1(n_6902),
.A2(n_6567),
.B(n_6611),
.Y(n_7133)
);

INVx1_ASAP7_75t_L g7134 ( 
.A(n_6897),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_6897),
.Y(n_7135)
);

INVx2_ASAP7_75t_L g7136 ( 
.A(n_7047),
.Y(n_7136)
);

NAND2xp5_ASAP7_75t_L g7137 ( 
.A(n_7111),
.B(n_6771),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6904),
.Y(n_7138)
);

AND2x2_ASAP7_75t_L g7139 ( 
.A(n_6867),
.B(n_6841),
.Y(n_7139)
);

NAND2xp5_ASAP7_75t_L g7140 ( 
.A(n_6908),
.B(n_6823),
.Y(n_7140)
);

AOI21xp5_ASAP7_75t_L g7141 ( 
.A1(n_6881),
.A2(n_6611),
.B(n_6802),
.Y(n_7141)
);

OAI22xp5_ASAP7_75t_L g7142 ( 
.A1(n_7072),
.A2(n_6595),
.B1(n_6717),
.B2(n_6843),
.Y(n_7142)
);

AND2x2_ASAP7_75t_L g7143 ( 
.A(n_6903),
.B(n_6765),
.Y(n_7143)
);

AND2x2_ASAP7_75t_L g7144 ( 
.A(n_6903),
.B(n_6885),
.Y(n_7144)
);

HB1xp67_ASAP7_75t_L g7145 ( 
.A(n_6889),
.Y(n_7145)
);

AOI21xp5_ASAP7_75t_L g7146 ( 
.A1(n_7011),
.A2(n_6802),
.B(n_6843),
.Y(n_7146)
);

BUFx2_ASAP7_75t_SL g7147 ( 
.A(n_7046),
.Y(n_7147)
);

NAND2xp5_ASAP7_75t_L g7148 ( 
.A(n_7119),
.B(n_6743),
.Y(n_7148)
);

OA21x2_ASAP7_75t_L g7149 ( 
.A1(n_6907),
.A2(n_6677),
.B(n_6592),
.Y(n_7149)
);

AOI221x1_ASAP7_75t_SL g7150 ( 
.A1(n_7083),
.A2(n_6832),
.B1(n_6696),
.B2(n_6715),
.C(n_190),
.Y(n_7150)
);

INVx2_ASAP7_75t_L g7151 ( 
.A(n_7047),
.Y(n_7151)
);

AOI221xp5_ASAP7_75t_L g7152 ( 
.A1(n_7072),
.A2(n_7069),
.B1(n_6928),
.B2(n_7055),
.C(n_6988),
.Y(n_7152)
);

AND2x2_ASAP7_75t_L g7153 ( 
.A(n_7071),
.B(n_6765),
.Y(n_7153)
);

NAND2xp5_ASAP7_75t_L g7154 ( 
.A(n_6957),
.B(n_6871),
.Y(n_7154)
);

AOI21x1_ASAP7_75t_SL g7155 ( 
.A1(n_6929),
.A2(n_6696),
.B(n_6837),
.Y(n_7155)
);

OAI22xp5_ASAP7_75t_L g7156 ( 
.A1(n_6964),
.A2(n_6669),
.B1(n_6802),
.B2(n_6822),
.Y(n_7156)
);

INVx2_ASAP7_75t_L g7157 ( 
.A(n_6997),
.Y(n_7157)
);

AND2x2_ASAP7_75t_L g7158 ( 
.A(n_7071),
.B(n_6680),
.Y(n_7158)
);

AND2x2_ASAP7_75t_L g7159 ( 
.A(n_7086),
.B(n_6680),
.Y(n_7159)
);

O2A1O1Ixp5_ASAP7_75t_L g7160 ( 
.A1(n_7012),
.A2(n_6865),
.B(n_6962),
.C(n_6950),
.Y(n_7160)
);

BUFx12f_ASAP7_75t_L g7161 ( 
.A(n_6927),
.Y(n_7161)
);

AOI21xp5_ASAP7_75t_L g7162 ( 
.A1(n_7085),
.A2(n_6847),
.B(n_6595),
.Y(n_7162)
);

BUFx2_ASAP7_75t_L g7163 ( 
.A(n_6935),
.Y(n_7163)
);

OAI22xp5_ASAP7_75t_L g7164 ( 
.A1(n_6926),
.A2(n_6822),
.B1(n_6680),
.B2(n_6684),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_L g7165 ( 
.A(n_6871),
.B(n_6634),
.Y(n_7165)
);

O2A1O1Ixp33_ASAP7_75t_L g7166 ( 
.A1(n_6933),
.A2(n_6847),
.B(n_6825),
.C(n_6845),
.Y(n_7166)
);

OA21x2_ASAP7_75t_L g7167 ( 
.A1(n_6866),
.A2(n_6835),
.B(n_6796),
.Y(n_7167)
);

OR2x2_ASAP7_75t_L g7168 ( 
.A(n_7005),
.B(n_6600),
.Y(n_7168)
);

HB1xp67_ASAP7_75t_L g7169 ( 
.A(n_6982),
.Y(n_7169)
);

AND2x2_ASAP7_75t_L g7170 ( 
.A(n_7086),
.B(n_6684),
.Y(n_7170)
);

OA21x2_ASAP7_75t_L g7171 ( 
.A1(n_6915),
.A2(n_6932),
.B(n_7116),
.Y(n_7171)
);

NAND2xp5_ASAP7_75t_L g7172 ( 
.A(n_6871),
.B(n_7050),
.Y(n_7172)
);

OR2x2_ASAP7_75t_L g7173 ( 
.A(n_6901),
.B(n_6600),
.Y(n_7173)
);

NAND2xp5_ASAP7_75t_L g7174 ( 
.A(n_7050),
.B(n_6780),
.Y(n_7174)
);

AND2x2_ASAP7_75t_L g7175 ( 
.A(n_6919),
.B(n_6684),
.Y(n_7175)
);

INVx3_ASAP7_75t_L g7176 ( 
.A(n_7013),
.Y(n_7176)
);

OAI22xp5_ASAP7_75t_L g7177 ( 
.A1(n_7039),
.A2(n_6822),
.B1(n_6701),
.B2(n_6728),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6904),
.Y(n_7178)
);

AOI21xp5_ASAP7_75t_L g7179 ( 
.A1(n_7100),
.A2(n_6825),
.B(n_6755),
.Y(n_7179)
);

AND2x2_ASAP7_75t_L g7180 ( 
.A(n_6919),
.B(n_6600),
.Y(n_7180)
);

AOI21xp5_ASAP7_75t_L g7181 ( 
.A1(n_7042),
.A2(n_6845),
.B(n_6755),
.Y(n_7181)
);

AND2x2_ASAP7_75t_L g7182 ( 
.A(n_6935),
.B(n_6711),
.Y(n_7182)
);

AOI21xp5_ASAP7_75t_SL g7183 ( 
.A1(n_6982),
.A2(n_6807),
.B(n_6654),
.Y(n_7183)
);

OA21x2_ASAP7_75t_L g7184 ( 
.A1(n_7116),
.A2(n_6790),
.B(n_6846),
.Y(n_7184)
);

INVx1_ASAP7_75t_L g7185 ( 
.A(n_6923),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_6923),
.Y(n_7186)
);

OR2x2_ASAP7_75t_L g7187 ( 
.A(n_7094),
.B(n_6780),
.Y(n_7187)
);

A2O1A1Ixp33_ASAP7_75t_L g7188 ( 
.A1(n_7006),
.A2(n_6731),
.B(n_6840),
.C(n_6860),
.Y(n_7188)
);

NAND2xp5_ASAP7_75t_L g7189 ( 
.A(n_7053),
.B(n_6780),
.Y(n_7189)
);

AOI21xp5_ASAP7_75t_L g7190 ( 
.A1(n_7051),
.A2(n_6604),
.B(n_6654),
.Y(n_7190)
);

AOI21xp5_ASAP7_75t_L g7191 ( 
.A1(n_7063),
.A2(n_6604),
.B(n_6807),
.Y(n_7191)
);

NOR2xp67_ASAP7_75t_L g7192 ( 
.A(n_7036),
.B(n_6801),
.Y(n_7192)
);

INVx3_ASAP7_75t_L g7193 ( 
.A(n_7013),
.Y(n_7193)
);

INVx2_ASAP7_75t_SL g7194 ( 
.A(n_7017),
.Y(n_7194)
);

BUFx3_ASAP7_75t_L g7195 ( 
.A(n_6874),
.Y(n_7195)
);

NOR2x1_ASAP7_75t_SL g7196 ( 
.A(n_6959),
.B(n_6591),
.Y(n_7196)
);

A2O1A1Ixp33_ASAP7_75t_L g7197 ( 
.A1(n_6905),
.A2(n_6862),
.B(n_6861),
.C(n_6808),
.Y(n_7197)
);

NOR2xp33_ASAP7_75t_L g7198 ( 
.A(n_7074),
.B(n_6629),
.Y(n_7198)
);

OA21x2_ASAP7_75t_L g7199 ( 
.A1(n_6995),
.A2(n_6720),
.B(n_6725),
.Y(n_7199)
);

INVx3_ASAP7_75t_L g7200 ( 
.A(n_6936),
.Y(n_7200)
);

NOR2xp67_ASAP7_75t_L g7201 ( 
.A(n_7036),
.B(n_6714),
.Y(n_7201)
);

AND2x2_ASAP7_75t_L g7202 ( 
.A(n_6912),
.B(n_6712),
.Y(n_7202)
);

A2O1A1Ixp33_ASAP7_75t_L g7203 ( 
.A1(n_7055),
.A2(n_6800),
.B(n_6752),
.C(n_6730),
.Y(n_7203)
);

AND2x2_ASAP7_75t_L g7204 ( 
.A(n_6894),
.B(n_6570),
.Y(n_7204)
);

NAND2xp5_ASAP7_75t_L g7205 ( 
.A(n_7053),
.B(n_6629),
.Y(n_7205)
);

OAI22xp5_ASAP7_75t_SL g7206 ( 
.A1(n_7064),
.A2(n_6850),
.B1(n_6570),
.B2(n_6730),
.Y(n_7206)
);

NAND2xp5_ASAP7_75t_L g7207 ( 
.A(n_6873),
.B(n_6752),
.Y(n_7207)
);

OAI211xp5_ASAP7_75t_SL g7208 ( 
.A1(n_7002),
.A2(n_6714),
.B(n_190),
.C(n_188),
.Y(n_7208)
);

BUFx2_ASAP7_75t_L g7209 ( 
.A(n_7029),
.Y(n_7209)
);

AOI221xp5_ASAP7_75t_L g7210 ( 
.A1(n_6988),
.A2(n_6591),
.B1(n_6638),
.B2(n_6752),
.C(n_6686),
.Y(n_7210)
);

INVx2_ASAP7_75t_L g7211 ( 
.A(n_6985),
.Y(n_7211)
);

HB1xp67_ASAP7_75t_L g7212 ( 
.A(n_7001),
.Y(n_7212)
);

INVx2_ASAP7_75t_L g7213 ( 
.A(n_6985),
.Y(n_7213)
);

O2A1O1Ixp33_ASAP7_75t_L g7214 ( 
.A1(n_6934),
.A2(n_6638),
.B(n_6850),
.C(n_6686),
.Y(n_7214)
);

AOI21xp5_ASAP7_75t_L g7215 ( 
.A1(n_7075),
.A2(n_6672),
.B(n_6587),
.Y(n_7215)
);

HB1xp67_ASAP7_75t_L g7216 ( 
.A(n_7001),
.Y(n_7216)
);

INVx2_ASAP7_75t_L g7217 ( 
.A(n_6987),
.Y(n_7217)
);

OAI22xp5_ASAP7_75t_L g7218 ( 
.A1(n_6884),
.A2(n_6941),
.B1(n_7029),
.B2(n_7118),
.Y(n_7218)
);

OR2x2_ASAP7_75t_L g7219 ( 
.A(n_6947),
.B(n_6587),
.Y(n_7219)
);

AND2x2_ASAP7_75t_L g7220 ( 
.A(n_6894),
.B(n_6781),
.Y(n_7220)
);

INVx2_ASAP7_75t_L g7221 ( 
.A(n_6987),
.Y(n_7221)
);

OAI22xp5_ASAP7_75t_L g7222 ( 
.A1(n_6884),
.A2(n_6672),
.B1(n_6642),
.B2(n_6617),
.Y(n_7222)
);

CKINVDCx20_ASAP7_75t_R g7223 ( 
.A(n_7102),
.Y(n_7223)
);

INVx2_ASAP7_75t_L g7224 ( 
.A(n_7023),
.Y(n_7224)
);

NAND2xp5_ASAP7_75t_L g7225 ( 
.A(n_6880),
.B(n_6788),
.Y(n_7225)
);

AND2x2_ASAP7_75t_L g7226 ( 
.A(n_7000),
.B(n_6786),
.Y(n_7226)
);

OAI22xp5_ASAP7_75t_L g7227 ( 
.A1(n_7093),
.A2(n_6642),
.B1(n_6617),
.B2(n_6660),
.Y(n_7227)
);

INVx2_ASAP7_75t_L g7228 ( 
.A(n_7023),
.Y(n_7228)
);

O2A1O1Ixp33_ASAP7_75t_L g7229 ( 
.A1(n_7057),
.A2(n_6705),
.B(n_190),
.C(n_191),
.Y(n_7229)
);

INVxp67_ASAP7_75t_L g7230 ( 
.A(n_6888),
.Y(n_7230)
);

AOI21xp5_ASAP7_75t_L g7231 ( 
.A1(n_6880),
.A2(n_6705),
.B(n_6660),
.Y(n_7231)
);

AND2x2_ASAP7_75t_L g7232 ( 
.A(n_7024),
.B(n_6746),
.Y(n_7232)
);

AND2x4_ASAP7_75t_L g7233 ( 
.A(n_6959),
.B(n_6762),
.Y(n_7233)
);

AND2x2_ASAP7_75t_L g7234 ( 
.A(n_6883),
.B(n_6756),
.Y(n_7234)
);

AOI21xp5_ASAP7_75t_SL g7235 ( 
.A1(n_6989),
.A2(n_6689),
.B(n_188),
.Y(n_7235)
);

OAI22xp5_ASAP7_75t_L g7236 ( 
.A1(n_7093),
.A2(n_6689),
.B1(n_6779),
.B2(n_6767),
.Y(n_7236)
);

AND2x2_ASAP7_75t_L g7237 ( 
.A(n_6883),
.B(n_6739),
.Y(n_7237)
);

O2A1O1Ixp33_ASAP7_75t_L g7238 ( 
.A1(n_7057),
.A2(n_192),
.B(n_193),
.C(n_191),
.Y(n_7238)
);

AOI22xp5_ASAP7_75t_L g7239 ( 
.A1(n_6891),
.A2(n_6690),
.B1(n_6719),
.B2(n_2959),
.Y(n_7239)
);

AND2x2_ASAP7_75t_L g7240 ( 
.A(n_7066),
.B(n_189),
.Y(n_7240)
);

NAND2xp5_ASAP7_75t_L g7241 ( 
.A(n_7067),
.B(n_398),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_6930),
.Y(n_7242)
);

AND2x2_ASAP7_75t_L g7243 ( 
.A(n_7066),
.B(n_192),
.Y(n_7243)
);

BUFx3_ASAP7_75t_L g7244 ( 
.A(n_7017),
.Y(n_7244)
);

CKINVDCx20_ASAP7_75t_R g7245 ( 
.A(n_6869),
.Y(n_7245)
);

AND2x2_ASAP7_75t_L g7246 ( 
.A(n_6913),
.B(n_192),
.Y(n_7246)
);

AOI21xp5_ASAP7_75t_L g7247 ( 
.A1(n_7067),
.A2(n_193),
.B(n_194),
.Y(n_7247)
);

O2A1O1Ixp33_ASAP7_75t_L g7248 ( 
.A1(n_7003),
.A2(n_195),
.B(n_197),
.C(n_194),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_6930),
.Y(n_7249)
);

OAI22xp5_ASAP7_75t_L g7250 ( 
.A1(n_7120),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_L g7251 ( 
.A(n_6879),
.B(n_399),
.Y(n_7251)
);

O2A1O1Ixp33_ASAP7_75t_L g7252 ( 
.A1(n_7097),
.A2(n_200),
.B(n_201),
.C(n_199),
.Y(n_7252)
);

NAND2xp5_ASAP7_75t_L g7253 ( 
.A(n_6879),
.B(n_401),
.Y(n_7253)
);

OAI22xp5_ASAP7_75t_L g7254 ( 
.A1(n_7128),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_7254)
);

A2O1A1Ixp33_ASAP7_75t_L g7255 ( 
.A1(n_7098),
.A2(n_202),
.B(n_198),
.C(n_201),
.Y(n_7255)
);

OA21x2_ASAP7_75t_L g7256 ( 
.A1(n_7127),
.A2(n_198),
.B(n_202),
.Y(n_7256)
);

AND2x2_ASAP7_75t_L g7257 ( 
.A(n_6953),
.B(n_202),
.Y(n_7257)
);

AND2x2_ASAP7_75t_L g7258 ( 
.A(n_6953),
.B(n_203),
.Y(n_7258)
);

AND2x4_ASAP7_75t_L g7259 ( 
.A(n_7065),
.B(n_203),
.Y(n_7259)
);

CKINVDCx20_ASAP7_75t_R g7260 ( 
.A(n_7043),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_6943),
.Y(n_7261)
);

OAI22xp5_ASAP7_75t_L g7262 ( 
.A1(n_7128),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_6943),
.Y(n_7263)
);

BUFx6f_ASAP7_75t_L g7264 ( 
.A(n_7058),
.Y(n_7264)
);

CKINVDCx5p33_ASAP7_75t_R g7265 ( 
.A(n_7088),
.Y(n_7265)
);

AOI21x1_ASAP7_75t_SL g7266 ( 
.A1(n_7035),
.A2(n_204),
.B(n_205),
.Y(n_7266)
);

INVxp67_ASAP7_75t_L g7267 ( 
.A(n_6996),
.Y(n_7267)
);

AND2x4_ASAP7_75t_L g7268 ( 
.A(n_7113),
.B(n_204),
.Y(n_7268)
);

O2A1O1Ixp5_ASAP7_75t_L g7269 ( 
.A1(n_7110),
.A2(n_207),
.B(n_205),
.C(n_206),
.Y(n_7269)
);

AND2x2_ASAP7_75t_L g7270 ( 
.A(n_6909),
.B(n_206),
.Y(n_7270)
);

AOI21xp5_ASAP7_75t_SL g7271 ( 
.A1(n_6989),
.A2(n_206),
.B(n_207),
.Y(n_7271)
);

O2A1O1Ixp5_ASAP7_75t_L g7272 ( 
.A1(n_6872),
.A2(n_210),
.B(n_207),
.C(n_209),
.Y(n_7272)
);

BUFx3_ASAP7_75t_L g7273 ( 
.A(n_7062),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_L g7274 ( 
.A(n_7101),
.B(n_401),
.Y(n_7274)
);

OA21x2_ASAP7_75t_L g7275 ( 
.A1(n_7127),
.A2(n_209),
.B(n_211),
.Y(n_7275)
);

OAI22xp5_ASAP7_75t_L g7276 ( 
.A1(n_6973),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_7276)
);

BUFx3_ASAP7_75t_L g7277 ( 
.A(n_6951),
.Y(n_7277)
);

HB1xp67_ASAP7_75t_L g7278 ( 
.A(n_6949),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_6949),
.Y(n_7279)
);

INVx1_ASAP7_75t_L g7280 ( 
.A(n_6956),
.Y(n_7280)
);

NAND2xp5_ASAP7_75t_L g7281 ( 
.A(n_7101),
.B(n_6918),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_6956),
.Y(n_7282)
);

O2A1O1Ixp5_ASAP7_75t_L g7283 ( 
.A1(n_6872),
.A2(n_213),
.B(n_211),
.C(n_212),
.Y(n_7283)
);

OR2x2_ASAP7_75t_L g7284 ( 
.A(n_6947),
.B(n_213),
.Y(n_7284)
);

CKINVDCx12_ASAP7_75t_R g7285 ( 
.A(n_7077),
.Y(n_7285)
);

OAI22xp5_ASAP7_75t_L g7286 ( 
.A1(n_6975),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_7286)
);

NAND2xp5_ASAP7_75t_L g7287 ( 
.A(n_6918),
.B(n_402),
.Y(n_7287)
);

INVx1_ASAP7_75t_SL g7288 ( 
.A(n_7035),
.Y(n_7288)
);

AND2x2_ASAP7_75t_L g7289 ( 
.A(n_7125),
.B(n_214),
.Y(n_7289)
);

AOI21xp5_ASAP7_75t_L g7290 ( 
.A1(n_6940),
.A2(n_214),
.B(n_215),
.Y(n_7290)
);

NAND2xp5_ASAP7_75t_L g7291 ( 
.A(n_6991),
.B(n_403),
.Y(n_7291)
);

AND2x2_ASAP7_75t_L g7292 ( 
.A(n_6948),
.B(n_215),
.Y(n_7292)
);

BUFx12f_ASAP7_75t_L g7293 ( 
.A(n_6969),
.Y(n_7293)
);

OA21x2_ASAP7_75t_L g7294 ( 
.A1(n_6937),
.A2(n_216),
.B(n_217),
.Y(n_7294)
);

NOR2xp67_ASAP7_75t_L g7295 ( 
.A(n_6868),
.B(n_6870),
.Y(n_7295)
);

AOI21xp5_ASAP7_75t_L g7296 ( 
.A1(n_6944),
.A2(n_217),
.B(n_218),
.Y(n_7296)
);

AOI21x1_ASAP7_75t_SL g7297 ( 
.A1(n_6948),
.A2(n_218),
.B(n_219),
.Y(n_7297)
);

O2A1O1Ixp33_ASAP7_75t_L g7298 ( 
.A1(n_7106),
.A2(n_221),
.B(n_222),
.C(n_220),
.Y(n_7298)
);

AOI21x1_ASAP7_75t_SL g7299 ( 
.A1(n_6992),
.A2(n_6911),
.B(n_7113),
.Y(n_7299)
);

AOI21xp5_ASAP7_75t_L g7300 ( 
.A1(n_6944),
.A2(n_218),
.B(n_220),
.Y(n_7300)
);

INVx2_ASAP7_75t_L g7301 ( 
.A(n_7041),
.Y(n_7301)
);

OR2x2_ASAP7_75t_L g7302 ( 
.A(n_6947),
.B(n_221),
.Y(n_7302)
);

AND2x2_ASAP7_75t_L g7303 ( 
.A(n_6931),
.B(n_221),
.Y(n_7303)
);

AND2x4_ASAP7_75t_L g7304 ( 
.A(n_6992),
.B(n_222),
.Y(n_7304)
);

AND2x4_ASAP7_75t_L g7305 ( 
.A(n_6963),
.B(n_223),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6958),
.Y(n_7306)
);

AOI21xp5_ASAP7_75t_SL g7307 ( 
.A1(n_6967),
.A2(n_223),
.B(n_224),
.Y(n_7307)
);

AND2x2_ASAP7_75t_L g7308 ( 
.A(n_6917),
.B(n_224),
.Y(n_7308)
);

NAND2xp5_ASAP7_75t_L g7309 ( 
.A(n_7004),
.B(n_404),
.Y(n_7309)
);

OAI22xp5_ASAP7_75t_L g7310 ( 
.A1(n_6967),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_7310)
);

INVx1_ASAP7_75t_L g7311 ( 
.A(n_6958),
.Y(n_7311)
);

AOI21xp5_ASAP7_75t_SL g7312 ( 
.A1(n_6952),
.A2(n_225),
.B(n_226),
.Y(n_7312)
);

AND2x2_ASAP7_75t_L g7313 ( 
.A(n_6895),
.B(n_226),
.Y(n_7313)
);

HB1xp67_ASAP7_75t_L g7314 ( 
.A(n_6966),
.Y(n_7314)
);

OR2x2_ASAP7_75t_L g7315 ( 
.A(n_6895),
.B(n_227),
.Y(n_7315)
);

OA21x2_ASAP7_75t_L g7316 ( 
.A1(n_7106),
.A2(n_228),
.B(n_229),
.Y(n_7316)
);

AND2x2_ASAP7_75t_L g7317 ( 
.A(n_7004),
.B(n_228),
.Y(n_7317)
);

AOI21x1_ASAP7_75t_SL g7318 ( 
.A1(n_6920),
.A2(n_229),
.B(n_230),
.Y(n_7318)
);

A2O1A1Ixp33_ASAP7_75t_L g7319 ( 
.A1(n_7114),
.A2(n_232),
.B(n_230),
.C(n_231),
.Y(n_7319)
);

OA21x2_ASAP7_75t_L g7320 ( 
.A1(n_7108),
.A2(n_231),
.B(n_232),
.Y(n_7320)
);

INVx2_ASAP7_75t_L g7321 ( 
.A(n_7041),
.Y(n_7321)
);

AOI21xp5_ASAP7_75t_L g7322 ( 
.A1(n_7020),
.A2(n_232),
.B(n_233),
.Y(n_7322)
);

AND2x2_ASAP7_75t_L g7323 ( 
.A(n_6966),
.B(n_6968),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_6968),
.Y(n_7324)
);

BUFx3_ASAP7_75t_L g7325 ( 
.A(n_7028),
.Y(n_7325)
);

AOI21x1_ASAP7_75t_SL g7326 ( 
.A1(n_7022),
.A2(n_233),
.B(n_234),
.Y(n_7326)
);

AND2x2_ASAP7_75t_L g7327 ( 
.A(n_6990),
.B(n_233),
.Y(n_7327)
);

HB1xp67_ASAP7_75t_L g7328 ( 
.A(n_6990),
.Y(n_7328)
);

OAI22xp5_ASAP7_75t_L g7329 ( 
.A1(n_7107),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_7329)
);

NAND2xp5_ASAP7_75t_L g7330 ( 
.A(n_6983),
.B(n_405),
.Y(n_7330)
);

INVx2_ASAP7_75t_L g7331 ( 
.A(n_7045),
.Y(n_7331)
);

BUFx3_ASAP7_75t_L g7332 ( 
.A(n_7076),
.Y(n_7332)
);

OAI22xp5_ASAP7_75t_L g7333 ( 
.A1(n_7052),
.A2(n_237),
.B1(n_234),
.B2(n_235),
.Y(n_7333)
);

AOI21xp5_ASAP7_75t_SL g7334 ( 
.A1(n_6952),
.A2(n_235),
.B(n_237),
.Y(n_7334)
);

OA21x2_ASAP7_75t_L g7335 ( 
.A1(n_7108),
.A2(n_238),
.B(n_239),
.Y(n_7335)
);

OAI22xp5_ASAP7_75t_L g7336 ( 
.A1(n_7059),
.A2(n_240),
.B1(n_238),
.B2(n_239),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_7045),
.Y(n_7337)
);

O2A1O1Ixp33_ASAP7_75t_L g7338 ( 
.A1(n_6955),
.A2(n_241),
.B(n_238),
.C(n_240),
.Y(n_7338)
);

HB1xp67_ASAP7_75t_L g7339 ( 
.A(n_6921),
.Y(n_7339)
);

OA21x2_ASAP7_75t_L g7340 ( 
.A1(n_6868),
.A2(n_6870),
.B(n_6890),
.Y(n_7340)
);

INVx3_ASAP7_75t_L g7341 ( 
.A(n_6998),
.Y(n_7341)
);

AOI21xp5_ASAP7_75t_L g7342 ( 
.A1(n_7020),
.A2(n_241),
.B(n_242),
.Y(n_7342)
);

OR2x2_ASAP7_75t_L g7343 ( 
.A(n_7015),
.B(n_6921),
.Y(n_7343)
);

NAND2xp5_ASAP7_75t_L g7344 ( 
.A(n_7099),
.B(n_409),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_7073),
.B(n_242),
.Y(n_7345)
);

INVx1_ASAP7_75t_L g7346 ( 
.A(n_7129),
.Y(n_7346)
);

AND2x2_ASAP7_75t_L g7347 ( 
.A(n_7084),
.B(n_243),
.Y(n_7347)
);

AOI21x1_ASAP7_75t_SL g7348 ( 
.A1(n_7037),
.A2(n_243),
.B(n_244),
.Y(n_7348)
);

AND2x2_ASAP7_75t_L g7349 ( 
.A(n_7090),
.B(n_244),
.Y(n_7349)
);

INVxp67_ASAP7_75t_L g7350 ( 
.A(n_6980),
.Y(n_7350)
);

OA21x2_ASAP7_75t_L g7351 ( 
.A1(n_6898),
.A2(n_244),
.B(n_245),
.Y(n_7351)
);

NAND2xp5_ASAP7_75t_L g7352 ( 
.A(n_7099),
.B(n_410),
.Y(n_7352)
);

OAI22xp5_ASAP7_75t_L g7353 ( 
.A1(n_6899),
.A2(n_247),
.B1(n_245),
.B2(n_246),
.Y(n_7353)
);

INVx1_ASAP7_75t_L g7354 ( 
.A(n_7129),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_7129),
.Y(n_7355)
);

OA21x2_ASAP7_75t_L g7356 ( 
.A1(n_7030),
.A2(n_246),
.B(n_247),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_7099),
.B(n_411),
.Y(n_7357)
);

OR2x2_ASAP7_75t_L g7358 ( 
.A(n_7092),
.B(n_246),
.Y(n_7358)
);

AND2x4_ASAP7_75t_L g7359 ( 
.A(n_6974),
.B(n_247),
.Y(n_7359)
);

O2A1O1Ixp5_ASAP7_75t_L g7360 ( 
.A1(n_6984),
.A2(n_251),
.B(n_248),
.C(n_249),
.Y(n_7360)
);

O2A1O1Ixp5_ASAP7_75t_L g7361 ( 
.A1(n_7009),
.A2(n_251),
.B(n_248),
.C(n_249),
.Y(n_7361)
);

O2A1O1Ixp33_ASAP7_75t_L g7362 ( 
.A1(n_6891),
.A2(n_252),
.B(n_249),
.C(n_251),
.Y(n_7362)
);

HB1xp67_ASAP7_75t_L g7363 ( 
.A(n_6876),
.Y(n_7363)
);

AND2x2_ASAP7_75t_L g7364 ( 
.A(n_6954),
.B(n_252),
.Y(n_7364)
);

INVx2_ASAP7_75t_L g7365 ( 
.A(n_7123),
.Y(n_7365)
);

INVxp67_ASAP7_75t_L g7366 ( 
.A(n_7049),
.Y(n_7366)
);

O2A1O1Ixp5_ASAP7_75t_L g7367 ( 
.A1(n_7009),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_7367)
);

BUFx3_ASAP7_75t_L g7368 ( 
.A(n_7081),
.Y(n_7368)
);

OA21x2_ASAP7_75t_L g7369 ( 
.A1(n_7014),
.A2(n_253),
.B(n_254),
.Y(n_7369)
);

OAI22xp5_ASAP7_75t_L g7370 ( 
.A1(n_7061),
.A2(n_256),
.B1(n_253),
.B2(n_255),
.Y(n_7370)
);

AND2x2_ASAP7_75t_L g7371 ( 
.A(n_6998),
.B(n_256),
.Y(n_7371)
);

OR2x2_ASAP7_75t_L g7372 ( 
.A(n_7010),
.B(n_256),
.Y(n_7372)
);

AOI21xp5_ASAP7_75t_SL g7373 ( 
.A1(n_7124),
.A2(n_6938),
.B(n_6977),
.Y(n_7373)
);

AOI21xp5_ASAP7_75t_L g7374 ( 
.A1(n_7010),
.A2(n_257),
.B(n_258),
.Y(n_7374)
);

INVx2_ASAP7_75t_L g7375 ( 
.A(n_7123),
.Y(n_7375)
);

AND2x2_ASAP7_75t_L g7376 ( 
.A(n_6922),
.B(n_257),
.Y(n_7376)
);

NAND2xp5_ASAP7_75t_L g7377 ( 
.A(n_7018),
.B(n_412),
.Y(n_7377)
);

HB1xp67_ASAP7_75t_L g7378 ( 
.A(n_7008),
.Y(n_7378)
);

OAI22xp5_ASAP7_75t_L g7379 ( 
.A1(n_7016),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_7379)
);

INVx1_ASAP7_75t_SL g7380 ( 
.A(n_7032),
.Y(n_7380)
);

OR2x6_ASAP7_75t_L g7381 ( 
.A(n_7312),
.B(n_7034),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_7209),
.B(n_6965),
.Y(n_7382)
);

INVx2_ASAP7_75t_L g7383 ( 
.A(n_7351),
.Y(n_7383)
);

BUFx2_ASAP7_75t_L g7384 ( 
.A(n_7132),
.Y(n_7384)
);

INVx1_ASAP7_75t_L g7385 ( 
.A(n_7278),
.Y(n_7385)
);

BUFx2_ASAP7_75t_L g7386 ( 
.A(n_7161),
.Y(n_7386)
);

OAI21xp5_ASAP7_75t_L g7387 ( 
.A1(n_7290),
.A2(n_7080),
.B(n_7091),
.Y(n_7387)
);

HB1xp67_ASAP7_75t_L g7388 ( 
.A(n_7212),
.Y(n_7388)
);

INVx2_ASAP7_75t_L g7389 ( 
.A(n_7351),
.Y(n_7389)
);

OA21x2_ASAP7_75t_L g7390 ( 
.A1(n_7165),
.A2(n_7152),
.B(n_7160),
.Y(n_7390)
);

BUFx12f_ASAP7_75t_L g7391 ( 
.A(n_7194),
.Y(n_7391)
);

HB1xp67_ASAP7_75t_L g7392 ( 
.A(n_7216),
.Y(n_7392)
);

INVx2_ASAP7_75t_L g7393 ( 
.A(n_7358),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7314),
.Y(n_7394)
);

INVx1_ASAP7_75t_L g7395 ( 
.A(n_7328),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_7372),
.Y(n_7396)
);

HB1xp67_ASAP7_75t_L g7397 ( 
.A(n_7371),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_7316),
.Y(n_7398)
);

INVx2_ASAP7_75t_SL g7399 ( 
.A(n_7264),
.Y(n_7399)
);

AND2x4_ASAP7_75t_L g7400 ( 
.A(n_7200),
.B(n_7032),
.Y(n_7400)
);

AOI22xp33_ASAP7_75t_L g7401 ( 
.A1(n_7208),
.A2(n_7080),
.B1(n_7019),
.B2(n_6906),
.Y(n_7401)
);

OAI21x1_ASAP7_75t_L g7402 ( 
.A1(n_7341),
.A2(n_6910),
.B(n_6925),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_7316),
.Y(n_7403)
);

INVx2_ASAP7_75t_L g7404 ( 
.A(n_7264),
.Y(n_7404)
);

AO21x2_ASAP7_75t_L g7405 ( 
.A1(n_7154),
.A2(n_7021),
.B(n_7018),
.Y(n_7405)
);

OA21x2_ASAP7_75t_L g7406 ( 
.A1(n_7281),
.A2(n_7021),
.B(n_7027),
.Y(n_7406)
);

OAI21x1_ASAP7_75t_L g7407 ( 
.A1(n_7341),
.A2(n_6914),
.B(n_7070),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_7320),
.Y(n_7408)
);

INVx2_ASAP7_75t_L g7409 ( 
.A(n_7264),
.Y(n_7409)
);

INVx2_ASAP7_75t_L g7410 ( 
.A(n_7273),
.Y(n_7410)
);

INVx3_ASAP7_75t_L g7411 ( 
.A(n_7293),
.Y(n_7411)
);

INVx2_ASAP7_75t_L g7412 ( 
.A(n_7277),
.Y(n_7412)
);

INVx2_ASAP7_75t_L g7413 ( 
.A(n_7359),
.Y(n_7413)
);

AND2x2_ASAP7_75t_L g7414 ( 
.A(n_7200),
.B(n_6999),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_7320),
.Y(n_7415)
);

HB1xp67_ASAP7_75t_L g7416 ( 
.A(n_7133),
.Y(n_7416)
);

INVxp67_ASAP7_75t_L g7417 ( 
.A(n_7287),
.Y(n_7417)
);

INVx2_ASAP7_75t_L g7418 ( 
.A(n_7359),
.Y(n_7418)
);

OAI21x1_ASAP7_75t_L g7419 ( 
.A1(n_7172),
.A2(n_7070),
.B(n_6961),
.Y(n_7419)
);

BUFx3_ASAP7_75t_L g7420 ( 
.A(n_7223),
.Y(n_7420)
);

AO21x2_ASAP7_75t_L g7421 ( 
.A1(n_7251),
.A2(n_7038),
.B(n_7027),
.Y(n_7421)
);

AND2x2_ASAP7_75t_L g7422 ( 
.A(n_7144),
.B(n_7007),
.Y(n_7422)
);

AND2x4_ASAP7_75t_L g7423 ( 
.A(n_7176),
.B(n_7032),
.Y(n_7423)
);

AND2x2_ASAP7_75t_L g7424 ( 
.A(n_7158),
.B(n_7040),
.Y(n_7424)
);

OR2x6_ASAP7_75t_L g7425 ( 
.A(n_7334),
.B(n_7034),
.Y(n_7425)
);

HB1xp67_ASAP7_75t_L g7426 ( 
.A(n_7133),
.Y(n_7426)
);

INVx2_ASAP7_75t_L g7427 ( 
.A(n_7288),
.Y(n_7427)
);

BUFx2_ASAP7_75t_L g7428 ( 
.A(n_7176),
.Y(n_7428)
);

INVx2_ASAP7_75t_L g7429 ( 
.A(n_7288),
.Y(n_7429)
);

AND2x4_ASAP7_75t_L g7430 ( 
.A(n_7193),
.B(n_7139),
.Y(n_7430)
);

AO21x2_ASAP7_75t_L g7431 ( 
.A1(n_7253),
.A2(n_7038),
.B(n_6945),
.Y(n_7431)
);

HB1xp67_ASAP7_75t_L g7432 ( 
.A(n_7169),
.Y(n_7432)
);

OR2x2_ASAP7_75t_L g7433 ( 
.A(n_7130),
.B(n_6938),
.Y(n_7433)
);

INVx1_ASAP7_75t_L g7434 ( 
.A(n_7335),
.Y(n_7434)
);

AND2x2_ASAP7_75t_L g7435 ( 
.A(n_7159),
.B(n_6994),
.Y(n_7435)
);

OR2x2_ASAP7_75t_L g7436 ( 
.A(n_7140),
.B(n_6970),
.Y(n_7436)
);

INVx1_ASAP7_75t_L g7437 ( 
.A(n_7335),
.Y(n_7437)
);

HB1xp67_ASAP7_75t_SL g7438 ( 
.A(n_7244),
.Y(n_7438)
);

HB1xp67_ASAP7_75t_L g7439 ( 
.A(n_7145),
.Y(n_7439)
);

AND2x2_ASAP7_75t_L g7440 ( 
.A(n_7170),
.B(n_7095),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_7337),
.Y(n_7441)
);

AO21x2_ASAP7_75t_L g7442 ( 
.A1(n_7274),
.A2(n_6945),
.B(n_6924),
.Y(n_7442)
);

AND2x4_ASAP7_75t_SL g7443 ( 
.A(n_7260),
.B(n_7245),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_7284),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_7302),
.Y(n_7445)
);

AOI21xp5_ASAP7_75t_SL g7446 ( 
.A1(n_7166),
.A2(n_7124),
.B(n_6977),
.Y(n_7446)
);

INVx1_ASAP7_75t_L g7447 ( 
.A(n_7256),
.Y(n_7447)
);

AOI22xp33_ASAP7_75t_L g7448 ( 
.A1(n_7142),
.A2(n_6906),
.B1(n_6970),
.B2(n_7056),
.Y(n_7448)
);

BUFx2_ASAP7_75t_L g7449 ( 
.A(n_7193),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_7256),
.Y(n_7450)
);

HB1xp67_ASAP7_75t_L g7451 ( 
.A(n_7378),
.Y(n_7451)
);

INVx1_ASAP7_75t_L g7452 ( 
.A(n_7275),
.Y(n_7452)
);

BUFx3_ASAP7_75t_L g7453 ( 
.A(n_7195),
.Y(n_7453)
);

INVx2_ASAP7_75t_L g7454 ( 
.A(n_7376),
.Y(n_7454)
);

INVx1_ASAP7_75t_SL g7455 ( 
.A(n_7147),
.Y(n_7455)
);

AND2x4_ASAP7_75t_L g7456 ( 
.A(n_7163),
.B(n_7143),
.Y(n_7456)
);

AO21x2_ASAP7_75t_L g7457 ( 
.A1(n_7339),
.A2(n_6993),
.B(n_6986),
.Y(n_7457)
);

BUFx2_ASAP7_75t_L g7458 ( 
.A(n_7230),
.Y(n_7458)
);

AND2x2_ASAP7_75t_L g7459 ( 
.A(n_7175),
.B(n_6916),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7275),
.Y(n_7460)
);

INVx2_ASAP7_75t_L g7461 ( 
.A(n_7305),
.Y(n_7461)
);

OAI21x1_ASAP7_75t_L g7462 ( 
.A1(n_7205),
.A2(n_6887),
.B(n_7126),
.Y(n_7462)
);

INVx2_ASAP7_75t_L g7463 ( 
.A(n_7305),
.Y(n_7463)
);

AND2x4_ASAP7_75t_L g7464 ( 
.A(n_7153),
.B(n_6939),
.Y(n_7464)
);

OR2x6_ASAP7_75t_L g7465 ( 
.A(n_7183),
.B(n_7031),
.Y(n_7465)
);

INVx2_ASAP7_75t_L g7466 ( 
.A(n_7211),
.Y(n_7466)
);

AO21x2_ASAP7_75t_L g7467 ( 
.A1(n_7136),
.A2(n_7082),
.B(n_7087),
.Y(n_7467)
);

INVx3_ASAP7_75t_L g7468 ( 
.A(n_7259),
.Y(n_7468)
);

INVx2_ASAP7_75t_L g7469 ( 
.A(n_7213),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_7134),
.Y(n_7470)
);

BUFx3_ASAP7_75t_L g7471 ( 
.A(n_7265),
.Y(n_7471)
);

AND2x4_ASAP7_75t_L g7472 ( 
.A(n_7240),
.B(n_7025),
.Y(n_7472)
);

OA21x2_ASAP7_75t_L g7473 ( 
.A1(n_7151),
.A2(n_6972),
.B(n_6878),
.Y(n_7473)
);

INVx1_ASAP7_75t_L g7474 ( 
.A(n_7135),
.Y(n_7474)
);

HB1xp67_ASAP7_75t_L g7475 ( 
.A(n_7295),
.Y(n_7475)
);

INVx3_ASAP7_75t_L g7476 ( 
.A(n_7259),
.Y(n_7476)
);

INVx2_ASAP7_75t_L g7477 ( 
.A(n_7217),
.Y(n_7477)
);

INVx1_ASAP7_75t_L g7478 ( 
.A(n_7138),
.Y(n_7478)
);

BUFx2_ASAP7_75t_L g7479 ( 
.A(n_7332),
.Y(n_7479)
);

INVx1_ASAP7_75t_L g7480 ( 
.A(n_7178),
.Y(n_7480)
);

NAND2xp5_ASAP7_75t_L g7481 ( 
.A(n_7162),
.B(n_7026),
.Y(n_7481)
);

NAND2xp5_ASAP7_75t_L g7482 ( 
.A(n_7323),
.B(n_7048),
.Y(n_7482)
);

INVx1_ASAP7_75t_L g7483 ( 
.A(n_7185),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_7186),
.Y(n_7484)
);

AND2x2_ASAP7_75t_L g7485 ( 
.A(n_7226),
.B(n_7089),
.Y(n_7485)
);

AND2x2_ASAP7_75t_L g7486 ( 
.A(n_7232),
.B(n_7060),
.Y(n_7486)
);

INVx2_ASAP7_75t_L g7487 ( 
.A(n_7221),
.Y(n_7487)
);

INVx3_ASAP7_75t_L g7488 ( 
.A(n_7304),
.Y(n_7488)
);

INVx2_ASAP7_75t_SL g7489 ( 
.A(n_7304),
.Y(n_7489)
);

INVx2_ASAP7_75t_L g7490 ( 
.A(n_7365),
.Y(n_7490)
);

INVx2_ASAP7_75t_L g7491 ( 
.A(n_7375),
.Y(n_7491)
);

INVx1_ASAP7_75t_L g7492 ( 
.A(n_7242),
.Y(n_7492)
);

NAND2x1_ASAP7_75t_L g7493 ( 
.A(n_7373),
.B(n_6971),
.Y(n_7493)
);

OA21x2_ASAP7_75t_L g7494 ( 
.A1(n_7190),
.A2(n_6960),
.B(n_6946),
.Y(n_7494)
);

INVx1_ASAP7_75t_L g7495 ( 
.A(n_7249),
.Y(n_7495)
);

INVx1_ASAP7_75t_SL g7496 ( 
.A(n_7325),
.Y(n_7496)
);

BUFx3_ASAP7_75t_L g7497 ( 
.A(n_7268),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_7261),
.Y(n_7498)
);

INVx1_ASAP7_75t_L g7499 ( 
.A(n_7263),
.Y(n_7499)
);

HB1xp67_ASAP7_75t_L g7500 ( 
.A(n_7295),
.Y(n_7500)
);

BUFx8_ASAP7_75t_SL g7501 ( 
.A(n_7364),
.Y(n_7501)
);

INVxp67_ASAP7_75t_L g7502 ( 
.A(n_7377),
.Y(n_7502)
);

BUFx6f_ASAP7_75t_L g7503 ( 
.A(n_7243),
.Y(n_7503)
);

INVx1_ASAP7_75t_L g7504 ( 
.A(n_7279),
.Y(n_7504)
);

OA21x2_ASAP7_75t_L g7505 ( 
.A1(n_7224),
.A2(n_6976),
.B(n_6900),
.Y(n_7505)
);

AO31x2_ASAP7_75t_L g7506 ( 
.A1(n_7228),
.A2(n_6875),
.A3(n_7105),
.B(n_7078),
.Y(n_7506)
);

INVx2_ASAP7_75t_L g7507 ( 
.A(n_7199),
.Y(n_7507)
);

INVxp33_ASAP7_75t_L g7508 ( 
.A(n_7198),
.Y(n_7508)
);

INVx2_ASAP7_75t_L g7509 ( 
.A(n_7199),
.Y(n_7509)
);

AND2x4_ASAP7_75t_L g7510 ( 
.A(n_7192),
.B(n_7068),
.Y(n_7510)
);

HB1xp67_ASAP7_75t_L g7511 ( 
.A(n_7369),
.Y(n_7511)
);

INVx1_ASAP7_75t_L g7512 ( 
.A(n_7280),
.Y(n_7512)
);

BUFx3_ASAP7_75t_L g7513 ( 
.A(n_7268),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7282),
.Y(n_7514)
);

OAI21x1_ASAP7_75t_L g7515 ( 
.A1(n_7299),
.A2(n_6896),
.B(n_6978),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_7306),
.Y(n_7516)
);

INVx2_ASAP7_75t_L g7517 ( 
.A(n_7356),
.Y(n_7517)
);

AOI22xp33_ASAP7_75t_L g7518 ( 
.A1(n_7142),
.A2(n_7079),
.B1(n_6882),
.B2(n_7078),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_7311),
.Y(n_7519)
);

INVx2_ASAP7_75t_L g7520 ( 
.A(n_7356),
.Y(n_7520)
);

NAND2xp5_ASAP7_75t_L g7521 ( 
.A(n_7296),
.B(n_6971),
.Y(n_7521)
);

INVx1_ASAP7_75t_L g7522 ( 
.A(n_7324),
.Y(n_7522)
);

HB1xp67_ASAP7_75t_L g7523 ( 
.A(n_7369),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_7315),
.Y(n_7524)
);

BUFx3_ASAP7_75t_L g7525 ( 
.A(n_7289),
.Y(n_7525)
);

INVx1_ASAP7_75t_L g7526 ( 
.A(n_7301),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7321),
.Y(n_7527)
);

AND2x2_ASAP7_75t_L g7528 ( 
.A(n_7202),
.B(n_6877),
.Y(n_7528)
);

INVx2_ASAP7_75t_L g7529 ( 
.A(n_7171),
.Y(n_7529)
);

NAND2x1_ASAP7_75t_L g7530 ( 
.A(n_7180),
.B(n_7157),
.Y(n_7530)
);

INVx2_ASAP7_75t_L g7531 ( 
.A(n_7171),
.Y(n_7531)
);

INVx1_ASAP7_75t_L g7532 ( 
.A(n_7331),
.Y(n_7532)
);

INVx1_ASAP7_75t_L g7533 ( 
.A(n_7344),
.Y(n_7533)
);

AO21x2_ASAP7_75t_L g7534 ( 
.A1(n_7191),
.A2(n_7103),
.B(n_7096),
.Y(n_7534)
);

AND2x2_ASAP7_75t_L g7535 ( 
.A(n_7350),
.B(n_7033),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7352),
.Y(n_7536)
);

INVx1_ASAP7_75t_L g7537 ( 
.A(n_7357),
.Y(n_7537)
);

HB1xp67_ASAP7_75t_L g7538 ( 
.A(n_7294),
.Y(n_7538)
);

AO21x2_ASAP7_75t_L g7539 ( 
.A1(n_7214),
.A2(n_6892),
.B(n_7044),
.Y(n_7539)
);

INVx1_ASAP7_75t_L g7540 ( 
.A(n_7317),
.Y(n_7540)
);

OAI21x1_ASAP7_75t_L g7541 ( 
.A1(n_7215),
.A2(n_6979),
.B(n_6981),
.Y(n_7541)
);

INVx1_ASAP7_75t_L g7542 ( 
.A(n_7327),
.Y(n_7542)
);

AND2x2_ASAP7_75t_L g7543 ( 
.A(n_7313),
.B(n_7104),
.Y(n_7543)
);

OR2x2_ASAP7_75t_L g7544 ( 
.A(n_7241),
.B(n_7105),
.Y(n_7544)
);

OAI21x1_ASAP7_75t_L g7545 ( 
.A1(n_7227),
.A2(n_7109),
.B(n_7115),
.Y(n_7545)
);

AND2x2_ASAP7_75t_L g7546 ( 
.A(n_7380),
.B(n_7112),
.Y(n_7546)
);

INVx2_ASAP7_75t_L g7547 ( 
.A(n_7294),
.Y(n_7547)
);

OA21x2_ASAP7_75t_L g7548 ( 
.A1(n_7141),
.A2(n_7054),
.B(n_7117),
.Y(n_7548)
);

INVx2_ASAP7_75t_L g7549 ( 
.A(n_7149),
.Y(n_7549)
);

INVx3_ASAP7_75t_L g7550 ( 
.A(n_7233),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7174),
.Y(n_7551)
);

INVx1_ASAP7_75t_L g7552 ( 
.A(n_7189),
.Y(n_7552)
);

INVx2_ASAP7_75t_L g7553 ( 
.A(n_7149),
.Y(n_7553)
);

INVx2_ASAP7_75t_L g7554 ( 
.A(n_7366),
.Y(n_7554)
);

OR2x2_ASAP7_75t_L g7555 ( 
.A(n_7148),
.B(n_7115),
.Y(n_7555)
);

INVx1_ASAP7_75t_L g7556 ( 
.A(n_7309),
.Y(n_7556)
);

INVx1_ASAP7_75t_L g7557 ( 
.A(n_7346),
.Y(n_7557)
);

INVx1_ASAP7_75t_L g7558 ( 
.A(n_7354),
.Y(n_7558)
);

INVx3_ASAP7_75t_L g7559 ( 
.A(n_7233),
.Y(n_7559)
);

HB1xp67_ASAP7_75t_L g7560 ( 
.A(n_7363),
.Y(n_7560)
);

INVx2_ASAP7_75t_L g7561 ( 
.A(n_7340),
.Y(n_7561)
);

INVx3_ASAP7_75t_L g7562 ( 
.A(n_7380),
.Y(n_7562)
);

OR2x2_ASAP7_75t_L g7563 ( 
.A(n_7207),
.B(n_7122),
.Y(n_7563)
);

INVx1_ASAP7_75t_SL g7564 ( 
.A(n_7270),
.Y(n_7564)
);

OR2x2_ASAP7_75t_L g7565 ( 
.A(n_7187),
.B(n_7122),
.Y(n_7565)
);

AO21x2_ASAP7_75t_L g7566 ( 
.A1(n_7300),
.A2(n_7121),
.B(n_7109),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_7355),
.Y(n_7567)
);

AO21x2_ASAP7_75t_L g7568 ( 
.A1(n_7343),
.A2(n_6882),
.B(n_6886),
.Y(n_7568)
);

INVx2_ASAP7_75t_L g7569 ( 
.A(n_7340),
.Y(n_7569)
);

INVx2_ASAP7_75t_L g7570 ( 
.A(n_7167),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_7203),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7330),
.Y(n_7572)
);

INVx2_ASAP7_75t_L g7573 ( 
.A(n_7167),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_7310),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_7345),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7347),
.Y(n_7576)
);

INVxp67_ASAP7_75t_L g7577 ( 
.A(n_7353),
.Y(n_7577)
);

INVx6_ASAP7_75t_SL g7578 ( 
.A(n_7285),
.Y(n_7578)
);

INVx2_ASAP7_75t_L g7579 ( 
.A(n_7368),
.Y(n_7579)
);

OR2x6_ASAP7_75t_L g7580 ( 
.A(n_7307),
.B(n_6886),
.Y(n_7580)
);

OAI21xp5_ASAP7_75t_L g7581 ( 
.A1(n_7362),
.A2(n_258),
.B(n_259),
.Y(n_7581)
);

INVx2_ASAP7_75t_L g7582 ( 
.A(n_7349),
.Y(n_7582)
);

INVx1_ASAP7_75t_L g7583 ( 
.A(n_7361),
.Y(n_7583)
);

INVx1_ASAP7_75t_L g7584 ( 
.A(n_7367),
.Y(n_7584)
);

OAI21x1_ASAP7_75t_L g7585 ( 
.A1(n_7227),
.A2(n_260),
.B(n_262),
.Y(n_7585)
);

HB1xp67_ASAP7_75t_L g7586 ( 
.A(n_7168),
.Y(n_7586)
);

INVx2_ASAP7_75t_L g7587 ( 
.A(n_7292),
.Y(n_7587)
);

OAI21xp5_ASAP7_75t_L g7588 ( 
.A1(n_7269),
.A2(n_260),
.B(n_263),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_7137),
.Y(n_7589)
);

NAND2xp5_ASAP7_75t_L g7590 ( 
.A(n_7179),
.B(n_263),
.Y(n_7590)
);

AND2x2_ASAP7_75t_L g7591 ( 
.A(n_7234),
.B(n_264),
.Y(n_7591)
);

INVx2_ASAP7_75t_L g7592 ( 
.A(n_7237),
.Y(n_7592)
);

HB1xp67_ASAP7_75t_L g7593 ( 
.A(n_7225),
.Y(n_7593)
);

HB1xp67_ASAP7_75t_L g7594 ( 
.A(n_7184),
.Y(n_7594)
);

NOR2xp33_ASAP7_75t_L g7595 ( 
.A(n_7267),
.B(n_264),
.Y(n_7595)
);

INVx3_ASAP7_75t_L g7596 ( 
.A(n_7182),
.Y(n_7596)
);

INVxp67_ASAP7_75t_L g7597 ( 
.A(n_7246),
.Y(n_7597)
);

INVx1_ASAP7_75t_L g7598 ( 
.A(n_7298),
.Y(n_7598)
);

INVx2_ASAP7_75t_L g7599 ( 
.A(n_7257),
.Y(n_7599)
);

HB1xp67_ASAP7_75t_L g7600 ( 
.A(n_7184),
.Y(n_7600)
);

INVx2_ASAP7_75t_L g7601 ( 
.A(n_7258),
.Y(n_7601)
);

NAND2xp5_ASAP7_75t_L g7602 ( 
.A(n_7146),
.B(n_265),
.Y(n_7602)
);

OR2x6_ASAP7_75t_L g7603 ( 
.A(n_7322),
.B(n_265),
.Y(n_7603)
);

OR2x2_ASAP7_75t_L g7604 ( 
.A(n_7131),
.B(n_7173),
.Y(n_7604)
);

INVx1_ASAP7_75t_L g7605 ( 
.A(n_7197),
.Y(n_7605)
);

INVx1_ASAP7_75t_L g7606 ( 
.A(n_7229),
.Y(n_7606)
);

NAND2xp5_ASAP7_75t_L g7607 ( 
.A(n_7181),
.B(n_266),
.Y(n_7607)
);

INVx1_ASAP7_75t_L g7608 ( 
.A(n_7238),
.Y(n_7608)
);

INVx2_ASAP7_75t_L g7609 ( 
.A(n_7196),
.Y(n_7609)
);

AO31x2_ASAP7_75t_L g7610 ( 
.A1(n_7218),
.A2(n_268),
.A3(n_266),
.B(n_267),
.Y(n_7610)
);

INVx2_ASAP7_75t_L g7611 ( 
.A(n_7308),
.Y(n_7611)
);

AND2x4_ASAP7_75t_L g7612 ( 
.A(n_7192),
.B(n_266),
.Y(n_7612)
);

INVx3_ASAP7_75t_L g7613 ( 
.A(n_7204),
.Y(n_7613)
);

HB1xp67_ASAP7_75t_L g7614 ( 
.A(n_7206),
.Y(n_7614)
);

INVx3_ASAP7_75t_L g7615 ( 
.A(n_7220),
.Y(n_7615)
);

AND2x2_ASAP7_75t_L g7616 ( 
.A(n_7430),
.B(n_7164),
.Y(n_7616)
);

OA21x2_ASAP7_75t_L g7617 ( 
.A1(n_7614),
.A2(n_7210),
.B(n_7231),
.Y(n_7617)
);

AND2x4_ASAP7_75t_L g7618 ( 
.A(n_7430),
.B(n_7342),
.Y(n_7618)
);

AOI22xp33_ASAP7_75t_L g7619 ( 
.A1(n_7580),
.A2(n_7206),
.B1(n_7219),
.B2(n_7276),
.Y(n_7619)
);

INVxp67_ASAP7_75t_L g7620 ( 
.A(n_7501),
.Y(n_7620)
);

INVx2_ASAP7_75t_SL g7621 ( 
.A(n_7443),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7432),
.Y(n_7622)
);

NAND2xp5_ASAP7_75t_L g7623 ( 
.A(n_7401),
.B(n_7150),
.Y(n_7623)
);

AND2x2_ASAP7_75t_L g7624 ( 
.A(n_7428),
.B(n_7303),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7432),
.Y(n_7625)
);

AND2x2_ASAP7_75t_L g7626 ( 
.A(n_7449),
.B(n_7177),
.Y(n_7626)
);

A2O1A1Ixp33_ASAP7_75t_L g7627 ( 
.A1(n_7614),
.A2(n_7150),
.B(n_7338),
.C(n_7252),
.Y(n_7627)
);

INVx1_ASAP7_75t_L g7628 ( 
.A(n_7439),
.Y(n_7628)
);

NOR2x1_ASAP7_75t_SL g7629 ( 
.A(n_7465),
.B(n_7156),
.Y(n_7629)
);

OAI21xp5_ASAP7_75t_L g7630 ( 
.A1(n_7521),
.A2(n_7283),
.B(n_7272),
.Y(n_7630)
);

INVx2_ASAP7_75t_L g7631 ( 
.A(n_7453),
.Y(n_7631)
);

AOI21xp5_ASAP7_75t_L g7632 ( 
.A1(n_7521),
.A2(n_7271),
.B(n_7222),
.Y(n_7632)
);

AO32x2_ASAP7_75t_L g7633 ( 
.A1(n_7489),
.A2(n_7329),
.A3(n_7222),
.B1(n_7336),
.B2(n_7333),
.Y(n_7633)
);

INVx2_ASAP7_75t_L g7634 ( 
.A(n_7453),
.Y(n_7634)
);

NOR2x1_ASAP7_75t_SL g7635 ( 
.A(n_7465),
.B(n_7250),
.Y(n_7635)
);

INVx1_ASAP7_75t_L g7636 ( 
.A(n_7439),
.Y(n_7636)
);

INVx3_ASAP7_75t_L g7637 ( 
.A(n_7420),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_7525),
.Y(n_7638)
);

OR2x6_ASAP7_75t_L g7639 ( 
.A(n_7384),
.B(n_7248),
.Y(n_7639)
);

CKINVDCx5p33_ASAP7_75t_R g7640 ( 
.A(n_7420),
.Y(n_7640)
);

AOI221xp5_ASAP7_75t_L g7641 ( 
.A1(n_7571),
.A2(n_7247),
.B1(n_7286),
.B2(n_7374),
.C(n_7255),
.Y(n_7641)
);

INVx1_ASAP7_75t_L g7642 ( 
.A(n_7526),
.Y(n_7642)
);

NAND2xp5_ASAP7_75t_L g7643 ( 
.A(n_7401),
.B(n_7250),
.Y(n_7643)
);

NOR2x1_ASAP7_75t_R g7644 ( 
.A(n_7386),
.B(n_7291),
.Y(n_7644)
);

OAI21xp5_ASAP7_75t_L g7645 ( 
.A1(n_7590),
.A2(n_7360),
.B(n_7319),
.Y(n_7645)
);

BUFx3_ASAP7_75t_L g7646 ( 
.A(n_7391),
.Y(n_7646)
);

OR2x2_ASAP7_75t_L g7647 ( 
.A(n_7397),
.B(n_7254),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_7527),
.Y(n_7648)
);

NAND2xp5_ASAP7_75t_L g7649 ( 
.A(n_7583),
.B(n_7254),
.Y(n_7649)
);

AND2x2_ASAP7_75t_L g7650 ( 
.A(n_7455),
.B(n_7201),
.Y(n_7650)
);

NAND2xp5_ASAP7_75t_L g7651 ( 
.A(n_7584),
.B(n_7262),
.Y(n_7651)
);

A2O1A1Ixp33_ASAP7_75t_L g7652 ( 
.A1(n_7511),
.A2(n_7201),
.B(n_7188),
.C(n_7370),
.Y(n_7652)
);

INVx2_ASAP7_75t_L g7653 ( 
.A(n_7503),
.Y(n_7653)
);

AND2x2_ASAP7_75t_L g7654 ( 
.A(n_7455),
.B(n_7262),
.Y(n_7654)
);

OR2x2_ASAP7_75t_L g7655 ( 
.A(n_7397),
.B(n_7236),
.Y(n_7655)
);

INVx3_ASAP7_75t_L g7656 ( 
.A(n_7578),
.Y(n_7656)
);

AOI22xp33_ASAP7_75t_SL g7657 ( 
.A1(n_7511),
.A2(n_7379),
.B1(n_7318),
.B2(n_7297),
.Y(n_7657)
);

AND2x2_ASAP7_75t_L g7658 ( 
.A(n_7458),
.B(n_7155),
.Y(n_7658)
);

AND2x2_ASAP7_75t_SL g7659 ( 
.A(n_7390),
.B(n_7326),
.Y(n_7659)
);

A2O1A1Ixp33_ASAP7_75t_L g7660 ( 
.A1(n_7523),
.A2(n_7239),
.B(n_7348),
.C(n_7266),
.Y(n_7660)
);

NOR2xp33_ASAP7_75t_L g7661 ( 
.A(n_7438),
.B(n_7235),
.Y(n_7661)
);

AOI21xp5_ASAP7_75t_L g7662 ( 
.A1(n_7481),
.A2(n_7239),
.B(n_267),
.Y(n_7662)
);

AND2x2_ASAP7_75t_L g7663 ( 
.A(n_7400),
.B(n_268),
.Y(n_7663)
);

OAI22xp5_ASAP7_75t_L g7664 ( 
.A1(n_7597),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_7664)
);

NAND2xp33_ASAP7_75t_L g7665 ( 
.A(n_7411),
.B(n_269),
.Y(n_7665)
);

AND2x2_ASAP7_75t_L g7666 ( 
.A(n_7400),
.B(n_7404),
.Y(n_7666)
);

INVx4_ASAP7_75t_SL g7667 ( 
.A(n_7471),
.Y(n_7667)
);

AND2x2_ASAP7_75t_L g7668 ( 
.A(n_7409),
.B(n_270),
.Y(n_7668)
);

AND2x2_ASAP7_75t_L g7669 ( 
.A(n_7410),
.B(n_270),
.Y(n_7669)
);

A2O1A1Ixp33_ASAP7_75t_L g7670 ( 
.A1(n_7523),
.A2(n_274),
.B(n_271),
.C(n_273),
.Y(n_7670)
);

NOR2xp33_ASAP7_75t_L g7671 ( 
.A(n_7438),
.B(n_271),
.Y(n_7671)
);

AND2x2_ASAP7_75t_L g7672 ( 
.A(n_7412),
.B(n_273),
.Y(n_7672)
);

INVx3_ASAP7_75t_SL g7673 ( 
.A(n_7411),
.Y(n_7673)
);

AO21x2_ASAP7_75t_L g7674 ( 
.A1(n_7590),
.A2(n_274),
.B(n_275),
.Y(n_7674)
);

NOR2xp33_ASAP7_75t_L g7675 ( 
.A(n_7501),
.B(n_274),
.Y(n_7675)
);

OAI21xp5_ASAP7_75t_L g7676 ( 
.A1(n_7607),
.A2(n_275),
.B(n_276),
.Y(n_7676)
);

AND2x2_ASAP7_75t_L g7677 ( 
.A(n_7440),
.B(n_275),
.Y(n_7677)
);

AND2x4_ASAP7_75t_L g7678 ( 
.A(n_7468),
.B(n_276),
.Y(n_7678)
);

NAND2xp5_ASAP7_75t_L g7679 ( 
.A(n_7496),
.B(n_277),
.Y(n_7679)
);

AND2x2_ASAP7_75t_L g7680 ( 
.A(n_7399),
.B(n_277),
.Y(n_7680)
);

AND2x2_ASAP7_75t_L g7681 ( 
.A(n_7456),
.B(n_277),
.Y(n_7681)
);

INVx1_ASAP7_75t_L g7682 ( 
.A(n_7532),
.Y(n_7682)
);

OAI21xp5_ASAP7_75t_L g7683 ( 
.A1(n_7607),
.A2(n_278),
.B(n_279),
.Y(n_7683)
);

OR2x2_ASAP7_75t_L g7684 ( 
.A(n_7427),
.B(n_279),
.Y(n_7684)
);

AOI21xp5_ASAP7_75t_L g7685 ( 
.A1(n_7481),
.A2(n_279),
.B(n_280),
.Y(n_7685)
);

BUFx8_ASAP7_75t_SL g7686 ( 
.A(n_7479),
.Y(n_7686)
);

NOR2xp33_ASAP7_75t_L g7687 ( 
.A(n_7496),
.B(n_280),
.Y(n_7687)
);

OAI22xp5_ASAP7_75t_L g7688 ( 
.A1(n_7597),
.A2(n_7580),
.B1(n_7493),
.B2(n_7564),
.Y(n_7688)
);

INVx1_ASAP7_75t_L g7689 ( 
.A(n_7398),
.Y(n_7689)
);

INVx3_ASAP7_75t_L g7690 ( 
.A(n_7578),
.Y(n_7690)
);

OR2x6_ASAP7_75t_L g7691 ( 
.A(n_7554),
.B(n_281),
.Y(n_7691)
);

BUFx6f_ASAP7_75t_L g7692 ( 
.A(n_7612),
.Y(n_7692)
);

AND2x4_ASAP7_75t_L g7693 ( 
.A(n_7497),
.B(n_281),
.Y(n_7693)
);

AO21x2_ASAP7_75t_L g7694 ( 
.A1(n_7416),
.A2(n_281),
.B(n_282),
.Y(n_7694)
);

NAND2xp5_ASAP7_75t_SL g7695 ( 
.A(n_7503),
.B(n_1751),
.Y(n_7695)
);

OAI21x1_ASAP7_75t_SL g7696 ( 
.A1(n_7602),
.A2(n_7390),
.B(n_7454),
.Y(n_7696)
);

AND2x2_ASAP7_75t_L g7697 ( 
.A(n_7456),
.B(n_282),
.Y(n_7697)
);

AO32x2_ASAP7_75t_L g7698 ( 
.A1(n_7417),
.A2(n_7577),
.A3(n_7605),
.B1(n_7502),
.B2(n_7444),
.Y(n_7698)
);

NAND2xp5_ASAP7_75t_L g7699 ( 
.A(n_7540),
.B(n_282),
.Y(n_7699)
);

OR2x2_ASAP7_75t_L g7700 ( 
.A(n_7429),
.B(n_283),
.Y(n_7700)
);

OAI22xp5_ASAP7_75t_L g7701 ( 
.A1(n_7580),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.Y(n_7701)
);

OR2x6_ASAP7_75t_L g7702 ( 
.A(n_7602),
.B(n_283),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7403),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7408),
.Y(n_7704)
);

AND2x2_ASAP7_75t_L g7705 ( 
.A(n_7424),
.B(n_284),
.Y(n_7705)
);

AND2x2_ASAP7_75t_L g7706 ( 
.A(n_7435),
.B(n_284),
.Y(n_7706)
);

NAND2xp33_ASAP7_75t_L g7707 ( 
.A(n_7564),
.B(n_285),
.Y(n_7707)
);

AOI22xp5_ASAP7_75t_L g7708 ( 
.A1(n_7577),
.A2(n_2959),
.B1(n_2985),
.B2(n_2895),
.Y(n_7708)
);

INVxp67_ASAP7_75t_L g7709 ( 
.A(n_7503),
.Y(n_7709)
);

AO21x2_ASAP7_75t_L g7710 ( 
.A1(n_7416),
.A2(n_285),
.B(n_286),
.Y(n_7710)
);

NOR2xp33_ASAP7_75t_L g7711 ( 
.A(n_7468),
.B(n_286),
.Y(n_7711)
);

INVx3_ASAP7_75t_L g7712 ( 
.A(n_7513),
.Y(n_7712)
);

OA21x2_ASAP7_75t_L g7713 ( 
.A1(n_7594),
.A2(n_287),
.B(n_288),
.Y(n_7713)
);

OAI22xp5_ASAP7_75t_L g7714 ( 
.A1(n_7475),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_7714)
);

OR2x6_ASAP7_75t_L g7715 ( 
.A(n_7612),
.B(n_287),
.Y(n_7715)
);

A2O1A1Ixp33_ASAP7_75t_L g7716 ( 
.A1(n_7538),
.A2(n_291),
.B(n_289),
.C(n_290),
.Y(n_7716)
);

INVx1_ASAP7_75t_L g7717 ( 
.A(n_7415),
.Y(n_7717)
);

OR2x6_ASAP7_75t_L g7718 ( 
.A(n_7611),
.B(n_290),
.Y(n_7718)
);

OA21x2_ASAP7_75t_L g7719 ( 
.A1(n_7594),
.A2(n_290),
.B(n_291),
.Y(n_7719)
);

AND2x4_ASAP7_75t_L g7720 ( 
.A(n_7476),
.B(n_291),
.Y(n_7720)
);

AND2x2_ASAP7_75t_L g7721 ( 
.A(n_7422),
.B(n_292),
.Y(n_7721)
);

CKINVDCx5p33_ASAP7_75t_R g7722 ( 
.A(n_7595),
.Y(n_7722)
);

AND2x2_ASAP7_75t_L g7723 ( 
.A(n_7591),
.B(n_292),
.Y(n_7723)
);

OA21x2_ASAP7_75t_L g7724 ( 
.A1(n_7600),
.A2(n_7437),
.B(n_7434),
.Y(n_7724)
);

NAND2xp5_ASAP7_75t_L g7725 ( 
.A(n_7542),
.B(n_293),
.Y(n_7725)
);

AND2x2_ASAP7_75t_L g7726 ( 
.A(n_7423),
.B(n_293),
.Y(n_7726)
);

NOR2xp33_ASAP7_75t_L g7727 ( 
.A(n_7476),
.B(n_293),
.Y(n_7727)
);

INVx3_ASAP7_75t_L g7728 ( 
.A(n_7488),
.Y(n_7728)
);

AND2x2_ASAP7_75t_L g7729 ( 
.A(n_7423),
.B(n_294),
.Y(n_7729)
);

NAND2xp5_ASAP7_75t_L g7730 ( 
.A(n_7417),
.B(n_294),
.Y(n_7730)
);

NAND2xp5_ASAP7_75t_L g7731 ( 
.A(n_7608),
.B(n_294),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7447),
.Y(n_7732)
);

INVx4_ASAP7_75t_L g7733 ( 
.A(n_7488),
.Y(n_7733)
);

AND2x2_ASAP7_75t_L g7734 ( 
.A(n_7414),
.B(n_7486),
.Y(n_7734)
);

INVx4_ASAP7_75t_L g7735 ( 
.A(n_7562),
.Y(n_7735)
);

AOI21xp5_ASAP7_75t_L g7736 ( 
.A1(n_7446),
.A2(n_295),
.B(n_296),
.Y(n_7736)
);

BUFx2_ASAP7_75t_L g7737 ( 
.A(n_7388),
.Y(n_7737)
);

A2O1A1Ixp33_ASAP7_75t_L g7738 ( 
.A1(n_7538),
.A2(n_298),
.B(n_295),
.C(n_297),
.Y(n_7738)
);

O2A1O1Ixp33_ASAP7_75t_L g7739 ( 
.A1(n_7588),
.A2(n_298),
.B(n_295),
.C(n_297),
.Y(n_7739)
);

CKINVDCx5p33_ASAP7_75t_R g7740 ( 
.A(n_7595),
.Y(n_7740)
);

INVx1_ASAP7_75t_L g7741 ( 
.A(n_7450),
.Y(n_7741)
);

INVx2_ASAP7_75t_L g7742 ( 
.A(n_7461),
.Y(n_7742)
);

A2O1A1Ixp33_ASAP7_75t_SL g7743 ( 
.A1(n_7570),
.A2(n_301),
.B(n_299),
.C(n_300),
.Y(n_7743)
);

AOI221xp5_ASAP7_75t_L g7744 ( 
.A1(n_7448),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.C(n_302),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7452),
.Y(n_7745)
);

OR2x2_ASAP7_75t_L g7746 ( 
.A(n_7524),
.B(n_299),
.Y(n_7746)
);

NOR2xp33_ASAP7_75t_L g7747 ( 
.A(n_7502),
.B(n_300),
.Y(n_7747)
);

INVx2_ASAP7_75t_SL g7748 ( 
.A(n_7587),
.Y(n_7748)
);

O2A1O1Ixp33_ASAP7_75t_SL g7749 ( 
.A1(n_7600),
.A2(n_303),
.B(n_301),
.C(n_302),
.Y(n_7749)
);

NOR2x1_ASAP7_75t_SL g7750 ( 
.A(n_7465),
.B(n_302),
.Y(n_7750)
);

BUFx4f_ASAP7_75t_SL g7751 ( 
.A(n_7579),
.Y(n_7751)
);

AND2x2_ASAP7_75t_L g7752 ( 
.A(n_7459),
.B(n_303),
.Y(n_7752)
);

NAND3xp33_ASAP7_75t_L g7753 ( 
.A(n_7448),
.B(n_304),
.C(n_305),
.Y(n_7753)
);

OR2x2_ASAP7_75t_L g7754 ( 
.A(n_7589),
.B(n_304),
.Y(n_7754)
);

AND2x2_ASAP7_75t_L g7755 ( 
.A(n_7485),
.B(n_7562),
.Y(n_7755)
);

NOR2xp33_ASAP7_75t_L g7756 ( 
.A(n_7508),
.B(n_304),
.Y(n_7756)
);

AND2x2_ASAP7_75t_L g7757 ( 
.A(n_7599),
.B(n_305),
.Y(n_7757)
);

AND2x2_ASAP7_75t_SL g7758 ( 
.A(n_7463),
.B(n_305),
.Y(n_7758)
);

AND2x2_ASAP7_75t_L g7759 ( 
.A(n_7601),
.B(n_306),
.Y(n_7759)
);

INVxp67_ASAP7_75t_L g7760 ( 
.A(n_7603),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7460),
.Y(n_7761)
);

INVx4_ASAP7_75t_L g7762 ( 
.A(n_7603),
.Y(n_7762)
);

NAND2xp33_ASAP7_75t_R g7763 ( 
.A(n_7381),
.B(n_306),
.Y(n_7763)
);

AOI221xp5_ASAP7_75t_L g7764 ( 
.A1(n_7441),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.C(n_310),
.Y(n_7764)
);

OAI21x1_ASAP7_75t_SL g7765 ( 
.A1(n_7387),
.A2(n_308),
.B(n_309),
.Y(n_7765)
);

AND2x2_ASAP7_75t_L g7766 ( 
.A(n_7382),
.B(n_309),
.Y(n_7766)
);

O2A1O1Ixp33_ASAP7_75t_SL g7767 ( 
.A1(n_7475),
.A2(n_7500),
.B(n_7387),
.C(n_7588),
.Y(n_7767)
);

AND2x2_ASAP7_75t_L g7768 ( 
.A(n_7592),
.B(n_7543),
.Y(n_7768)
);

AOI221xp5_ASAP7_75t_L g7769 ( 
.A1(n_7573),
.A2(n_7537),
.B1(n_7536),
.B2(n_7533),
.C(n_7606),
.Y(n_7769)
);

OR2x6_ASAP7_75t_L g7770 ( 
.A(n_7581),
.B(n_310),
.Y(n_7770)
);

OR2x2_ASAP7_75t_L g7771 ( 
.A(n_7556),
.B(n_310),
.Y(n_7771)
);

OR2x2_ASAP7_75t_L g7772 ( 
.A(n_7482),
.B(n_311),
.Y(n_7772)
);

NOR2xp33_ASAP7_75t_L g7773 ( 
.A(n_7508),
.B(n_311),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_7396),
.Y(n_7774)
);

AND2x2_ASAP7_75t_L g7775 ( 
.A(n_7615),
.B(n_7546),
.Y(n_7775)
);

AOI22xp5_ASAP7_75t_L g7776 ( 
.A1(n_7574),
.A2(n_2959),
.B1(n_2985),
.B2(n_2895),
.Y(n_7776)
);

INVx3_ASAP7_75t_L g7777 ( 
.A(n_7550),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7557),
.Y(n_7778)
);

AND2x2_ASAP7_75t_L g7779 ( 
.A(n_7615),
.B(n_311),
.Y(n_7779)
);

INVx1_ASAP7_75t_L g7780 ( 
.A(n_7558),
.Y(n_7780)
);

AND2x2_ASAP7_75t_L g7781 ( 
.A(n_7528),
.B(n_312),
.Y(n_7781)
);

AND2x2_ASAP7_75t_L g7782 ( 
.A(n_7613),
.B(n_312),
.Y(n_7782)
);

NOR2xp33_ASAP7_75t_R g7783 ( 
.A(n_7598),
.B(n_312),
.Y(n_7783)
);

AND2x2_ASAP7_75t_L g7784 ( 
.A(n_7613),
.B(n_313),
.Y(n_7784)
);

NAND2xp5_ASAP7_75t_L g7785 ( 
.A(n_7572),
.B(n_314),
.Y(n_7785)
);

AND2x2_ASAP7_75t_L g7786 ( 
.A(n_7535),
.B(n_314),
.Y(n_7786)
);

AO21x1_ASAP7_75t_L g7787 ( 
.A1(n_7426),
.A2(n_314),
.B(n_315),
.Y(n_7787)
);

O2A1O1Ixp33_ASAP7_75t_L g7788 ( 
.A1(n_7547),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_7788)
);

NAND3xp33_ASAP7_75t_L g7789 ( 
.A(n_7426),
.B(n_7518),
.C(n_7500),
.Y(n_7789)
);

AOI22xp5_ASAP7_75t_L g7790 ( 
.A1(n_7539),
.A2(n_3029),
.B1(n_2985),
.B2(n_1766),
.Y(n_7790)
);

A2O1A1Ixp33_ASAP7_75t_L g7791 ( 
.A1(n_7517),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_7791)
);

AND2x4_ASAP7_75t_L g7792 ( 
.A(n_7490),
.B(n_318),
.Y(n_7792)
);

INVx1_ASAP7_75t_L g7793 ( 
.A(n_7567),
.Y(n_7793)
);

AND2x4_ASAP7_75t_L g7794 ( 
.A(n_7491),
.B(n_318),
.Y(n_7794)
);

BUFx12f_ASAP7_75t_L g7795 ( 
.A(n_7603),
.Y(n_7795)
);

NAND2xp5_ASAP7_75t_L g7796 ( 
.A(n_7575),
.B(n_319),
.Y(n_7796)
);

INVx1_ASAP7_75t_L g7797 ( 
.A(n_7388),
.Y(n_7797)
);

HB1xp67_ASAP7_75t_L g7798 ( 
.A(n_7610),
.Y(n_7798)
);

INVx2_ASAP7_75t_L g7799 ( 
.A(n_7413),
.Y(n_7799)
);

A2O1A1Ixp33_ASAP7_75t_L g7800 ( 
.A1(n_7520),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_7800)
);

AND2x2_ASAP7_75t_L g7801 ( 
.A(n_7464),
.B(n_319),
.Y(n_7801)
);

OR2x2_ASAP7_75t_L g7802 ( 
.A(n_7482),
.B(n_320),
.Y(n_7802)
);

A2O1A1Ixp33_ASAP7_75t_L g7803 ( 
.A1(n_7581),
.A2(n_322),
.B(n_320),
.C(n_321),
.Y(n_7803)
);

AO21x2_ASAP7_75t_L g7804 ( 
.A1(n_7696),
.A2(n_7392),
.B(n_7529),
.Y(n_7804)
);

INVx2_ASAP7_75t_L g7805 ( 
.A(n_7637),
.Y(n_7805)
);

OR2x2_ASAP7_75t_L g7806 ( 
.A(n_7647),
.B(n_7451),
.Y(n_7806)
);

HB1xp67_ASAP7_75t_L g7807 ( 
.A(n_7724),
.Y(n_7807)
);

INVx2_ASAP7_75t_L g7808 ( 
.A(n_7692),
.Y(n_7808)
);

AND2x2_ASAP7_75t_L g7809 ( 
.A(n_7621),
.B(n_7464),
.Y(n_7809)
);

INVx1_ASAP7_75t_L g7810 ( 
.A(n_7724),
.Y(n_7810)
);

AND2x4_ASAP7_75t_L g7811 ( 
.A(n_7656),
.B(n_7576),
.Y(n_7811)
);

BUFx2_ASAP7_75t_L g7812 ( 
.A(n_7686),
.Y(n_7812)
);

INVx1_ASAP7_75t_L g7813 ( 
.A(n_7713),
.Y(n_7813)
);

INVx2_ASAP7_75t_L g7814 ( 
.A(n_7692),
.Y(n_7814)
);

AND2x2_ASAP7_75t_L g7815 ( 
.A(n_7690),
.B(n_7385),
.Y(n_7815)
);

AND2x2_ASAP7_75t_L g7816 ( 
.A(n_7620),
.B(n_7394),
.Y(n_7816)
);

INVx2_ASAP7_75t_L g7817 ( 
.A(n_7640),
.Y(n_7817)
);

OR2x2_ASAP7_75t_L g7818 ( 
.A(n_7772),
.B(n_7451),
.Y(n_7818)
);

INVx2_ASAP7_75t_L g7819 ( 
.A(n_7715),
.Y(n_7819)
);

NAND2xp5_ASAP7_75t_L g7820 ( 
.A(n_7713),
.B(n_7392),
.Y(n_7820)
);

NAND2xp5_ASAP7_75t_L g7821 ( 
.A(n_7719),
.B(n_7659),
.Y(n_7821)
);

NOR2xp33_ASAP7_75t_L g7822 ( 
.A(n_7646),
.B(n_7582),
.Y(n_7822)
);

OAI31xp33_ASAP7_75t_SL g7823 ( 
.A1(n_7688),
.A2(n_7609),
.A3(n_7515),
.B(n_7395),
.Y(n_7823)
);

OR2x2_ASAP7_75t_L g7824 ( 
.A(n_7802),
.B(n_7649),
.Y(n_7824)
);

AOI221xp5_ASAP7_75t_L g7825 ( 
.A1(n_7623),
.A2(n_7767),
.B1(n_7627),
.B2(n_7630),
.C(n_7789),
.Y(n_7825)
);

CKINVDCx20_ASAP7_75t_R g7826 ( 
.A(n_7751),
.Y(n_7826)
);

INVx1_ASAP7_75t_L g7827 ( 
.A(n_7719),
.Y(n_7827)
);

AND2x2_ASAP7_75t_L g7828 ( 
.A(n_7673),
.B(n_7596),
.Y(n_7828)
);

INVx2_ASAP7_75t_L g7829 ( 
.A(n_7698),
.Y(n_7829)
);

OAI31xp33_ASAP7_75t_L g7830 ( 
.A1(n_7753),
.A2(n_7445),
.A3(n_7518),
.B(n_7544),
.Y(n_7830)
);

NAND2xp5_ASAP7_75t_L g7831 ( 
.A(n_7694),
.B(n_7421),
.Y(n_7831)
);

INVxp67_ASAP7_75t_SL g7832 ( 
.A(n_7787),
.Y(n_7832)
);

INVx2_ASAP7_75t_L g7833 ( 
.A(n_7698),
.Y(n_7833)
);

INVx1_ASAP7_75t_L g7834 ( 
.A(n_7679),
.Y(n_7834)
);

CKINVDCx20_ASAP7_75t_R g7835 ( 
.A(n_7722),
.Y(n_7835)
);

BUFx2_ASAP7_75t_L g7836 ( 
.A(n_7624),
.Y(n_7836)
);

INVx2_ASAP7_75t_L g7837 ( 
.A(n_7715),
.Y(n_7837)
);

INVx1_ASAP7_75t_L g7838 ( 
.A(n_7746),
.Y(n_7838)
);

INVx2_ASAP7_75t_L g7839 ( 
.A(n_7758),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7737),
.Y(n_7840)
);

AND2x2_ASAP7_75t_L g7841 ( 
.A(n_7654),
.B(n_7596),
.Y(n_7841)
);

INVx1_ASAP7_75t_L g7842 ( 
.A(n_7737),
.Y(n_7842)
);

INVx1_ASAP7_75t_L g7843 ( 
.A(n_7689),
.Y(n_7843)
);

INVx1_ASAP7_75t_L g7844 ( 
.A(n_7703),
.Y(n_7844)
);

INVx2_ASAP7_75t_SL g7845 ( 
.A(n_7631),
.Y(n_7845)
);

BUFx6f_ASAP7_75t_L g7846 ( 
.A(n_7675),
.Y(n_7846)
);

INVx2_ASAP7_75t_SL g7847 ( 
.A(n_7634),
.Y(n_7847)
);

AND2x2_ASAP7_75t_L g7848 ( 
.A(n_7755),
.B(n_7472),
.Y(n_7848)
);

BUFx4f_ASAP7_75t_L g7849 ( 
.A(n_7693),
.Y(n_7849)
);

HB1xp67_ASAP7_75t_L g7850 ( 
.A(n_7710),
.Y(n_7850)
);

INVxp67_ASAP7_75t_SL g7851 ( 
.A(n_7671),
.Y(n_7851)
);

AND2x2_ASAP7_75t_L g7852 ( 
.A(n_7752),
.B(n_7472),
.Y(n_7852)
);

INVx2_ASAP7_75t_L g7853 ( 
.A(n_7750),
.Y(n_7853)
);

AO31x2_ASAP7_75t_L g7854 ( 
.A1(n_7704),
.A2(n_7531),
.A3(n_7569),
.B(n_7561),
.Y(n_7854)
);

AND2x2_ASAP7_75t_L g7855 ( 
.A(n_7712),
.B(n_7781),
.Y(n_7855)
);

OR2x2_ASAP7_75t_L g7856 ( 
.A(n_7651),
.B(n_7610),
.Y(n_7856)
);

INVx2_ASAP7_75t_L g7857 ( 
.A(n_7718),
.Y(n_7857)
);

INVxp67_ASAP7_75t_SL g7858 ( 
.A(n_7701),
.Y(n_7858)
);

INVx2_ASAP7_75t_L g7859 ( 
.A(n_7718),
.Y(n_7859)
);

HB1xp67_ASAP7_75t_L g7860 ( 
.A(n_7643),
.Y(n_7860)
);

INVx2_ASAP7_75t_L g7861 ( 
.A(n_7691),
.Y(n_7861)
);

NAND2xp5_ASAP7_75t_L g7862 ( 
.A(n_7685),
.B(n_7421),
.Y(n_7862)
);

INVx2_ASAP7_75t_L g7863 ( 
.A(n_7691),
.Y(n_7863)
);

HB1xp67_ASAP7_75t_L g7864 ( 
.A(n_7639),
.Y(n_7864)
);

INVx2_ASAP7_75t_L g7865 ( 
.A(n_7795),
.Y(n_7865)
);

INVx1_ASAP7_75t_L g7866 ( 
.A(n_7717),
.Y(n_7866)
);

INVx1_ASAP7_75t_L g7867 ( 
.A(n_7732),
.Y(n_7867)
);

AND2x2_ASAP7_75t_L g7868 ( 
.A(n_7666),
.B(n_7550),
.Y(n_7868)
);

INVx2_ASAP7_75t_L g7869 ( 
.A(n_7792),
.Y(n_7869)
);

INVx2_ASAP7_75t_L g7870 ( 
.A(n_7792),
.Y(n_7870)
);

AND2x2_ASAP7_75t_L g7871 ( 
.A(n_7616),
.B(n_7559),
.Y(n_7871)
);

INVx2_ASAP7_75t_L g7872 ( 
.A(n_7794),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_7741),
.Y(n_7873)
);

INVx1_ASAP7_75t_L g7874 ( 
.A(n_7745),
.Y(n_7874)
);

INVxp67_ASAP7_75t_R g7875 ( 
.A(n_7681),
.Y(n_7875)
);

AOI22xp33_ASAP7_75t_SL g7876 ( 
.A1(n_7635),
.A2(n_7632),
.B1(n_7617),
.B2(n_7633),
.Y(n_7876)
);

INVx1_ASAP7_75t_L g7877 ( 
.A(n_7761),
.Y(n_7877)
);

INVx2_ASAP7_75t_L g7878 ( 
.A(n_7794),
.Y(n_7878)
);

INVx1_ASAP7_75t_L g7879 ( 
.A(n_7771),
.Y(n_7879)
);

OR2x2_ASAP7_75t_L g7880 ( 
.A(n_7785),
.B(n_7610),
.Y(n_7880)
);

INVxp67_ASAP7_75t_L g7881 ( 
.A(n_7644),
.Y(n_7881)
);

INVx1_ASAP7_75t_L g7882 ( 
.A(n_7730),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_7731),
.Y(n_7883)
);

INVxp67_ASAP7_75t_L g7884 ( 
.A(n_7756),
.Y(n_7884)
);

INVx3_ASAP7_75t_L g7885 ( 
.A(n_7733),
.Y(n_7885)
);

AND2x2_ASAP7_75t_L g7886 ( 
.A(n_7667),
.B(n_7559),
.Y(n_7886)
);

INVx2_ASAP7_75t_L g7887 ( 
.A(n_7678),
.Y(n_7887)
);

INVx3_ASAP7_75t_L g7888 ( 
.A(n_7678),
.Y(n_7888)
);

OR2x2_ASAP7_75t_L g7889 ( 
.A(n_7748),
.B(n_7433),
.Y(n_7889)
);

OR2x2_ASAP7_75t_L g7890 ( 
.A(n_7796),
.B(n_7555),
.Y(n_7890)
);

INVx1_ASAP7_75t_L g7891 ( 
.A(n_7699),
.Y(n_7891)
);

INVx1_ASAP7_75t_L g7892 ( 
.A(n_7725),
.Y(n_7892)
);

INVx2_ASAP7_75t_L g7893 ( 
.A(n_7720),
.Y(n_7893)
);

BUFx2_ASAP7_75t_L g7894 ( 
.A(n_7721),
.Y(n_7894)
);

INVx3_ASAP7_75t_L g7895 ( 
.A(n_7720),
.Y(n_7895)
);

INVx1_ASAP7_75t_L g7896 ( 
.A(n_7754),
.Y(n_7896)
);

AND2x2_ASAP7_75t_L g7897 ( 
.A(n_7667),
.B(n_7548),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_7622),
.Y(n_7898)
);

INVx1_ASAP7_75t_L g7899 ( 
.A(n_7625),
.Y(n_7899)
);

AND2x2_ASAP7_75t_L g7900 ( 
.A(n_7734),
.B(n_7548),
.Y(n_7900)
);

AND2x4_ASAP7_75t_L g7901 ( 
.A(n_7638),
.B(n_7418),
.Y(n_7901)
);

OR2x2_ASAP7_75t_L g7902 ( 
.A(n_7702),
.B(n_7593),
.Y(n_7902)
);

INVx2_ASAP7_75t_L g7903 ( 
.A(n_7762),
.Y(n_7903)
);

INVxp67_ASAP7_75t_L g7904 ( 
.A(n_7773),
.Y(n_7904)
);

INVx2_ASAP7_75t_L g7905 ( 
.A(n_7697),
.Y(n_7905)
);

AO21x1_ASAP7_75t_SL g7906 ( 
.A1(n_7628),
.A2(n_7560),
.B(n_7474),
.Y(n_7906)
);

INVx2_ASAP7_75t_L g7907 ( 
.A(n_7698),
.Y(n_7907)
);

INVx1_ASAP7_75t_L g7908 ( 
.A(n_7797),
.Y(n_7908)
);

AND2x2_ASAP7_75t_L g7909 ( 
.A(n_7618),
.B(n_7470),
.Y(n_7909)
);

AOI33xp33_ASAP7_75t_L g7910 ( 
.A1(n_7619),
.A2(n_7551),
.A3(n_7552),
.B1(n_7553),
.B2(n_7549),
.B3(n_7509),
.Y(n_7910)
);

AND2x2_ASAP7_75t_L g7911 ( 
.A(n_7618),
.B(n_7478),
.Y(n_7911)
);

AND2x2_ASAP7_75t_L g7912 ( 
.A(n_7775),
.B(n_7480),
.Y(n_7912)
);

OR2x2_ASAP7_75t_L g7913 ( 
.A(n_7702),
.B(n_7593),
.Y(n_7913)
);

INVx1_ASAP7_75t_L g7914 ( 
.A(n_7636),
.Y(n_7914)
);

NOR2xp33_ASAP7_75t_L g7915 ( 
.A(n_7740),
.B(n_7534),
.Y(n_7915)
);

BUFx2_ASAP7_75t_L g7916 ( 
.A(n_7677),
.Y(n_7916)
);

OR2x2_ASAP7_75t_L g7917 ( 
.A(n_7684),
.B(n_7483),
.Y(n_7917)
);

INVx2_ASAP7_75t_L g7918 ( 
.A(n_7735),
.Y(n_7918)
);

INVx2_ASAP7_75t_L g7919 ( 
.A(n_7728),
.Y(n_7919)
);

INVx2_ASAP7_75t_L g7920 ( 
.A(n_7777),
.Y(n_7920)
);

INVx1_ASAP7_75t_L g7921 ( 
.A(n_7798),
.Y(n_7921)
);

INVx1_ASAP7_75t_L g7922 ( 
.A(n_7757),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_7759),
.Y(n_7923)
);

AND2x4_ASAP7_75t_SL g7924 ( 
.A(n_7726),
.B(n_7381),
.Y(n_7924)
);

INVx2_ASAP7_75t_L g7925 ( 
.A(n_7663),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_7723),
.Y(n_7926)
);

AND2x2_ASAP7_75t_L g7927 ( 
.A(n_7626),
.B(n_7484),
.Y(n_7927)
);

AND2x2_ASAP7_75t_L g7928 ( 
.A(n_7658),
.B(n_7801),
.Y(n_7928)
);

INVx2_ASAP7_75t_L g7929 ( 
.A(n_7729),
.Y(n_7929)
);

AOI21xp5_ASAP7_75t_L g7930 ( 
.A1(n_7707),
.A2(n_7539),
.B(n_7425),
.Y(n_7930)
);

INVx1_ASAP7_75t_L g7931 ( 
.A(n_7700),
.Y(n_7931)
);

BUFx3_ASAP7_75t_L g7932 ( 
.A(n_7669),
.Y(n_7932)
);

AND2x4_ASAP7_75t_L g7933 ( 
.A(n_7709),
.B(n_7510),
.Y(n_7933)
);

AND2x2_ASAP7_75t_L g7934 ( 
.A(n_7653),
.B(n_7492),
.Y(n_7934)
);

INVx2_ASAP7_75t_L g7935 ( 
.A(n_7633),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_7687),
.Y(n_7936)
);

AND2x2_ASAP7_75t_L g7937 ( 
.A(n_7768),
.B(n_7705),
.Y(n_7937)
);

INVx2_ASAP7_75t_SL g7938 ( 
.A(n_7672),
.Y(n_7938)
);

INVx2_ASAP7_75t_L g7939 ( 
.A(n_7765),
.Y(n_7939)
);

AND2x2_ASAP7_75t_L g7940 ( 
.A(n_7706),
.B(n_7495),
.Y(n_7940)
);

INVx1_ASAP7_75t_L g7941 ( 
.A(n_7778),
.Y(n_7941)
);

INVx1_ASAP7_75t_L g7942 ( 
.A(n_7780),
.Y(n_7942)
);

INVx1_ASAP7_75t_L g7943 ( 
.A(n_7793),
.Y(n_7943)
);

INVx4_ASAP7_75t_L g7944 ( 
.A(n_7680),
.Y(n_7944)
);

INVx2_ASAP7_75t_SL g7945 ( 
.A(n_7782),
.Y(n_7945)
);

OR2x2_ASAP7_75t_L g7946 ( 
.A(n_7774),
.B(n_7498),
.Y(n_7946)
);

INVx1_ASAP7_75t_L g7947 ( 
.A(n_7642),
.Y(n_7947)
);

INVx1_ASAP7_75t_L g7948 ( 
.A(n_7648),
.Y(n_7948)
);

INVx4_ASAP7_75t_L g7949 ( 
.A(n_7668),
.Y(n_7949)
);

INVx2_ASAP7_75t_L g7950 ( 
.A(n_7633),
.Y(n_7950)
);

INVx2_ASAP7_75t_L g7951 ( 
.A(n_7784),
.Y(n_7951)
);

OAI21xp33_ASAP7_75t_L g7952 ( 
.A1(n_7876),
.A2(n_7652),
.B(n_7650),
.Y(n_7952)
);

AOI22xp5_ASAP7_75t_L g7953 ( 
.A1(n_7935),
.A2(n_7950),
.B1(n_7876),
.B2(n_7832),
.Y(n_7953)
);

AND2x2_ASAP7_75t_L g7954 ( 
.A(n_7812),
.B(n_7766),
.Y(n_7954)
);

NAND2xp5_ASAP7_75t_L g7955 ( 
.A(n_7832),
.B(n_7894),
.Y(n_7955)
);

AND2x2_ASAP7_75t_L g7956 ( 
.A(n_7875),
.B(n_7836),
.Y(n_7956)
);

OAI21xp5_ASAP7_75t_L g7957 ( 
.A1(n_7930),
.A2(n_7736),
.B(n_7660),
.Y(n_7957)
);

NAND2xp5_ASAP7_75t_L g7958 ( 
.A(n_7916),
.B(n_7657),
.Y(n_7958)
);

NOR3xp33_ASAP7_75t_L g7959 ( 
.A(n_7825),
.B(n_7769),
.C(n_7744),
.Y(n_7959)
);

NAND2xp5_ASAP7_75t_L g7960 ( 
.A(n_7938),
.B(n_7674),
.Y(n_7960)
);

AND2x2_ASAP7_75t_L g7961 ( 
.A(n_7855),
.B(n_7779),
.Y(n_7961)
);

NAND2xp5_ASAP7_75t_L g7962 ( 
.A(n_7945),
.B(n_7786),
.Y(n_7962)
);

AND2x2_ASAP7_75t_L g7963 ( 
.A(n_7928),
.B(n_7881),
.Y(n_7963)
);

NOR2xp33_ASAP7_75t_L g7964 ( 
.A(n_7826),
.B(n_7835),
.Y(n_7964)
);

OAI221xp5_ASAP7_75t_L g7965 ( 
.A1(n_7935),
.A2(n_7645),
.B1(n_7763),
.B2(n_7617),
.C(n_7641),
.Y(n_7965)
);

AOI21xp33_ASAP7_75t_SL g7966 ( 
.A1(n_7950),
.A2(n_7661),
.B(n_7639),
.Y(n_7966)
);

AOI22xp33_ASAP7_75t_SL g7967 ( 
.A1(n_7829),
.A2(n_7629),
.B1(n_7442),
.B2(n_7534),
.Y(n_7967)
);

AND2x2_ASAP7_75t_L g7968 ( 
.A(n_7881),
.B(n_7676),
.Y(n_7968)
);

AOI22xp33_ASAP7_75t_L g7969 ( 
.A1(n_7829),
.A2(n_7568),
.B1(n_7442),
.B2(n_7507),
.Y(n_7969)
);

NOR3xp33_ASAP7_75t_L g7970 ( 
.A(n_7825),
.B(n_7760),
.C(n_7727),
.Y(n_7970)
);

NOR2xp33_ASAP7_75t_R g7971 ( 
.A(n_7826),
.B(n_7665),
.Y(n_7971)
);

AND2x2_ASAP7_75t_L g7972 ( 
.A(n_7871),
.B(n_7683),
.Y(n_7972)
);

OAI21xp5_ASAP7_75t_SL g7973 ( 
.A1(n_7823),
.A2(n_7739),
.B(n_7655),
.Y(n_7973)
);

NAND3xp33_ASAP7_75t_L g7974 ( 
.A(n_7833),
.B(n_7716),
.C(n_7670),
.Y(n_7974)
);

NAND2xp5_ASAP7_75t_L g7975 ( 
.A(n_7940),
.B(n_7749),
.Y(n_7975)
);

NAND4xp25_ASAP7_75t_L g7976 ( 
.A(n_7823),
.B(n_7682),
.C(n_7743),
.D(n_7711),
.Y(n_7976)
);

NAND4xp25_ASAP7_75t_SL g7977 ( 
.A(n_7910),
.B(n_7764),
.C(n_7738),
.D(n_7788),
.Y(n_7977)
);

AOI22xp33_ASAP7_75t_L g7978 ( 
.A1(n_7833),
.A2(n_7568),
.B1(n_7662),
.B2(n_7466),
.Y(n_7978)
);

NAND2xp5_ASAP7_75t_L g7979 ( 
.A(n_7937),
.B(n_7747),
.Y(n_7979)
);

INVx1_ASAP7_75t_L g7980 ( 
.A(n_7807),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_L g7981 ( 
.A(n_7926),
.B(n_7791),
.Y(n_7981)
);

OAI21xp5_ASAP7_75t_SL g7982 ( 
.A1(n_7930),
.A2(n_7790),
.B(n_7560),
.Y(n_7982)
);

OA21x2_ASAP7_75t_L g7983 ( 
.A1(n_7907),
.A2(n_7545),
.B(n_7419),
.Y(n_7983)
);

NAND3xp33_ASAP7_75t_L g7984 ( 
.A(n_7907),
.B(n_7800),
.C(n_7714),
.Y(n_7984)
);

NAND2xp5_ASAP7_75t_L g7985 ( 
.A(n_7860),
.B(n_7742),
.Y(n_7985)
);

OAI21xp5_ASAP7_75t_L g7986 ( 
.A1(n_7821),
.A2(n_7585),
.B(n_7803),
.Y(n_7986)
);

NAND2xp5_ASAP7_75t_L g7987 ( 
.A(n_7860),
.B(n_7770),
.Y(n_7987)
);

NAND4xp25_ASAP7_75t_L g7988 ( 
.A(n_7897),
.B(n_7604),
.C(n_7436),
.D(n_7504),
.Y(n_7988)
);

NOR3xp33_ASAP7_75t_L g7989 ( 
.A(n_7865),
.B(n_7695),
.C(n_7664),
.Y(n_7989)
);

NAND2xp5_ASAP7_75t_SL g7990 ( 
.A(n_7849),
.B(n_7510),
.Y(n_7990)
);

OAI21xp33_ASAP7_75t_SL g7991 ( 
.A1(n_7821),
.A2(n_7407),
.B(n_7402),
.Y(n_7991)
);

NAND2xp5_ASAP7_75t_L g7992 ( 
.A(n_7949),
.B(n_7770),
.Y(n_7992)
);

NOR2xp33_ASAP7_75t_L g7993 ( 
.A(n_7835),
.B(n_7799),
.Y(n_7993)
);

NAND2xp5_ASAP7_75t_L g7994 ( 
.A(n_7949),
.B(n_7846),
.Y(n_7994)
);

OAI21xp5_ASAP7_75t_SL g7995 ( 
.A1(n_7807),
.A2(n_7586),
.B(n_7512),
.Y(n_7995)
);

NAND2xp5_ASAP7_75t_L g7996 ( 
.A(n_7846),
.B(n_7783),
.Y(n_7996)
);

AOI22xp5_ASAP7_75t_L g7997 ( 
.A1(n_7915),
.A2(n_7566),
.B1(n_7425),
.B2(n_7381),
.Y(n_7997)
);

OAI221xp5_ASAP7_75t_SL g7998 ( 
.A1(n_7910),
.A2(n_7425),
.B1(n_7586),
.B2(n_7563),
.C(n_7487),
.Y(n_7998)
);

NAND2xp5_ASAP7_75t_L g7999 ( 
.A(n_7846),
.B(n_7457),
.Y(n_7999)
);

AOI21xp33_ASAP7_75t_L g8000 ( 
.A1(n_7862),
.A2(n_7477),
.B(n_7469),
.Y(n_8000)
);

NAND2xp5_ASAP7_75t_L g8001 ( 
.A(n_7888),
.B(n_7457),
.Y(n_8001)
);

NAND3xp33_ASAP7_75t_L g8002 ( 
.A(n_7810),
.B(n_7406),
.C(n_7708),
.Y(n_8002)
);

AND2x2_ASAP7_75t_SL g8003 ( 
.A(n_7924),
.B(n_7393),
.Y(n_8003)
);

NAND2xp5_ASAP7_75t_L g8004 ( 
.A(n_7888),
.B(n_7895),
.Y(n_8004)
);

NOR2xp33_ASAP7_75t_L g8005 ( 
.A(n_7944),
.B(n_7566),
.Y(n_8005)
);

INVx1_ASAP7_75t_L g8006 ( 
.A(n_7850),
.Y(n_8006)
);

AND2x2_ASAP7_75t_L g8007 ( 
.A(n_7841),
.B(n_7499),
.Y(n_8007)
);

AND2x2_ASAP7_75t_L g8008 ( 
.A(n_7848),
.B(n_7868),
.Y(n_8008)
);

AND2x2_ASAP7_75t_L g8009 ( 
.A(n_7886),
.B(n_7514),
.Y(n_8009)
);

AND2x2_ASAP7_75t_L g8010 ( 
.A(n_7927),
.B(n_7516),
.Y(n_8010)
);

OAI221xp5_ASAP7_75t_L g8011 ( 
.A1(n_7830),
.A2(n_7915),
.B1(n_7862),
.B2(n_7831),
.C(n_7850),
.Y(n_8011)
);

AOI32xp33_ASAP7_75t_L g8012 ( 
.A1(n_7858),
.A2(n_7541),
.A3(n_7389),
.B1(n_7383),
.B2(n_7462),
.Y(n_8012)
);

NAND2xp5_ASAP7_75t_L g8013 ( 
.A(n_7895),
.B(n_7776),
.Y(n_8013)
);

NAND3xp33_ASAP7_75t_L g8014 ( 
.A(n_7830),
.B(n_7406),
.C(n_7494),
.Y(n_8014)
);

AND2x2_ASAP7_75t_L g8015 ( 
.A(n_7828),
.B(n_7519),
.Y(n_8015)
);

AND2x2_ASAP7_75t_SL g8016 ( 
.A(n_7924),
.B(n_7494),
.Y(n_8016)
);

NAND2xp5_ASAP7_75t_L g8017 ( 
.A(n_7922),
.B(n_7467),
.Y(n_8017)
);

NAND2xp5_ASAP7_75t_L g8018 ( 
.A(n_7923),
.B(n_7467),
.Y(n_8018)
);

NAND2xp5_ASAP7_75t_L g8019 ( 
.A(n_7932),
.B(n_7522),
.Y(n_8019)
);

AND2x2_ASAP7_75t_L g8020 ( 
.A(n_7809),
.B(n_7530),
.Y(n_8020)
);

NAND2xp5_ASAP7_75t_L g8021 ( 
.A(n_7932),
.B(n_7431),
.Y(n_8021)
);

OAI21xp33_ASAP7_75t_L g8022 ( 
.A1(n_7822),
.A2(n_7815),
.B(n_7903),
.Y(n_8022)
);

NAND2xp33_ASAP7_75t_SL g8023 ( 
.A(n_7806),
.B(n_7565),
.Y(n_8023)
);

AND2x2_ASAP7_75t_L g8024 ( 
.A(n_7811),
.B(n_7431),
.Y(n_8024)
);

NAND2xp5_ASAP7_75t_L g8025 ( 
.A(n_7951),
.B(n_7405),
.Y(n_8025)
);

AND2x2_ASAP7_75t_L g8026 ( 
.A(n_7811),
.B(n_7505),
.Y(n_8026)
);

NOR3xp33_ASAP7_75t_SL g8027 ( 
.A(n_7822),
.B(n_7405),
.C(n_7505),
.Y(n_8027)
);

AOI21xp5_ASAP7_75t_SL g8028 ( 
.A1(n_7820),
.A2(n_7473),
.B(n_322),
.Y(n_8028)
);

NAND3xp33_ASAP7_75t_L g8029 ( 
.A(n_7864),
.B(n_7473),
.C(n_7506),
.Y(n_8029)
);

AND2x2_ASAP7_75t_L g8030 ( 
.A(n_7944),
.B(n_7506),
.Y(n_8030)
);

NAND2xp5_ASAP7_75t_SL g8031 ( 
.A(n_7849),
.B(n_7506),
.Y(n_8031)
);

HB1xp67_ASAP7_75t_L g8032 ( 
.A(n_7864),
.Y(n_8032)
);

OAI22xp5_ASAP7_75t_L g8033 ( 
.A1(n_7858),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_8033)
);

OAI221xp5_ASAP7_75t_L g8034 ( 
.A1(n_7831),
.A2(n_7827),
.B1(n_7813),
.B2(n_7820),
.C(n_7856),
.Y(n_8034)
);

OAI22xp5_ASAP7_75t_L g8035 ( 
.A1(n_7853),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.Y(n_8035)
);

NAND2xp5_ASAP7_75t_L g8036 ( 
.A(n_7838),
.B(n_323),
.Y(n_8036)
);

NAND2xp5_ASAP7_75t_L g8037 ( 
.A(n_7936),
.B(n_324),
.Y(n_8037)
);

OAI22xp5_ASAP7_75t_L g8038 ( 
.A1(n_7925),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_8038)
);

NAND2xp5_ASAP7_75t_L g8039 ( 
.A(n_7879),
.B(n_326),
.Y(n_8039)
);

OAI21xp5_ASAP7_75t_L g8040 ( 
.A1(n_7884),
.A2(n_326),
.B(n_327),
.Y(n_8040)
);

NAND2xp33_ASAP7_75t_L g8041 ( 
.A(n_7817),
.B(n_327),
.Y(n_8041)
);

NAND2xp5_ASAP7_75t_L g8042 ( 
.A(n_7896),
.B(n_328),
.Y(n_8042)
);

NAND2xp5_ASAP7_75t_L g8043 ( 
.A(n_7905),
.B(n_328),
.Y(n_8043)
);

NAND2xp5_ASAP7_75t_L g8044 ( 
.A(n_7887),
.B(n_329),
.Y(n_8044)
);

NAND2xp5_ASAP7_75t_SL g8045 ( 
.A(n_7893),
.B(n_7852),
.Y(n_8045)
);

INVx1_ASAP7_75t_L g8046 ( 
.A(n_7921),
.Y(n_8046)
);

NAND4xp25_ASAP7_75t_L g8047 ( 
.A(n_7816),
.B(n_331),
.C(n_329),
.D(n_330),
.Y(n_8047)
);

NAND2xp5_ASAP7_75t_L g8048 ( 
.A(n_7929),
.B(n_7912),
.Y(n_8048)
);

OAI21xp5_ASAP7_75t_SL g8049 ( 
.A1(n_7900),
.A2(n_329),
.B(n_330),
.Y(n_8049)
);

NAND2xp5_ASAP7_75t_SL g8050 ( 
.A(n_7933),
.B(n_1751),
.Y(n_8050)
);

AOI22xp33_ASAP7_75t_L g8051 ( 
.A1(n_7839),
.A2(n_3029),
.B1(n_2985),
.B2(n_1781),
.Y(n_8051)
);

NAND3xp33_ASAP7_75t_L g8052 ( 
.A(n_7840),
.B(n_330),
.C(n_332),
.Y(n_8052)
);

OAI21xp5_ASAP7_75t_SL g8053 ( 
.A1(n_7933),
.A2(n_332),
.B(n_333),
.Y(n_8053)
);

NAND4xp25_ASAP7_75t_L g8054 ( 
.A(n_7805),
.B(n_334),
.C(n_332),
.D(n_333),
.Y(n_8054)
);

NAND2xp5_ASAP7_75t_L g8055 ( 
.A(n_7884),
.B(n_334),
.Y(n_8055)
);

AND2x2_ASAP7_75t_L g8056 ( 
.A(n_7845),
.B(n_7847),
.Y(n_8056)
);

NAND2xp5_ASAP7_75t_L g8057 ( 
.A(n_7904),
.B(n_334),
.Y(n_8057)
);

NAND2xp5_ASAP7_75t_L g8058 ( 
.A(n_7904),
.B(n_335),
.Y(n_8058)
);

OA21x2_ASAP7_75t_L g8059 ( 
.A1(n_7842),
.A2(n_7851),
.B(n_7844),
.Y(n_8059)
);

AOI22xp33_ASAP7_75t_L g8060 ( 
.A1(n_7834),
.A2(n_7931),
.B1(n_7851),
.B2(n_7880),
.Y(n_8060)
);

OAI21xp5_ASAP7_75t_SL g8061 ( 
.A1(n_7885),
.A2(n_335),
.B(n_336),
.Y(n_8061)
);

AND2x2_ASAP7_75t_L g8062 ( 
.A(n_7885),
.B(n_335),
.Y(n_8062)
);

AOI221xp5_ASAP7_75t_L g8063 ( 
.A1(n_7883),
.A2(n_7804),
.B1(n_7882),
.B2(n_7892),
.C(n_7891),
.Y(n_8063)
);

OAI22xp5_ASAP7_75t_L g8064 ( 
.A1(n_7808),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_8064)
);

NAND4xp25_ASAP7_75t_L g8065 ( 
.A(n_7918),
.B(n_339),
.C(n_337),
.D(n_338),
.Y(n_8065)
);

NAND3xp33_ASAP7_75t_L g8066 ( 
.A(n_7902),
.B(n_7913),
.C(n_7824),
.Y(n_8066)
);

NAND2xp5_ASAP7_75t_L g8067 ( 
.A(n_7901),
.B(n_339),
.Y(n_8067)
);

NAND2xp5_ASAP7_75t_L g8068 ( 
.A(n_7901),
.B(n_340),
.Y(n_8068)
);

NAND4xp25_ASAP7_75t_L g8069 ( 
.A(n_7919),
.B(n_340),
.C(n_341),
.D(n_413),
.Y(n_8069)
);

NAND2xp5_ASAP7_75t_L g8070 ( 
.A(n_7909),
.B(n_340),
.Y(n_8070)
);

NAND2xp5_ASAP7_75t_L g8071 ( 
.A(n_7911),
.B(n_7934),
.Y(n_8071)
);

NAND3xp33_ASAP7_75t_L g8072 ( 
.A(n_7814),
.B(n_341),
.C(n_414),
.Y(n_8072)
);

AND2x2_ASAP7_75t_L g8073 ( 
.A(n_7920),
.B(n_341),
.Y(n_8073)
);

NAND2xp5_ASAP7_75t_L g8074 ( 
.A(n_7819),
.B(n_415),
.Y(n_8074)
);

INVx1_ASAP7_75t_L g8075 ( 
.A(n_7854),
.Y(n_8075)
);

OAI21xp33_ASAP7_75t_SL g8076 ( 
.A1(n_7843),
.A2(n_417),
.B(n_418),
.Y(n_8076)
);

NOR2xp33_ASAP7_75t_L g8077 ( 
.A(n_7939),
.B(n_418),
.Y(n_8077)
);

AOI22xp33_ASAP7_75t_L g8078 ( 
.A1(n_7861),
.A2(n_3029),
.B1(n_2985),
.B2(n_1781),
.Y(n_8078)
);

NAND2xp5_ASAP7_75t_L g8079 ( 
.A(n_7837),
.B(n_419),
.Y(n_8079)
);

NAND3xp33_ASAP7_75t_L g8080 ( 
.A(n_7898),
.B(n_419),
.C(n_420),
.Y(n_8080)
);

NAND4xp25_ASAP7_75t_L g8081 ( 
.A(n_7818),
.B(n_423),
.C(n_421),
.D(n_422),
.Y(n_8081)
);

AND2x2_ASAP7_75t_L g8082 ( 
.A(n_7906),
.B(n_422),
.Y(n_8082)
);

NAND2xp5_ASAP7_75t_SL g8083 ( 
.A(n_7890),
.B(n_1766),
.Y(n_8083)
);

NAND2xp5_ASAP7_75t_L g8084 ( 
.A(n_7857),
.B(n_7859),
.Y(n_8084)
);

AOI21xp33_ASAP7_75t_L g8085 ( 
.A1(n_7917),
.A2(n_423),
.B(n_424),
.Y(n_8085)
);

NAND2xp5_ASAP7_75t_L g8086 ( 
.A(n_7869),
.B(n_424),
.Y(n_8086)
);

NAND2xp5_ASAP7_75t_L g8087 ( 
.A(n_7870),
.B(n_425),
.Y(n_8087)
);

AOI22xp5_ASAP7_75t_L g8088 ( 
.A1(n_7863),
.A2(n_3029),
.B1(n_1781),
.B2(n_1825),
.Y(n_8088)
);

OAI22xp5_ASAP7_75t_L g8089 ( 
.A1(n_7889),
.A2(n_429),
.B1(n_426),
.B2(n_428),
.Y(n_8089)
);

NAND2xp33_ASAP7_75t_L g8090 ( 
.A(n_7946),
.B(n_3029),
.Y(n_8090)
);

AND2x2_ASAP7_75t_L g8091 ( 
.A(n_7804),
.B(n_430),
.Y(n_8091)
);

AND2x2_ASAP7_75t_L g8092 ( 
.A(n_7899),
.B(n_430),
.Y(n_8092)
);

AND2x2_ASAP7_75t_L g8093 ( 
.A(n_7908),
.B(n_431),
.Y(n_8093)
);

INVx1_ASAP7_75t_L g8094 ( 
.A(n_8059),
.Y(n_8094)
);

AND2x4_ASAP7_75t_L g8095 ( 
.A(n_8008),
.B(n_7872),
.Y(n_8095)
);

AND2x2_ASAP7_75t_L g8096 ( 
.A(n_7964),
.B(n_7914),
.Y(n_8096)
);

BUFx2_ASAP7_75t_L g8097 ( 
.A(n_7971),
.Y(n_8097)
);

INVx2_ASAP7_75t_L g8098 ( 
.A(n_8003),
.Y(n_8098)
);

OR2x2_ASAP7_75t_L g8099 ( 
.A(n_7955),
.B(n_7854),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_8059),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_7953),
.Y(n_8101)
);

AND2x2_ASAP7_75t_L g8102 ( 
.A(n_7954),
.B(n_7947),
.Y(n_8102)
);

INVx2_ASAP7_75t_L g8103 ( 
.A(n_7956),
.Y(n_8103)
);

AND2x4_ASAP7_75t_L g8104 ( 
.A(n_7961),
.B(n_7878),
.Y(n_8104)
);

INVx1_ASAP7_75t_L g8105 ( 
.A(n_8091),
.Y(n_8105)
);

OR2x2_ASAP7_75t_L g8106 ( 
.A(n_8032),
.B(n_7854),
.Y(n_8106)
);

HB1xp67_ASAP7_75t_L g8107 ( 
.A(n_7963),
.Y(n_8107)
);

BUFx2_ASAP7_75t_L g8108 ( 
.A(n_8082),
.Y(n_8108)
);

INVx1_ASAP7_75t_L g8109 ( 
.A(n_8075),
.Y(n_8109)
);

INVx2_ASAP7_75t_L g8110 ( 
.A(n_8056),
.Y(n_8110)
);

NOR2xp33_ASAP7_75t_L g8111 ( 
.A(n_8076),
.B(n_7941),
.Y(n_8111)
);

INVx4_ASAP7_75t_L g8112 ( 
.A(n_8062),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7985),
.Y(n_8113)
);

INVx2_ASAP7_75t_L g8114 ( 
.A(n_8030),
.Y(n_8114)
);

AND2x2_ASAP7_75t_L g8115 ( 
.A(n_8020),
.B(n_7948),
.Y(n_8115)
);

INVx1_ASAP7_75t_L g8116 ( 
.A(n_7987),
.Y(n_8116)
);

NAND2xp5_ASAP7_75t_L g8117 ( 
.A(n_8061),
.B(n_7942),
.Y(n_8117)
);

INVx1_ASAP7_75t_L g8118 ( 
.A(n_8006),
.Y(n_8118)
);

INVxp33_ASAP7_75t_SL g8119 ( 
.A(n_7993),
.Y(n_8119)
);

OR2x2_ASAP7_75t_L g8120 ( 
.A(n_8066),
.B(n_7943),
.Y(n_8120)
);

INVxp67_ASAP7_75t_L g8121 ( 
.A(n_7996),
.Y(n_8121)
);

AND2x2_ASAP7_75t_L g8122 ( 
.A(n_8007),
.B(n_7866),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_8084),
.Y(n_8123)
);

INVx1_ASAP7_75t_L g8124 ( 
.A(n_8067),
.Y(n_8124)
);

AND2x2_ASAP7_75t_L g8125 ( 
.A(n_8010),
.B(n_7867),
.Y(n_8125)
);

AND2x2_ASAP7_75t_L g8126 ( 
.A(n_8015),
.B(n_7873),
.Y(n_8126)
);

OAI22xp5_ASAP7_75t_L g8127 ( 
.A1(n_8014),
.A2(n_7877),
.B1(n_7874),
.B2(n_434),
.Y(n_8127)
);

AND2x2_ASAP7_75t_L g8128 ( 
.A(n_8045),
.B(n_431),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_8068),
.Y(n_8129)
);

AND2x2_ASAP7_75t_L g8130 ( 
.A(n_8009),
.B(n_432),
.Y(n_8130)
);

INVx1_ASAP7_75t_L g8131 ( 
.A(n_8044),
.Y(n_8131)
);

OR2x2_ASAP7_75t_L g8132 ( 
.A(n_7958),
.B(n_432),
.Y(n_8132)
);

AND2x2_ASAP7_75t_L g8133 ( 
.A(n_8071),
.B(n_434),
.Y(n_8133)
);

HB1xp67_ASAP7_75t_L g8134 ( 
.A(n_7994),
.Y(n_8134)
);

NOR2xp33_ASAP7_75t_L g8135 ( 
.A(n_8047),
.B(n_8053),
.Y(n_8135)
);

NOR2xp33_ASAP7_75t_L g8136 ( 
.A(n_8054),
.B(n_435),
.Y(n_8136)
);

OR2x2_ASAP7_75t_L g8137 ( 
.A(n_8019),
.B(n_436),
.Y(n_8137)
);

HB1xp67_ASAP7_75t_L g8138 ( 
.A(n_7983),
.Y(n_8138)
);

HB1xp67_ASAP7_75t_L g8139 ( 
.A(n_7983),
.Y(n_8139)
);

INVx2_ASAP7_75t_L g8140 ( 
.A(n_8092),
.Y(n_8140)
);

BUFx2_ASAP7_75t_L g8141 ( 
.A(n_7972),
.Y(n_8141)
);

BUFx3_ASAP7_75t_L g8142 ( 
.A(n_7992),
.Y(n_8142)
);

AND2x4_ASAP7_75t_L g8143 ( 
.A(n_7990),
.B(n_436),
.Y(n_8143)
);

INVx2_ASAP7_75t_L g8144 ( 
.A(n_8093),
.Y(n_8144)
);

AND2x4_ASAP7_75t_L g8145 ( 
.A(n_8073),
.B(n_437),
.Y(n_8145)
);

BUFx2_ASAP7_75t_SL g8146 ( 
.A(n_7968),
.Y(n_8146)
);

INVx2_ASAP7_75t_L g8147 ( 
.A(n_8026),
.Y(n_8147)
);

INVx2_ASAP7_75t_L g8148 ( 
.A(n_8016),
.Y(n_8148)
);

INVx4_ASAP7_75t_L g8149 ( 
.A(n_8024),
.Y(n_8149)
);

INVx2_ASAP7_75t_L g8150 ( 
.A(n_8004),
.Y(n_8150)
);

NAND2x1p5_ASAP7_75t_L g8151 ( 
.A(n_8077),
.B(n_437),
.Y(n_8151)
);

INVx1_ASAP7_75t_L g8152 ( 
.A(n_8086),
.Y(n_8152)
);

AND2x2_ASAP7_75t_L g8153 ( 
.A(n_8022),
.B(n_438),
.Y(n_8153)
);

OR2x2_ASAP7_75t_L g8154 ( 
.A(n_7979),
.B(n_438),
.Y(n_8154)
);

INVx1_ASAP7_75t_L g8155 ( 
.A(n_8087),
.Y(n_8155)
);

INVx1_ASAP7_75t_L g8156 ( 
.A(n_8070),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_7960),
.Y(n_8157)
);

INVx1_ASAP7_75t_L g8158 ( 
.A(n_7980),
.Y(n_8158)
);

AND2x4_ASAP7_75t_L g8159 ( 
.A(n_7962),
.B(n_439),
.Y(n_8159)
);

AND2x2_ASAP7_75t_L g8160 ( 
.A(n_8048),
.B(n_440),
.Y(n_8160)
);

INVx1_ASAP7_75t_L g8161 ( 
.A(n_8036),
.Y(n_8161)
);

HB1xp67_ASAP7_75t_L g8162 ( 
.A(n_7975),
.Y(n_8162)
);

INVx1_ASAP7_75t_L g8163 ( 
.A(n_8039),
.Y(n_8163)
);

INVx1_ASAP7_75t_L g8164 ( 
.A(n_8042),
.Y(n_8164)
);

AND2x4_ASAP7_75t_L g8165 ( 
.A(n_8031),
.B(n_440),
.Y(n_8165)
);

OR2x2_ASAP7_75t_L g8166 ( 
.A(n_8049),
.B(n_441),
.Y(n_8166)
);

AND2x2_ASAP7_75t_L g8167 ( 
.A(n_7952),
.B(n_441),
.Y(n_8167)
);

INVxp67_ASAP7_75t_L g8168 ( 
.A(n_7965),
.Y(n_8168)
);

AND2x2_ASAP7_75t_L g8169 ( 
.A(n_7957),
.B(n_442),
.Y(n_8169)
);

INVxp67_ASAP7_75t_L g8170 ( 
.A(n_8005),
.Y(n_8170)
);

INVxp67_ASAP7_75t_L g8171 ( 
.A(n_8041),
.Y(n_8171)
);

AND2x4_ASAP7_75t_L g8172 ( 
.A(n_7989),
.B(n_444),
.Y(n_8172)
);

INVx2_ASAP7_75t_L g8173 ( 
.A(n_8055),
.Y(n_8173)
);

AOI22xp33_ASAP7_75t_L g8174 ( 
.A1(n_7959),
.A2(n_3029),
.B1(n_1781),
.B2(n_1825),
.Y(n_8174)
);

NAND2xp5_ASAP7_75t_L g8175 ( 
.A(n_7970),
.B(n_444),
.Y(n_8175)
);

NAND2xp5_ASAP7_75t_L g8176 ( 
.A(n_7978),
.B(n_445),
.Y(n_8176)
);

NOR2xp33_ASAP7_75t_L g8177 ( 
.A(n_8065),
.B(n_447),
.Y(n_8177)
);

INVx1_ASAP7_75t_SL g8178 ( 
.A(n_8023),
.Y(n_8178)
);

INVx1_ASAP7_75t_L g8179 ( 
.A(n_8034),
.Y(n_8179)
);

AND2x4_ASAP7_75t_L g8180 ( 
.A(n_8052),
.B(n_448),
.Y(n_8180)
);

OR2x2_ASAP7_75t_L g8181 ( 
.A(n_7988),
.B(n_449),
.Y(n_8181)
);

INVx2_ASAP7_75t_L g8182 ( 
.A(n_8057),
.Y(n_8182)
);

AND2x4_ASAP7_75t_L g8183 ( 
.A(n_8052),
.B(n_449),
.Y(n_8183)
);

AND2x2_ASAP7_75t_L g8184 ( 
.A(n_8046),
.B(n_8040),
.Y(n_8184)
);

NAND2xp5_ASAP7_75t_L g8185 ( 
.A(n_7967),
.B(n_450),
.Y(n_8185)
);

INVx2_ASAP7_75t_L g8186 ( 
.A(n_8058),
.Y(n_8186)
);

AND2x2_ASAP7_75t_L g8187 ( 
.A(n_7986),
.B(n_451),
.Y(n_8187)
);

NOR2xp67_ASAP7_75t_L g8188 ( 
.A(n_8080),
.B(n_453),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_8011),
.Y(n_8189)
);

INVx1_ASAP7_75t_L g8190 ( 
.A(n_8080),
.Y(n_8190)
);

INVx2_ASAP7_75t_L g8191 ( 
.A(n_8037),
.Y(n_8191)
);

HB1xp67_ASAP7_75t_L g8192 ( 
.A(n_8001),
.Y(n_8192)
);

INVx2_ASAP7_75t_L g8193 ( 
.A(n_7999),
.Y(n_8193)
);

INVx3_ASAP7_75t_L g8194 ( 
.A(n_8043),
.Y(n_8194)
);

INVx2_ASAP7_75t_L g8195 ( 
.A(n_8074),
.Y(n_8195)
);

AND2x2_ASAP7_75t_L g8196 ( 
.A(n_8060),
.B(n_453),
.Y(n_8196)
);

INVx1_ASAP7_75t_L g8197 ( 
.A(n_7974),
.Y(n_8197)
);

NOR2xp33_ASAP7_75t_L g8198 ( 
.A(n_8081),
.B(n_454),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_7974),
.Y(n_8199)
);

NAND2xp5_ASAP7_75t_L g8200 ( 
.A(n_8028),
.B(n_454),
.Y(n_8200)
);

INVxp67_ASAP7_75t_SL g8201 ( 
.A(n_7998),
.Y(n_8201)
);

INVx1_ASAP7_75t_L g8202 ( 
.A(n_8029),
.Y(n_8202)
);

AND2x2_ASAP7_75t_L g8203 ( 
.A(n_7995),
.B(n_455),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_8033),
.Y(n_8204)
);

AND2x2_ASAP7_75t_L g8205 ( 
.A(n_8063),
.B(n_455),
.Y(n_8205)
);

AND2x2_ASAP7_75t_L g8206 ( 
.A(n_7991),
.B(n_456),
.Y(n_8206)
);

INVx1_ASAP7_75t_L g8207 ( 
.A(n_7984),
.Y(n_8207)
);

INVx3_ASAP7_75t_L g8208 ( 
.A(n_8079),
.Y(n_8208)
);

AND2x2_ASAP7_75t_L g8209 ( 
.A(n_8027),
.B(n_7973),
.Y(n_8209)
);

INVx1_ASAP7_75t_L g8210 ( 
.A(n_7984),
.Y(n_8210)
);

INVx3_ASAP7_75t_L g8211 ( 
.A(n_8025),
.Y(n_8211)
);

AND2x2_ASAP7_75t_L g8212 ( 
.A(n_7981),
.B(n_460),
.Y(n_8212)
);

NAND2xp5_ASAP7_75t_L g8213 ( 
.A(n_8035),
.B(n_461),
.Y(n_8213)
);

AND2x2_ASAP7_75t_L g8214 ( 
.A(n_7966),
.B(n_462),
.Y(n_8214)
);

INVx2_ASAP7_75t_L g8215 ( 
.A(n_8021),
.Y(n_8215)
);

NAND2xp5_ASAP7_75t_L g8216 ( 
.A(n_8089),
.B(n_463),
.Y(n_8216)
);

OAI21x1_ASAP7_75t_L g8217 ( 
.A1(n_8094),
.A2(n_7969),
.B(n_7997),
.Y(n_8217)
);

INVx2_ASAP7_75t_L g8218 ( 
.A(n_8151),
.Y(n_8218)
);

INVx1_ASAP7_75t_L g8219 ( 
.A(n_8094),
.Y(n_8219)
);

OA21x2_ASAP7_75t_L g8220 ( 
.A1(n_8100),
.A2(n_7982),
.B(n_8000),
.Y(n_8220)
);

INVx1_ASAP7_75t_L g8221 ( 
.A(n_8100),
.Y(n_8221)
);

INVx1_ASAP7_75t_L g8222 ( 
.A(n_8138),
.Y(n_8222)
);

INVx1_ASAP7_75t_L g8223 ( 
.A(n_8139),
.Y(n_8223)
);

OAI21x1_ASAP7_75t_L g8224 ( 
.A1(n_8106),
.A2(n_8018),
.B(n_8017),
.Y(n_8224)
);

OA21x2_ASAP7_75t_L g8225 ( 
.A1(n_8197),
.A2(n_7976),
.B(n_8002),
.Y(n_8225)
);

INVx1_ASAP7_75t_L g8226 ( 
.A(n_8107),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_8146),
.Y(n_8227)
);

NAND2xp5_ASAP7_75t_SL g8228 ( 
.A(n_8119),
.B(n_8012),
.Y(n_8228)
);

INVx1_ASAP7_75t_L g8229 ( 
.A(n_8141),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_8197),
.Y(n_8230)
);

OAI21x1_ASAP7_75t_L g8231 ( 
.A1(n_8098),
.A2(n_8050),
.B(n_8013),
.Y(n_8231)
);

NAND2xp5_ASAP7_75t_L g8232 ( 
.A(n_8112),
.B(n_8085),
.Y(n_8232)
);

INVx2_ASAP7_75t_L g8233 ( 
.A(n_8095),
.Y(n_8233)
);

INVx2_ASAP7_75t_L g8234 ( 
.A(n_8095),
.Y(n_8234)
);

INVx2_ASAP7_75t_L g8235 ( 
.A(n_8112),
.Y(n_8235)
);

OAI21x1_ASAP7_75t_L g8236 ( 
.A1(n_8099),
.A2(n_8083),
.B(n_8038),
.Y(n_8236)
);

BUFx3_ASAP7_75t_L g8237 ( 
.A(n_8097),
.Y(n_8237)
);

NOR2x1p5_ASAP7_75t_L g8238 ( 
.A(n_8103),
.B(n_8069),
.Y(n_8238)
);

OAI21x1_ASAP7_75t_L g8239 ( 
.A1(n_8101),
.A2(n_8002),
.B(n_8064),
.Y(n_8239)
);

INVx1_ASAP7_75t_SL g8240 ( 
.A(n_8178),
.Y(n_8240)
);

AND2x4_ASAP7_75t_L g8241 ( 
.A(n_8104),
.B(n_8072),
.Y(n_8241)
);

INVxp67_ASAP7_75t_SL g8242 ( 
.A(n_8207),
.Y(n_8242)
);

INVx2_ASAP7_75t_SL g8243 ( 
.A(n_8104),
.Y(n_8243)
);

HB1xp67_ASAP7_75t_L g8244 ( 
.A(n_8207),
.Y(n_8244)
);

INVx1_ASAP7_75t_L g8245 ( 
.A(n_8199),
.Y(n_8245)
);

INVxp67_ASAP7_75t_SL g8246 ( 
.A(n_8210),
.Y(n_8246)
);

INVx1_ASAP7_75t_L g8247 ( 
.A(n_8199),
.Y(n_8247)
);

NOR2xp33_ASAP7_75t_L g8248 ( 
.A(n_8171),
.B(n_7977),
.Y(n_8248)
);

OA21x2_ASAP7_75t_L g8249 ( 
.A1(n_8210),
.A2(n_8088),
.B(n_8051),
.Y(n_8249)
);

AOI21xp33_ASAP7_75t_L g8250 ( 
.A1(n_8101),
.A2(n_8090),
.B(n_8078),
.Y(n_8250)
);

INVx2_ASAP7_75t_L g8251 ( 
.A(n_8145),
.Y(n_8251)
);

INVx4_ASAP7_75t_SL g8252 ( 
.A(n_8142),
.Y(n_8252)
);

INVx2_ASAP7_75t_L g8253 ( 
.A(n_8145),
.Y(n_8253)
);

INVxp67_ASAP7_75t_L g8254 ( 
.A(n_8108),
.Y(n_8254)
);

INVx1_ASAP7_75t_L g8255 ( 
.A(n_8102),
.Y(n_8255)
);

OAI21x1_ASAP7_75t_L g8256 ( 
.A1(n_8206),
.A2(n_463),
.B(n_464),
.Y(n_8256)
);

AND2x2_ASAP7_75t_L g8257 ( 
.A(n_8115),
.B(n_465),
.Y(n_8257)
);

BUFx2_ASAP7_75t_L g8258 ( 
.A(n_8159),
.Y(n_8258)
);

HB1xp67_ASAP7_75t_L g8259 ( 
.A(n_8180),
.Y(n_8259)
);

INVx1_ASAP7_75t_SL g8260 ( 
.A(n_8166),
.Y(n_8260)
);

BUFx2_ASAP7_75t_L g8261 ( 
.A(n_8159),
.Y(n_8261)
);

INVx1_ASAP7_75t_L g8262 ( 
.A(n_8105),
.Y(n_8262)
);

INVx1_ASAP7_75t_L g8263 ( 
.A(n_8180),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_8105),
.Y(n_8264)
);

NAND2xp5_ASAP7_75t_SL g8265 ( 
.A(n_8183),
.B(n_1766),
.Y(n_8265)
);

NAND3xp33_ASAP7_75t_SL g8266 ( 
.A(n_8209),
.B(n_466),
.C(n_468),
.Y(n_8266)
);

OAI21xp5_ASAP7_75t_L g8267 ( 
.A1(n_8201),
.A2(n_8169),
.B(n_8167),
.Y(n_8267)
);

AND2x2_ASAP7_75t_L g8268 ( 
.A(n_8126),
.B(n_466),
.Y(n_8268)
);

INVx2_ASAP7_75t_L g8269 ( 
.A(n_8130),
.Y(n_8269)
);

OR2x6_ASAP7_75t_L g8270 ( 
.A(n_8121),
.B(n_2433),
.Y(n_8270)
);

INVxp67_ASAP7_75t_SL g8271 ( 
.A(n_8200),
.Y(n_8271)
);

INVx1_ASAP7_75t_L g8272 ( 
.A(n_8125),
.Y(n_8272)
);

BUFx2_ASAP7_75t_L g8273 ( 
.A(n_8128),
.Y(n_8273)
);

BUFx2_ASAP7_75t_L g8274 ( 
.A(n_8122),
.Y(n_8274)
);

INVx2_ASAP7_75t_L g8275 ( 
.A(n_8154),
.Y(n_8275)
);

INVx1_ASAP7_75t_L g8276 ( 
.A(n_8183),
.Y(n_8276)
);

INVx1_ASAP7_75t_L g8277 ( 
.A(n_8212),
.Y(n_8277)
);

INVx1_ASAP7_75t_SL g8278 ( 
.A(n_8120),
.Y(n_8278)
);

INVx4_ASAP7_75t_L g8279 ( 
.A(n_8134),
.Y(n_8279)
);

OA21x2_ASAP7_75t_L g8280 ( 
.A1(n_8202),
.A2(n_468),
.B(n_469),
.Y(n_8280)
);

NOR2x1p5_ASAP7_75t_L g8281 ( 
.A(n_8110),
.B(n_469),
.Y(n_8281)
);

INVx1_ASAP7_75t_L g8282 ( 
.A(n_8160),
.Y(n_8282)
);

INVx3_ASAP7_75t_L g8283 ( 
.A(n_8143),
.Y(n_8283)
);

OAI21x1_ASAP7_75t_L g8284 ( 
.A1(n_8185),
.A2(n_471),
.B(n_472),
.Y(n_8284)
);

INVx1_ASAP7_75t_L g8285 ( 
.A(n_8133),
.Y(n_8285)
);

INVx1_ASAP7_75t_L g8286 ( 
.A(n_8208),
.Y(n_8286)
);

INVx5_ASAP7_75t_L g8287 ( 
.A(n_8143),
.Y(n_8287)
);

INVx2_ASAP7_75t_SL g8288 ( 
.A(n_8096),
.Y(n_8288)
);

NAND2xp5_ASAP7_75t_L g8289 ( 
.A(n_8188),
.B(n_473),
.Y(n_8289)
);

OR2x2_ASAP7_75t_SL g8290 ( 
.A(n_8162),
.B(n_475),
.Y(n_8290)
);

NOR2xp33_ASAP7_75t_L g8291 ( 
.A(n_8190),
.B(n_476),
.Y(n_8291)
);

OR2x2_ASAP7_75t_L g8292 ( 
.A(n_8181),
.B(n_476),
.Y(n_8292)
);

INVx1_ASAP7_75t_L g8293 ( 
.A(n_8208),
.Y(n_8293)
);

INVx2_ASAP7_75t_L g8294 ( 
.A(n_8140),
.Y(n_8294)
);

INVx4_ASAP7_75t_L g8295 ( 
.A(n_8137),
.Y(n_8295)
);

INVx2_ASAP7_75t_L g8296 ( 
.A(n_8144),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_8194),
.Y(n_8297)
);

INVx1_ASAP7_75t_L g8298 ( 
.A(n_8194),
.Y(n_8298)
);

NAND2xp33_ASAP7_75t_R g8299 ( 
.A(n_8172),
.B(n_8187),
.Y(n_8299)
);

NOR3xp33_ASAP7_75t_SL g8300 ( 
.A(n_8127),
.B(n_477),
.C(n_479),
.Y(n_8300)
);

AND2x2_ASAP7_75t_L g8301 ( 
.A(n_8184),
.B(n_8150),
.Y(n_8301)
);

AND2x2_ASAP7_75t_L g8302 ( 
.A(n_8147),
.B(n_477),
.Y(n_8302)
);

NAND2xp5_ASAP7_75t_L g8303 ( 
.A(n_8135),
.B(n_479),
.Y(n_8303)
);

INVx1_ASAP7_75t_L g8304 ( 
.A(n_8190),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_8175),
.Y(n_8305)
);

AND2x2_ASAP7_75t_L g8306 ( 
.A(n_8203),
.B(n_8113),
.Y(n_8306)
);

AND2x4_ASAP7_75t_L g8307 ( 
.A(n_8153),
.B(n_480),
.Y(n_8307)
);

INVx1_ASAP7_75t_L g8308 ( 
.A(n_8123),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_8252),
.B(n_8148),
.Y(n_8309)
);

AND2x2_ASAP7_75t_L g8310 ( 
.A(n_8252),
.B(n_8111),
.Y(n_8310)
);

INVx1_ASAP7_75t_L g8311 ( 
.A(n_8244),
.Y(n_8311)
);

INVx1_ASAP7_75t_L g8312 ( 
.A(n_8242),
.Y(n_8312)
);

INVx1_ASAP7_75t_L g8313 ( 
.A(n_8246),
.Y(n_8313)
);

AND2x2_ASAP7_75t_L g8314 ( 
.A(n_8274),
.B(n_8117),
.Y(n_8314)
);

OR2x2_ASAP7_75t_L g8315 ( 
.A(n_8243),
.B(n_8179),
.Y(n_8315)
);

AND2x2_ASAP7_75t_L g8316 ( 
.A(n_8237),
.B(n_8114),
.Y(n_8316)
);

INVx2_ASAP7_75t_SL g8317 ( 
.A(n_8287),
.Y(n_8317)
);

INVx1_ASAP7_75t_L g8318 ( 
.A(n_8258),
.Y(n_8318)
);

INVx1_ASAP7_75t_L g8319 ( 
.A(n_8261),
.Y(n_8319)
);

AND2x2_ASAP7_75t_L g8320 ( 
.A(n_8229),
.B(n_8172),
.Y(n_8320)
);

INVx2_ASAP7_75t_L g8321 ( 
.A(n_8290),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_8259),
.Y(n_8322)
);

AND2x2_ASAP7_75t_L g8323 ( 
.A(n_8240),
.B(n_8149),
.Y(n_8323)
);

AND2x4_ASAP7_75t_L g8324 ( 
.A(n_8233),
.B(n_8116),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_8234),
.Y(n_8325)
);

AND2x4_ASAP7_75t_L g8326 ( 
.A(n_8287),
.B(n_8156),
.Y(n_8326)
);

OR2x2_ASAP7_75t_L g8327 ( 
.A(n_8279),
.B(n_8179),
.Y(n_8327)
);

INVx2_ASAP7_75t_SL g8328 ( 
.A(n_8287),
.Y(n_8328)
);

AND2x2_ASAP7_75t_L g8329 ( 
.A(n_8288),
.B(n_8149),
.Y(n_8329)
);

INVx1_ASAP7_75t_L g8330 ( 
.A(n_8273),
.Y(n_8330)
);

OR2x2_ASAP7_75t_L g8331 ( 
.A(n_8279),
.B(n_8278),
.Y(n_8331)
);

INVx2_ASAP7_75t_L g8332 ( 
.A(n_8281),
.Y(n_8332)
);

AND2x2_ASAP7_75t_L g8333 ( 
.A(n_8227),
.B(n_8196),
.Y(n_8333)
);

OR2x2_ASAP7_75t_L g8334 ( 
.A(n_8230),
.B(n_8132),
.Y(n_8334)
);

AND2x4_ASAP7_75t_L g8335 ( 
.A(n_8283),
.B(n_8235),
.Y(n_8335)
);

INVx4_ASAP7_75t_L g8336 ( 
.A(n_8283),
.Y(n_8336)
);

AND2x2_ASAP7_75t_L g8337 ( 
.A(n_8255),
.B(n_8158),
.Y(n_8337)
);

INVx1_ASAP7_75t_L g8338 ( 
.A(n_8301),
.Y(n_8338)
);

INVx1_ASAP7_75t_L g8339 ( 
.A(n_8263),
.Y(n_8339)
);

BUFx2_ASAP7_75t_L g8340 ( 
.A(n_8241),
.Y(n_8340)
);

INVx1_ASAP7_75t_L g8341 ( 
.A(n_8263),
.Y(n_8341)
);

OR2x2_ASAP7_75t_L g8342 ( 
.A(n_8245),
.B(n_8247),
.Y(n_8342)
);

HB1xp67_ASAP7_75t_L g8343 ( 
.A(n_8220),
.Y(n_8343)
);

AND2x2_ASAP7_75t_L g8344 ( 
.A(n_8272),
.B(n_8165),
.Y(n_8344)
);

INVx1_ASAP7_75t_SL g8345 ( 
.A(n_8257),
.Y(n_8345)
);

BUFx2_ASAP7_75t_L g8346 ( 
.A(n_8241),
.Y(n_8346)
);

NAND2xp5_ASAP7_75t_L g8347 ( 
.A(n_8268),
.B(n_8177),
.Y(n_8347)
);

NAND2xp5_ASAP7_75t_L g8348 ( 
.A(n_8295),
.B(n_8136),
.Y(n_8348)
);

INVx2_ASAP7_75t_L g8349 ( 
.A(n_8295),
.Y(n_8349)
);

AND2x2_ASAP7_75t_L g8350 ( 
.A(n_8254),
.B(n_8165),
.Y(n_8350)
);

OR2x2_ASAP7_75t_L g8351 ( 
.A(n_8225),
.B(n_8157),
.Y(n_8351)
);

NAND2xp5_ASAP7_75t_L g8352 ( 
.A(n_8307),
.B(n_8198),
.Y(n_8352)
);

NAND2xp5_ASAP7_75t_L g8353 ( 
.A(n_8307),
.B(n_8204),
.Y(n_8353)
);

BUFx2_ASAP7_75t_L g8354 ( 
.A(n_8220),
.Y(n_8354)
);

OR2x2_ASAP7_75t_L g8355 ( 
.A(n_8225),
.B(n_8202),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_8280),
.Y(n_8356)
);

INVxp67_ASAP7_75t_L g8357 ( 
.A(n_8299),
.Y(n_8357)
);

OR2x2_ASAP7_75t_L g8358 ( 
.A(n_8226),
.B(n_8176),
.Y(n_8358)
);

AND2x4_ASAP7_75t_L g8359 ( 
.A(n_8294),
.B(n_8161),
.Y(n_8359)
);

NOR2xp33_ASAP7_75t_L g8360 ( 
.A(n_8266),
.B(n_8204),
.Y(n_8360)
);

INVx1_ASAP7_75t_L g8361 ( 
.A(n_8280),
.Y(n_8361)
);

INVx1_ASAP7_75t_L g8362 ( 
.A(n_8277),
.Y(n_8362)
);

INVx2_ASAP7_75t_SL g8363 ( 
.A(n_8238),
.Y(n_8363)
);

HB1xp67_ASAP7_75t_L g8364 ( 
.A(n_8276),
.Y(n_8364)
);

INVx2_ASAP7_75t_SL g8365 ( 
.A(n_8302),
.Y(n_8365)
);

AND2x2_ASAP7_75t_L g8366 ( 
.A(n_8306),
.B(n_8118),
.Y(n_8366)
);

AND2x2_ASAP7_75t_L g8367 ( 
.A(n_8228),
.B(n_8205),
.Y(n_8367)
);

INVx1_ASAP7_75t_L g8368 ( 
.A(n_8271),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_8285),
.Y(n_8369)
);

INVx1_ASAP7_75t_L g8370 ( 
.A(n_8222),
.Y(n_8370)
);

INVx1_ASAP7_75t_L g8371 ( 
.A(n_8289),
.Y(n_8371)
);

INVx1_ASAP7_75t_L g8372 ( 
.A(n_8282),
.Y(n_8372)
);

NAND2xp5_ASAP7_75t_L g8373 ( 
.A(n_8269),
.B(n_8275),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_8222),
.Y(n_8374)
);

HB1xp67_ASAP7_75t_L g8375 ( 
.A(n_8304),
.Y(n_8375)
);

NAND2xp5_ASAP7_75t_L g8376 ( 
.A(n_8260),
.B(n_8131),
.Y(n_8376)
);

INVx1_ASAP7_75t_L g8377 ( 
.A(n_8223),
.Y(n_8377)
);

AND2x2_ASAP7_75t_L g8378 ( 
.A(n_8262),
.B(n_8163),
.Y(n_8378)
);

INVx3_ASAP7_75t_L g8379 ( 
.A(n_8296),
.Y(n_8379)
);

OR2x2_ASAP7_75t_L g8380 ( 
.A(n_8304),
.B(n_8264),
.Y(n_8380)
);

INVx1_ASAP7_75t_L g8381 ( 
.A(n_8223),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_8219),
.Y(n_8382)
);

INVx2_ASAP7_75t_L g8383 ( 
.A(n_8251),
.Y(n_8383)
);

AND2x2_ASAP7_75t_L g8384 ( 
.A(n_8297),
.B(n_8164),
.Y(n_8384)
);

OR2x2_ASAP7_75t_L g8385 ( 
.A(n_8298),
.B(n_8211),
.Y(n_8385)
);

INVx2_ASAP7_75t_L g8386 ( 
.A(n_8253),
.Y(n_8386)
);

OR2x6_ASAP7_75t_L g8387 ( 
.A(n_8286),
.B(n_8214),
.Y(n_8387)
);

INVx1_ASAP7_75t_L g8388 ( 
.A(n_8354),
.Y(n_8388)
);

NAND2xp5_ASAP7_75t_L g8389 ( 
.A(n_8340),
.B(n_8218),
.Y(n_8389)
);

INVx1_ASAP7_75t_L g8390 ( 
.A(n_8343),
.Y(n_8390)
);

OAI22xp5_ASAP7_75t_L g8391 ( 
.A1(n_8355),
.A2(n_8293),
.B1(n_8308),
.B2(n_8300),
.Y(n_8391)
);

INVx1_ASAP7_75t_L g8392 ( 
.A(n_8375),
.Y(n_8392)
);

NAND2xp5_ASAP7_75t_L g8393 ( 
.A(n_8346),
.B(n_8291),
.Y(n_8393)
);

INVx1_ASAP7_75t_L g8394 ( 
.A(n_8356),
.Y(n_8394)
);

INVx1_ASAP7_75t_L g8395 ( 
.A(n_8361),
.Y(n_8395)
);

OR2x2_ASAP7_75t_L g8396 ( 
.A(n_8331),
.B(n_8239),
.Y(n_8396)
);

OAI211xp5_ASAP7_75t_L g8397 ( 
.A1(n_8351),
.A2(n_8221),
.B(n_8219),
.C(n_8170),
.Y(n_8397)
);

INVx1_ASAP7_75t_L g8398 ( 
.A(n_8379),
.Y(n_8398)
);

OAI33xp33_ASAP7_75t_L g8399 ( 
.A1(n_8370),
.A2(n_8189),
.A3(n_8221),
.B1(n_8232),
.B2(n_8168),
.B3(n_8109),
.Y(n_8399)
);

INVx2_ASAP7_75t_L g8400 ( 
.A(n_8310),
.Y(n_8400)
);

OAI31xp33_ASAP7_75t_L g8401 ( 
.A1(n_8311),
.A2(n_8189),
.A3(n_8192),
.B(n_8211),
.Y(n_8401)
);

OAI32xp33_ASAP7_75t_L g8402 ( 
.A1(n_8311),
.A2(n_8248),
.A3(n_8303),
.B1(n_8215),
.B2(n_8305),
.Y(n_8402)
);

AND2x4_ASAP7_75t_L g8403 ( 
.A(n_8379),
.B(n_8124),
.Y(n_8403)
);

AND2x2_ASAP7_75t_L g8404 ( 
.A(n_8323),
.B(n_8267),
.Y(n_8404)
);

INVx1_ASAP7_75t_L g8405 ( 
.A(n_8353),
.Y(n_8405)
);

OR2x2_ASAP7_75t_L g8406 ( 
.A(n_8327),
.B(n_8338),
.Y(n_8406)
);

HB1xp67_ASAP7_75t_L g8407 ( 
.A(n_8317),
.Y(n_8407)
);

OR2x2_ASAP7_75t_L g8408 ( 
.A(n_8336),
.B(n_8318),
.Y(n_8408)
);

AND2x2_ASAP7_75t_L g8409 ( 
.A(n_8314),
.B(n_8305),
.Y(n_8409)
);

INVx2_ASAP7_75t_L g8410 ( 
.A(n_8336),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_8364),
.Y(n_8411)
);

AOI22xp5_ASAP7_75t_L g8412 ( 
.A1(n_8345),
.A2(n_8129),
.B1(n_8191),
.B2(n_8182),
.Y(n_8412)
);

INVx1_ASAP7_75t_L g8413 ( 
.A(n_8380),
.Y(n_8413)
);

AOI21xp5_ASAP7_75t_L g8414 ( 
.A1(n_8312),
.A2(n_8217),
.B(n_8216),
.Y(n_8414)
);

INVx1_ASAP7_75t_L g8415 ( 
.A(n_8316),
.Y(n_8415)
);

NAND2xp5_ASAP7_75t_L g8416 ( 
.A(n_8326),
.B(n_8152),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_8328),
.Y(n_8417)
);

INVx1_ASAP7_75t_L g8418 ( 
.A(n_8312),
.Y(n_8418)
);

OR2x2_ASAP7_75t_L g8419 ( 
.A(n_8319),
.B(n_8292),
.Y(n_8419)
);

NAND2xp5_ASAP7_75t_L g8420 ( 
.A(n_8326),
.B(n_8155),
.Y(n_8420)
);

INVx1_ASAP7_75t_L g8421 ( 
.A(n_8370),
.Y(n_8421)
);

OR2x2_ASAP7_75t_L g8422 ( 
.A(n_8315),
.B(n_8224),
.Y(n_8422)
);

OR2x2_ASAP7_75t_L g8423 ( 
.A(n_8357),
.B(n_8349),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_8313),
.Y(n_8424)
);

NOR2xp67_ASAP7_75t_SL g8425 ( 
.A(n_8330),
.B(n_8265),
.Y(n_8425)
);

OR2x2_ASAP7_75t_L g8426 ( 
.A(n_8322),
.B(n_8173),
.Y(n_8426)
);

INVx3_ASAP7_75t_L g8427 ( 
.A(n_8335),
.Y(n_8427)
);

INVx1_ASAP7_75t_L g8428 ( 
.A(n_8313),
.Y(n_8428)
);

NAND2xp5_ASAP7_75t_L g8429 ( 
.A(n_8365),
.B(n_8186),
.Y(n_8429)
);

INVx2_ASAP7_75t_SL g8430 ( 
.A(n_8335),
.Y(n_8430)
);

INVx1_ASAP7_75t_L g8431 ( 
.A(n_8377),
.Y(n_8431)
);

INVx2_ASAP7_75t_L g8432 ( 
.A(n_8334),
.Y(n_8432)
);

NAND2xp5_ASAP7_75t_L g8433 ( 
.A(n_8324),
.B(n_8256),
.Y(n_8433)
);

AND2x2_ASAP7_75t_L g8434 ( 
.A(n_8366),
.B(n_8344),
.Y(n_8434)
);

INVx2_ASAP7_75t_L g8435 ( 
.A(n_8332),
.Y(n_8435)
);

NOR2xp67_ASAP7_75t_L g8436 ( 
.A(n_8363),
.B(n_8213),
.Y(n_8436)
);

NAND2xp5_ASAP7_75t_L g8437 ( 
.A(n_8324),
.B(n_8195),
.Y(n_8437)
);

AND2x2_ASAP7_75t_L g8438 ( 
.A(n_8350),
.B(n_8231),
.Y(n_8438)
);

AND2x2_ASAP7_75t_L g8439 ( 
.A(n_8329),
.B(n_8236),
.Y(n_8439)
);

INVx1_ASAP7_75t_L g8440 ( 
.A(n_8382),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_8359),
.B(n_8284),
.Y(n_8441)
);

NAND2xp5_ASAP7_75t_L g8442 ( 
.A(n_8359),
.B(n_8193),
.Y(n_8442)
);

INVx1_ASAP7_75t_L g8443 ( 
.A(n_8382),
.Y(n_8443)
);

AND2x2_ASAP7_75t_L g8444 ( 
.A(n_8320),
.B(n_8270),
.Y(n_8444)
);

INVx1_ASAP7_75t_L g8445 ( 
.A(n_8342),
.Y(n_8445)
);

AND2x2_ASAP7_75t_L g8446 ( 
.A(n_8309),
.B(n_8270),
.Y(n_8446)
);

INVx1_ASAP7_75t_L g8447 ( 
.A(n_8383),
.Y(n_8447)
);

INVx1_ASAP7_75t_L g8448 ( 
.A(n_8386),
.Y(n_8448)
);

AND2x2_ASAP7_75t_L g8449 ( 
.A(n_8333),
.B(n_8337),
.Y(n_8449)
);

INVx2_ASAP7_75t_L g8450 ( 
.A(n_8321),
.Y(n_8450)
);

INVx1_ASAP7_75t_L g8451 ( 
.A(n_8377),
.Y(n_8451)
);

AND2x2_ASAP7_75t_L g8452 ( 
.A(n_8378),
.B(n_8249),
.Y(n_8452)
);

OAI21xp33_ASAP7_75t_L g8453 ( 
.A1(n_8360),
.A2(n_8250),
.B(n_8174),
.Y(n_8453)
);

INVx2_ASAP7_75t_L g8454 ( 
.A(n_8387),
.Y(n_8454)
);

INVx1_ASAP7_75t_L g8455 ( 
.A(n_8427),
.Y(n_8455)
);

AND2x2_ASAP7_75t_L g8456 ( 
.A(n_8449),
.B(n_8384),
.Y(n_8456)
);

INVx2_ASAP7_75t_L g8457 ( 
.A(n_8427),
.Y(n_8457)
);

AND2x2_ASAP7_75t_L g8458 ( 
.A(n_8434),
.B(n_8362),
.Y(n_8458)
);

INVx2_ASAP7_75t_L g8459 ( 
.A(n_8430),
.Y(n_8459)
);

INVx2_ASAP7_75t_L g8460 ( 
.A(n_8452),
.Y(n_8460)
);

NOR2xp67_ASAP7_75t_L g8461 ( 
.A(n_8396),
.B(n_8381),
.Y(n_8461)
);

INVx1_ASAP7_75t_L g8462 ( 
.A(n_8422),
.Y(n_8462)
);

OR2x2_ASAP7_75t_L g8463 ( 
.A(n_8432),
.B(n_8339),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_8390),
.Y(n_8464)
);

INVx1_ASAP7_75t_L g8465 ( 
.A(n_8390),
.Y(n_8465)
);

NOR2xp67_ASAP7_75t_SL g8466 ( 
.A(n_8406),
.B(n_8368),
.Y(n_8466)
);

BUFx2_ASAP7_75t_R g8467 ( 
.A(n_8389),
.Y(n_8467)
);

INVx2_ASAP7_75t_L g8468 ( 
.A(n_8403),
.Y(n_8468)
);

INVx1_ASAP7_75t_L g8469 ( 
.A(n_8437),
.Y(n_8469)
);

NAND2xp5_ASAP7_75t_L g8470 ( 
.A(n_8403),
.B(n_8341),
.Y(n_8470)
);

INVx1_ASAP7_75t_L g8471 ( 
.A(n_8407),
.Y(n_8471)
);

INVx3_ASAP7_75t_SL g8472 ( 
.A(n_8408),
.Y(n_8472)
);

AND2x2_ASAP7_75t_L g8473 ( 
.A(n_8439),
.B(n_8369),
.Y(n_8473)
);

OR2x2_ASAP7_75t_SL g8474 ( 
.A(n_8400),
.B(n_8385),
.Y(n_8474)
);

OR2x2_ASAP7_75t_L g8475 ( 
.A(n_8393),
.B(n_8376),
.Y(n_8475)
);

INVx1_ASAP7_75t_L g8476 ( 
.A(n_8409),
.Y(n_8476)
);

INVx2_ASAP7_75t_L g8477 ( 
.A(n_8419),
.Y(n_8477)
);

NAND2xp5_ASAP7_75t_L g8478 ( 
.A(n_8388),
.B(n_8381),
.Y(n_8478)
);

OAI22xp33_ASAP7_75t_L g8479 ( 
.A1(n_8433),
.A2(n_8387),
.B1(n_8358),
.B2(n_8347),
.Y(n_8479)
);

OAI21xp33_ASAP7_75t_L g8480 ( 
.A1(n_8411),
.A2(n_8373),
.B(n_8372),
.Y(n_8480)
);

AND2x2_ASAP7_75t_L g8481 ( 
.A(n_8404),
.B(n_8325),
.Y(n_8481)
);

INVx1_ASAP7_75t_L g8482 ( 
.A(n_8392),
.Y(n_8482)
);

OR2x2_ASAP7_75t_L g8483 ( 
.A(n_8415),
.B(n_8374),
.Y(n_8483)
);

INVx1_ASAP7_75t_L g8484 ( 
.A(n_8392),
.Y(n_8484)
);

NAND2xp5_ASAP7_75t_L g8485 ( 
.A(n_8421),
.B(n_8367),
.Y(n_8485)
);

NAND2xp5_ASAP7_75t_L g8486 ( 
.A(n_8421),
.B(n_8348),
.Y(n_8486)
);

NAND2xp5_ASAP7_75t_L g8487 ( 
.A(n_8431),
.B(n_8371),
.Y(n_8487)
);

INVx1_ASAP7_75t_L g8488 ( 
.A(n_8442),
.Y(n_8488)
);

AOI32xp33_ASAP7_75t_L g8489 ( 
.A1(n_8438),
.A2(n_8352),
.A3(n_8249),
.B1(n_483),
.B2(n_481),
.Y(n_8489)
);

AND2x2_ASAP7_75t_L g8490 ( 
.A(n_8445),
.B(n_482),
.Y(n_8490)
);

OAI221xp5_ASAP7_75t_SL g8491 ( 
.A1(n_8401),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.C(n_486),
.Y(n_8491)
);

INVxp67_ASAP7_75t_SL g8492 ( 
.A(n_8436),
.Y(n_8492)
);

AND2x2_ASAP7_75t_L g8493 ( 
.A(n_8413),
.B(n_484),
.Y(n_8493)
);

NOR2x1p5_ASAP7_75t_L g8494 ( 
.A(n_8416),
.B(n_486),
.Y(n_8494)
);

AND2x2_ASAP7_75t_L g8495 ( 
.A(n_8405),
.B(n_487),
.Y(n_8495)
);

OAI21xp5_ASAP7_75t_L g8496 ( 
.A1(n_8414),
.A2(n_488),
.B(n_489),
.Y(n_8496)
);

INVx1_ASAP7_75t_L g8497 ( 
.A(n_8431),
.Y(n_8497)
);

INVxp67_ASAP7_75t_SL g8498 ( 
.A(n_8441),
.Y(n_8498)
);

INVxp67_ASAP7_75t_SL g8499 ( 
.A(n_8420),
.Y(n_8499)
);

INVx1_ASAP7_75t_L g8500 ( 
.A(n_8447),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_8448),
.Y(n_8501)
);

AND2x2_ASAP7_75t_L g8502 ( 
.A(n_8398),
.B(n_488),
.Y(n_8502)
);

BUFx2_ASAP7_75t_L g8503 ( 
.A(n_8410),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_8394),
.Y(n_8504)
);

NAND2x1_ASAP7_75t_L g8505 ( 
.A(n_8395),
.B(n_489),
.Y(n_8505)
);

NAND2xp5_ASAP7_75t_L g8506 ( 
.A(n_8456),
.B(n_8450),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_8481),
.Y(n_8507)
);

OAI22xp5_ASAP7_75t_L g8508 ( 
.A1(n_8460),
.A2(n_8463),
.B1(n_8462),
.B2(n_8485),
.Y(n_8508)
);

INVx1_ASAP7_75t_L g8509 ( 
.A(n_8458),
.Y(n_8509)
);

OR2x6_ASAP7_75t_L g8510 ( 
.A(n_8457),
.B(n_8454),
.Y(n_8510)
);

INVxp67_ASAP7_75t_SL g8511 ( 
.A(n_8461),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8473),
.Y(n_8512)
);

INVx1_ASAP7_75t_L g8513 ( 
.A(n_8467),
.Y(n_8513)
);

INVx1_ASAP7_75t_L g8514 ( 
.A(n_8492),
.Y(n_8514)
);

AOI322xp5_ASAP7_75t_L g8515 ( 
.A1(n_8498),
.A2(n_8465),
.A3(n_8464),
.B1(n_8479),
.B2(n_8485),
.C1(n_8435),
.C2(n_8480),
.Y(n_8515)
);

INVx1_ASAP7_75t_L g8516 ( 
.A(n_8461),
.Y(n_8516)
);

INVx1_ASAP7_75t_L g8517 ( 
.A(n_8470),
.Y(n_8517)
);

OR2x2_ASAP7_75t_L g8518 ( 
.A(n_8474),
.B(n_8426),
.Y(n_8518)
);

AOI22xp5_ASAP7_75t_L g8519 ( 
.A1(n_8477),
.A2(n_8391),
.B1(n_8399),
.B2(n_8397),
.Y(n_8519)
);

INVx2_ASAP7_75t_L g8520 ( 
.A(n_8494),
.Y(n_8520)
);

INVx2_ASAP7_75t_L g8521 ( 
.A(n_8475),
.Y(n_8521)
);

INVx1_ASAP7_75t_L g8522 ( 
.A(n_8503),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_8499),
.Y(n_8523)
);

OAI211xp5_ASAP7_75t_L g8524 ( 
.A1(n_8480),
.A2(n_8402),
.B(n_8417),
.C(n_8418),
.Y(n_8524)
);

NOR2xp67_ASAP7_75t_L g8525 ( 
.A(n_8476),
.B(n_8451),
.Y(n_8525)
);

INVx2_ASAP7_75t_SL g8526 ( 
.A(n_8468),
.Y(n_8526)
);

AOI22xp5_ASAP7_75t_L g8527 ( 
.A1(n_8500),
.A2(n_8412),
.B1(n_8429),
.B2(n_8428),
.Y(n_8527)
);

INVx2_ASAP7_75t_L g8528 ( 
.A(n_8505),
.Y(n_8528)
);

AOI22xp33_ASAP7_75t_L g8529 ( 
.A1(n_8501),
.A2(n_8424),
.B1(n_8443),
.B2(n_8440),
.Y(n_8529)
);

OAI21xp33_ASAP7_75t_L g8530 ( 
.A1(n_8471),
.A2(n_8423),
.B(n_8446),
.Y(n_8530)
);

OR2x2_ASAP7_75t_L g8531 ( 
.A(n_8472),
.B(n_8444),
.Y(n_8531)
);

AOI21xp33_ASAP7_75t_SL g8532 ( 
.A1(n_8455),
.A2(n_8496),
.B(n_8489),
.Y(n_8532)
);

NAND2x1_ASAP7_75t_L g8533 ( 
.A(n_8466),
.B(n_8425),
.Y(n_8533)
);

OAI322xp33_ASAP7_75t_L g8534 ( 
.A1(n_8478),
.A2(n_8402),
.A3(n_8453),
.B1(n_492),
.B2(n_493),
.C1(n_494),
.C2(n_496),
.Y(n_8534)
);

INVx1_ASAP7_75t_L g8535 ( 
.A(n_8483),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_L g8536 ( 
.A(n_8493),
.B(n_8490),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_8459),
.Y(n_8537)
);

AOI22xp5_ASAP7_75t_L g8538 ( 
.A1(n_8486),
.A2(n_8504),
.B1(n_8484),
.B2(n_8482),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_8478),
.Y(n_8539)
);

INVx1_ASAP7_75t_SL g8540 ( 
.A(n_8518),
.Y(n_8540)
);

NAND3x2_ASAP7_75t_L g8541 ( 
.A(n_8531),
.B(n_8488),
.C(n_8469),
.Y(n_8541)
);

OAI22xp33_ASAP7_75t_L g8542 ( 
.A1(n_8538),
.A2(n_8486),
.B1(n_8487),
.B2(n_8497),
.Y(n_8542)
);

NAND2xp5_ASAP7_75t_L g8543 ( 
.A(n_8521),
.B(n_8495),
.Y(n_8543)
);

AND2x2_ASAP7_75t_L g8544 ( 
.A(n_8513),
.B(n_8507),
.Y(n_8544)
);

OAI21xp5_ASAP7_75t_L g8545 ( 
.A1(n_8506),
.A2(n_8496),
.B(n_8487),
.Y(n_8545)
);

NAND2xp5_ASAP7_75t_L g8546 ( 
.A(n_8522),
.B(n_8502),
.Y(n_8546)
);

NOR2x1_ASAP7_75t_L g8547 ( 
.A(n_8533),
.B(n_8491),
.Y(n_8547)
);

AOI22xp5_ASAP7_75t_L g8548 ( 
.A1(n_8511),
.A2(n_2433),
.B1(n_493),
.B2(n_490),
.Y(n_8548)
);

INVx2_ASAP7_75t_L g8549 ( 
.A(n_8528),
.Y(n_8549)
);

NAND2xp5_ASAP7_75t_L g8550 ( 
.A(n_8526),
.B(n_490),
.Y(n_8550)
);

INVxp67_ASAP7_75t_L g8551 ( 
.A(n_8510),
.Y(n_8551)
);

NAND2xp5_ASAP7_75t_L g8552 ( 
.A(n_8512),
.B(n_491),
.Y(n_8552)
);

AOI22xp5_ASAP7_75t_L g8553 ( 
.A1(n_8516),
.A2(n_8525),
.B1(n_8535),
.B2(n_8539),
.Y(n_8553)
);

NAND2xp5_ASAP7_75t_L g8554 ( 
.A(n_8515),
.B(n_496),
.Y(n_8554)
);

NAND2xp5_ASAP7_75t_L g8555 ( 
.A(n_8509),
.B(n_497),
.Y(n_8555)
);

OR2x2_ASAP7_75t_L g8556 ( 
.A(n_8508),
.B(n_498),
.Y(n_8556)
);

AOI322xp5_ASAP7_75t_L g8557 ( 
.A1(n_8519),
.A2(n_499),
.A3(n_500),
.B1(n_501),
.B2(n_502),
.C1(n_503),
.C2(n_505),
.Y(n_8557)
);

A2O1A1Ixp33_ASAP7_75t_L g8558 ( 
.A1(n_8514),
.A2(n_505),
.B(n_500),
.C(n_503),
.Y(n_8558)
);

INVx1_ASAP7_75t_L g8559 ( 
.A(n_8510),
.Y(n_8559)
);

AND2x2_ASAP7_75t_L g8560 ( 
.A(n_8537),
.B(n_507),
.Y(n_8560)
);

INVx1_ASAP7_75t_L g8561 ( 
.A(n_8536),
.Y(n_8561)
);

INVx2_ASAP7_75t_L g8562 ( 
.A(n_8520),
.Y(n_8562)
);

INVx1_ASAP7_75t_L g8563 ( 
.A(n_8523),
.Y(n_8563)
);

INVx1_ASAP7_75t_L g8564 ( 
.A(n_8527),
.Y(n_8564)
);

INVx1_ASAP7_75t_L g8565 ( 
.A(n_8524),
.Y(n_8565)
);

INVx1_ASAP7_75t_L g8566 ( 
.A(n_8534),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_8517),
.Y(n_8567)
);

AOI21xp33_ASAP7_75t_L g8568 ( 
.A1(n_8529),
.A2(n_507),
.B(n_508),
.Y(n_8568)
);

INVxp67_ASAP7_75t_SL g8569 ( 
.A(n_8530),
.Y(n_8569)
);

OAI21xp5_ASAP7_75t_SL g8570 ( 
.A1(n_8532),
.A2(n_508),
.B(n_509),
.Y(n_8570)
);

BUFx2_ASAP7_75t_L g8571 ( 
.A(n_8510),
.Y(n_8571)
);

INVx1_ASAP7_75t_L g8572 ( 
.A(n_8506),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_8506),
.Y(n_8573)
);

INVx1_ASAP7_75t_L g8574 ( 
.A(n_8571),
.Y(n_8574)
);

INVxp67_ASAP7_75t_L g8575 ( 
.A(n_8559),
.Y(n_8575)
);

NOR2xp33_ASAP7_75t_L g8576 ( 
.A(n_8551),
.B(n_509),
.Y(n_8576)
);

AND2x2_ASAP7_75t_L g8577 ( 
.A(n_8540),
.B(n_510),
.Y(n_8577)
);

AO221x1_ASAP7_75t_L g8578 ( 
.A1(n_8542),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.C(n_513),
.Y(n_8578)
);

AOI22xp33_ASAP7_75t_L g8579 ( 
.A1(n_8565),
.A2(n_1825),
.B1(n_1878),
.B2(n_1781),
.Y(n_8579)
);

OAI32xp33_ASAP7_75t_L g8580 ( 
.A1(n_8572),
.A2(n_514),
.A3(n_511),
.B1(n_513),
.B2(n_515),
.Y(n_8580)
);

INVx1_ASAP7_75t_L g8581 ( 
.A(n_8564),
.Y(n_8581)
);

AOI21xp33_ASAP7_75t_L g8582 ( 
.A1(n_8543),
.A2(n_514),
.B(n_515),
.Y(n_8582)
);

O2A1O1Ixp33_ASAP7_75t_L g8583 ( 
.A1(n_8554),
.A2(n_8545),
.B(n_8549),
.C(n_8573),
.Y(n_8583)
);

INVx2_ASAP7_75t_SL g8584 ( 
.A(n_8544),
.Y(n_8584)
);

AOI22xp5_ASAP7_75t_L g8585 ( 
.A1(n_8553),
.A2(n_2433),
.B1(n_520),
.B2(n_516),
.Y(n_8585)
);

XOR2x2_ASAP7_75t_L g8586 ( 
.A(n_8547),
.B(n_516),
.Y(n_8586)
);

OR2x2_ASAP7_75t_L g8587 ( 
.A(n_8541),
.B(n_517),
.Y(n_8587)
);

OR2x2_ASAP7_75t_L g8588 ( 
.A(n_8556),
.B(n_521),
.Y(n_8588)
);

INVx1_ASAP7_75t_L g8589 ( 
.A(n_8560),
.Y(n_8589)
);

OAI21xp33_ASAP7_75t_L g8590 ( 
.A1(n_8569),
.A2(n_522),
.B(n_523),
.Y(n_8590)
);

OAI221xp5_ASAP7_75t_L g8591 ( 
.A1(n_8553),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.C(n_525),
.Y(n_8591)
);

INVxp67_ASAP7_75t_L g8592 ( 
.A(n_8546),
.Y(n_8592)
);

INVx1_ASAP7_75t_L g8593 ( 
.A(n_8550),
.Y(n_8593)
);

BUFx2_ASAP7_75t_L g8594 ( 
.A(n_8567),
.Y(n_8594)
);

AOI21xp33_ASAP7_75t_SL g8595 ( 
.A1(n_8568),
.A2(n_524),
.B(n_526),
.Y(n_8595)
);

AND2x2_ASAP7_75t_L g8596 ( 
.A(n_8561),
.B(n_527),
.Y(n_8596)
);

O2A1O1Ixp33_ASAP7_75t_SL g8597 ( 
.A1(n_8563),
.A2(n_533),
.B(n_530),
.C(n_531),
.Y(n_8597)
);

OR2x2_ASAP7_75t_L g8598 ( 
.A(n_8562),
.B(n_530),
.Y(n_8598)
);

INVx2_ASAP7_75t_L g8599 ( 
.A(n_8566),
.Y(n_8599)
);

INVx1_ASAP7_75t_L g8600 ( 
.A(n_8552),
.Y(n_8600)
);

INVx1_ASAP7_75t_L g8601 ( 
.A(n_8555),
.Y(n_8601)
);

INVx2_ASAP7_75t_L g8602 ( 
.A(n_8548),
.Y(n_8602)
);

HB1xp67_ASAP7_75t_L g8603 ( 
.A(n_8570),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_8558),
.Y(n_8604)
);

OAI21xp5_ASAP7_75t_L g8605 ( 
.A1(n_8557),
.A2(n_533),
.B(n_534),
.Y(n_8605)
);

INVx1_ASAP7_75t_SL g8606 ( 
.A(n_8540),
.Y(n_8606)
);

OR2x2_ASAP7_75t_L g8607 ( 
.A(n_8540),
.B(n_534),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_8571),
.Y(n_8608)
);

INVx1_ASAP7_75t_L g8609 ( 
.A(n_8571),
.Y(n_8609)
);

OAI22xp5_ASAP7_75t_L g8610 ( 
.A1(n_8540),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_8610)
);

INVx1_ASAP7_75t_SL g8611 ( 
.A(n_8606),
.Y(n_8611)
);

AOI22xp5_ASAP7_75t_L g8612 ( 
.A1(n_8594),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_8612)
);

AOI21xp5_ASAP7_75t_L g8613 ( 
.A1(n_8584),
.A2(n_538),
.B(n_539),
.Y(n_8613)
);

OAI321xp33_ASAP7_75t_L g8614 ( 
.A1(n_8574),
.A2(n_1977),
.A3(n_1949),
.B1(n_1878),
.B2(n_1825),
.C(n_542),
.Y(n_8614)
);

INVx1_ASAP7_75t_L g8615 ( 
.A(n_8581),
.Y(n_8615)
);

INVxp67_ASAP7_75t_L g8616 ( 
.A(n_8574),
.Y(n_8616)
);

AOI311xp33_ASAP7_75t_L g8617 ( 
.A1(n_8592),
.A2(n_540),
.A3(n_538),
.B(n_539),
.C(n_541),
.Y(n_8617)
);

AOI211xp5_ASAP7_75t_L g8618 ( 
.A1(n_8583),
.A2(n_8587),
.B(n_8599),
.C(n_8608),
.Y(n_8618)
);

AOI21xp5_ASAP7_75t_L g8619 ( 
.A1(n_8597),
.A2(n_540),
.B(n_541),
.Y(n_8619)
);

NAND2xp5_ASAP7_75t_L g8620 ( 
.A(n_8609),
.B(n_544),
.Y(n_8620)
);

NAND2xp5_ASAP7_75t_L g8621 ( 
.A(n_8578),
.B(n_545),
.Y(n_8621)
);

AOI21xp5_ASAP7_75t_L g8622 ( 
.A1(n_8610),
.A2(n_545),
.B(n_546),
.Y(n_8622)
);

OR2x2_ASAP7_75t_L g8623 ( 
.A(n_8607),
.B(n_549),
.Y(n_8623)
);

AOI22xp5_ASAP7_75t_L g8624 ( 
.A1(n_8586),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.Y(n_8624)
);

INVx1_ASAP7_75t_L g8625 ( 
.A(n_8577),
.Y(n_8625)
);

OAI22xp5_ASAP7_75t_L g8626 ( 
.A1(n_8603),
.A2(n_553),
.B1(n_550),
.B2(n_552),
.Y(n_8626)
);

AOI221xp5_ASAP7_75t_L g8627 ( 
.A1(n_8595),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.C(n_556),
.Y(n_8627)
);

O2A1O1Ixp33_ASAP7_75t_L g8628 ( 
.A1(n_8575),
.A2(n_558),
.B(n_554),
.C(n_557),
.Y(n_8628)
);

OAI221xp5_ASAP7_75t_L g8629 ( 
.A1(n_8590),
.A2(n_561),
.B1(n_557),
.B2(n_559),
.C(n_562),
.Y(n_8629)
);

AOI21xp33_ASAP7_75t_L g8630 ( 
.A1(n_8588),
.A2(n_563),
.B(n_564),
.Y(n_8630)
);

NOR3xp33_ASAP7_75t_L g8631 ( 
.A(n_8589),
.B(n_563),
.C(n_564),
.Y(n_8631)
);

INVx1_ASAP7_75t_L g8632 ( 
.A(n_8596),
.Y(n_8632)
);

OAI21xp33_ASAP7_75t_L g8633 ( 
.A1(n_8604),
.A2(n_566),
.B(n_567),
.Y(n_8633)
);

OAI22xp5_ASAP7_75t_L g8634 ( 
.A1(n_8591),
.A2(n_570),
.B1(n_566),
.B2(n_569),
.Y(n_8634)
);

NAND3xp33_ASAP7_75t_SL g8635 ( 
.A(n_8598),
.B(n_572),
.C(n_573),
.Y(n_8635)
);

AOI221xp5_ASAP7_75t_L g8636 ( 
.A1(n_8605),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.C(n_576),
.Y(n_8636)
);

AOI222xp33_ASAP7_75t_L g8637 ( 
.A1(n_8600),
.A2(n_574),
.B1(n_576),
.B2(n_577),
.C1(n_578),
.C2(n_579),
.Y(n_8637)
);

OAI221xp5_ASAP7_75t_L g8638 ( 
.A1(n_8585),
.A2(n_578),
.B1(n_580),
.B2(n_581),
.C(n_582),
.Y(n_8638)
);

INVx2_ASAP7_75t_L g8639 ( 
.A(n_8601),
.Y(n_8639)
);

AOI31xp33_ASAP7_75t_L g8640 ( 
.A1(n_8582),
.A2(n_585),
.A3(n_583),
.B(n_584),
.Y(n_8640)
);

AOI211xp5_ASAP7_75t_L g8641 ( 
.A1(n_8580),
.A2(n_587),
.B(n_585),
.C(n_586),
.Y(n_8641)
);

O2A1O1Ixp33_ASAP7_75t_L g8642 ( 
.A1(n_8576),
.A2(n_589),
.B(n_587),
.C(n_588),
.Y(n_8642)
);

AOI211xp5_ASAP7_75t_L g8643 ( 
.A1(n_8593),
.A2(n_8602),
.B(n_8579),
.C(n_592),
.Y(n_8643)
);

AOI221x1_ASAP7_75t_L g8644 ( 
.A1(n_8599),
.A2(n_590),
.B1(n_591),
.B2(n_593),
.C(n_594),
.Y(n_8644)
);

OAI222xp33_ASAP7_75t_L g8645 ( 
.A1(n_8606),
.A2(n_591),
.B1(n_593),
.B2(n_594),
.C1(n_595),
.C2(n_596),
.Y(n_8645)
);

AOI221xp5_ASAP7_75t_L g8646 ( 
.A1(n_8616),
.A2(n_598),
.B1(n_599),
.B2(n_600),
.C(n_603),
.Y(n_8646)
);

OAI22xp33_ASAP7_75t_L g8647 ( 
.A1(n_8611),
.A2(n_604),
.B1(n_598),
.B2(n_599),
.Y(n_8647)
);

OAI211xp5_ASAP7_75t_SL g8648 ( 
.A1(n_8618),
.A2(n_608),
.B(n_606),
.C(n_607),
.Y(n_8648)
);

AOI221xp5_ASAP7_75t_L g8649 ( 
.A1(n_8619),
.A2(n_606),
.B1(n_608),
.B2(n_609),
.C(n_610),
.Y(n_8649)
);

OAI21xp5_ASAP7_75t_L g8650 ( 
.A1(n_8615),
.A2(n_609),
.B(n_611),
.Y(n_8650)
);

OAI21xp33_ASAP7_75t_L g8651 ( 
.A1(n_8621),
.A2(n_613),
.B(n_614),
.Y(n_8651)
);

OAI21xp5_ASAP7_75t_SL g8652 ( 
.A1(n_8624),
.A2(n_613),
.B(n_615),
.Y(n_8652)
);

NAND2xp5_ASAP7_75t_SL g8653 ( 
.A(n_8617),
.B(n_1825),
.Y(n_8653)
);

NAND2xp5_ASAP7_75t_L g8654 ( 
.A(n_8632),
.B(n_616),
.Y(n_8654)
);

AOI21xp5_ASAP7_75t_L g8655 ( 
.A1(n_8613),
.A2(n_616),
.B(n_617),
.Y(n_8655)
);

NAND2xp5_ASAP7_75t_L g8656 ( 
.A(n_8644),
.B(n_617),
.Y(n_8656)
);

NAND2xp5_ASAP7_75t_SL g8657 ( 
.A(n_8637),
.B(n_1878),
.Y(n_8657)
);

O2A1O1Ixp33_ASAP7_75t_L g8658 ( 
.A1(n_8639),
.A2(n_620),
.B(n_618),
.C(n_619),
.Y(n_8658)
);

NAND2xp5_ASAP7_75t_L g8659 ( 
.A(n_8625),
.B(n_619),
.Y(n_8659)
);

AOI221xp5_ASAP7_75t_L g8660 ( 
.A1(n_8636),
.A2(n_620),
.B1(n_621),
.B2(n_623),
.C(n_624),
.Y(n_8660)
);

AOI21xp33_ASAP7_75t_SL g8661 ( 
.A1(n_8640),
.A2(n_625),
.B(n_626),
.Y(n_8661)
);

NAND2xp5_ASAP7_75t_L g8662 ( 
.A(n_8623),
.B(n_626),
.Y(n_8662)
);

OAI21xp5_ASAP7_75t_L g8663 ( 
.A1(n_8622),
.A2(n_628),
.B(n_630),
.Y(n_8663)
);

AOI22xp5_ASAP7_75t_L g8664 ( 
.A1(n_8634),
.A2(n_632),
.B1(n_628),
.B2(n_631),
.Y(n_8664)
);

AOI22xp5_ASAP7_75t_L g8665 ( 
.A1(n_8635),
.A2(n_634),
.B1(n_631),
.B2(n_633),
.Y(n_8665)
);

OAI321xp33_ASAP7_75t_L g8666 ( 
.A1(n_8643),
.A2(n_633),
.A3(n_636),
.B1(n_637),
.B2(n_638),
.C(n_639),
.Y(n_8666)
);

AOI22x1_ASAP7_75t_L g8667 ( 
.A1(n_8641),
.A2(n_638),
.B1(n_636),
.B2(n_637),
.Y(n_8667)
);

NAND2xp5_ASAP7_75t_L g8668 ( 
.A(n_8631),
.B(n_640),
.Y(n_8668)
);

AOI222xp33_ASAP7_75t_L g8669 ( 
.A1(n_8627),
.A2(n_641),
.B1(n_642),
.B2(n_643),
.C1(n_645),
.C2(n_646),
.Y(n_8669)
);

OAI221xp5_ASAP7_75t_L g8670 ( 
.A1(n_8633),
.A2(n_641),
.B1(n_645),
.B2(n_646),
.C(n_647),
.Y(n_8670)
);

OAI21xp33_ASAP7_75t_L g8671 ( 
.A1(n_8629),
.A2(n_648),
.B(n_649),
.Y(n_8671)
);

AOI22xp5_ASAP7_75t_L g8672 ( 
.A1(n_8620),
.A2(n_651),
.B1(n_648),
.B2(n_650),
.Y(n_8672)
);

AOI221xp5_ASAP7_75t_L g8673 ( 
.A1(n_8630),
.A2(n_652),
.B1(n_653),
.B2(n_654),
.C(n_655),
.Y(n_8673)
);

AOI311xp33_ASAP7_75t_L g8674 ( 
.A1(n_8638),
.A2(n_652),
.A3(n_653),
.B(n_657),
.C(n_658),
.Y(n_8674)
);

AOI21xp5_ASAP7_75t_L g8675 ( 
.A1(n_8628),
.A2(n_657),
.B(n_660),
.Y(n_8675)
);

AOI21xp5_ASAP7_75t_L g8676 ( 
.A1(n_8645),
.A2(n_661),
.B(n_662),
.Y(n_8676)
);

AOI22xp5_ASAP7_75t_L g8677 ( 
.A1(n_8612),
.A2(n_661),
.B1(n_665),
.B2(n_667),
.Y(n_8677)
);

AOI21xp5_ASAP7_75t_L g8678 ( 
.A1(n_8626),
.A2(n_667),
.B(n_668),
.Y(n_8678)
);

OAI221xp5_ASAP7_75t_L g8679 ( 
.A1(n_8649),
.A2(n_8642),
.B1(n_8614),
.B2(n_671),
.C(n_672),
.Y(n_8679)
);

NAND3xp33_ASAP7_75t_L g8680 ( 
.A(n_8653),
.B(n_1949),
.C(n_1878),
.Y(n_8680)
);

AOI21xp33_ASAP7_75t_SL g8681 ( 
.A1(n_8656),
.A2(n_8647),
.B(n_8662),
.Y(n_8681)
);

NOR2xp33_ASAP7_75t_L g8682 ( 
.A(n_8661),
.B(n_8648),
.Y(n_8682)
);

AOI221xp5_ASAP7_75t_L g8683 ( 
.A1(n_8651),
.A2(n_669),
.B1(n_670),
.B2(n_671),
.C(n_672),
.Y(n_8683)
);

O2A1O1Ixp33_ASAP7_75t_L g8684 ( 
.A1(n_8659),
.A2(n_673),
.B(n_674),
.C(n_675),
.Y(n_8684)
);

OAI21xp33_ASAP7_75t_SL g8685 ( 
.A1(n_8663),
.A2(n_674),
.B(n_675),
.Y(n_8685)
);

AOI221xp5_ASAP7_75t_L g8686 ( 
.A1(n_8676),
.A2(n_676),
.B1(n_677),
.B2(n_679),
.C(n_680),
.Y(n_8686)
);

NOR3x1_ASAP7_75t_L g8687 ( 
.A(n_8650),
.B(n_8670),
.C(n_8652),
.Y(n_8687)
);

HB1xp67_ASAP7_75t_L g8688 ( 
.A(n_8654),
.Y(n_8688)
);

OAI21xp5_ASAP7_75t_SL g8689 ( 
.A1(n_8665),
.A2(n_676),
.B(n_680),
.Y(n_8689)
);

NAND2xp5_ASAP7_75t_SL g8690 ( 
.A(n_8666),
.B(n_1878),
.Y(n_8690)
);

O2A1O1Ixp5_ASAP7_75t_L g8691 ( 
.A1(n_8655),
.A2(n_681),
.B(n_682),
.C(n_683),
.Y(n_8691)
);

NAND3x1_ASAP7_75t_L g8692 ( 
.A(n_8668),
.B(n_681),
.C(n_682),
.Y(n_8692)
);

AOI221xp5_ASAP7_75t_L g8693 ( 
.A1(n_8658),
.A2(n_685),
.B1(n_686),
.B2(n_687),
.C(n_688),
.Y(n_8693)
);

AOI31xp33_ASAP7_75t_L g8694 ( 
.A1(n_8673),
.A2(n_689),
.A3(n_690),
.B(n_691),
.Y(n_8694)
);

NAND2xp5_ASAP7_75t_SL g8695 ( 
.A(n_8674),
.B(n_1949),
.Y(n_8695)
);

AOI21xp5_ASAP7_75t_L g8696 ( 
.A1(n_8657),
.A2(n_689),
.B(n_691),
.Y(n_8696)
);

AOI21xp33_ASAP7_75t_SL g8697 ( 
.A1(n_8667),
.A2(n_692),
.B(n_693),
.Y(n_8697)
);

NAND2xp5_ASAP7_75t_L g8698 ( 
.A(n_8675),
.B(n_692),
.Y(n_8698)
);

NAND4xp25_ASAP7_75t_SL g8699 ( 
.A(n_8669),
.B(n_693),
.C(n_695),
.D(n_697),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8672),
.Y(n_8700)
);

AOI221x1_ASAP7_75t_L g8701 ( 
.A1(n_8671),
.A2(n_695),
.B1(n_698),
.B2(n_699),
.C(n_700),
.Y(n_8701)
);

AOI211xp5_ASAP7_75t_L g8702 ( 
.A1(n_8660),
.A2(n_8678),
.B(n_8646),
.C(n_8677),
.Y(n_8702)
);

OAI22xp5_ASAP7_75t_L g8703 ( 
.A1(n_8664),
.A2(n_701),
.B1(n_702),
.B2(n_703),
.Y(n_8703)
);

OAI22xp33_ASAP7_75t_L g8704 ( 
.A1(n_8677),
.A2(n_702),
.B1(n_703),
.B2(n_705),
.Y(n_8704)
);

AOI222xp33_ASAP7_75t_L g8705 ( 
.A1(n_8656),
.A2(n_705),
.B1(n_706),
.B2(n_707),
.C1(n_708),
.C2(n_709),
.Y(n_8705)
);

OAI21xp33_ASAP7_75t_L g8706 ( 
.A1(n_8682),
.A2(n_706),
.B(n_707),
.Y(n_8706)
);

O2A1O1Ixp33_ASAP7_75t_L g8707 ( 
.A1(n_8681),
.A2(n_708),
.B(n_710),
.C(n_711),
.Y(n_8707)
);

NAND2xp5_ASAP7_75t_L g8708 ( 
.A(n_8688),
.B(n_711),
.Y(n_8708)
);

AOI31xp33_ASAP7_75t_L g8709 ( 
.A1(n_8705),
.A2(n_712),
.A3(n_713),
.B(n_714),
.Y(n_8709)
);

NAND3xp33_ASAP7_75t_L g8710 ( 
.A(n_8695),
.B(n_1977),
.C(n_1949),
.Y(n_8710)
);

INVx1_ASAP7_75t_L g8711 ( 
.A(n_8692),
.Y(n_8711)
);

NOR2xp33_ASAP7_75t_L g8712 ( 
.A(n_8685),
.B(n_715),
.Y(n_8712)
);

INVx2_ASAP7_75t_L g8713 ( 
.A(n_8691),
.Y(n_8713)
);

OR2x2_ASAP7_75t_L g8714 ( 
.A(n_8698),
.B(n_715),
.Y(n_8714)
);

INVxp67_ASAP7_75t_L g8715 ( 
.A(n_8690),
.Y(n_8715)
);

AOI211xp5_ASAP7_75t_L g8716 ( 
.A1(n_8704),
.A2(n_716),
.B(n_718),
.C(n_719),
.Y(n_8716)
);

NAND3xp33_ASAP7_75t_L g8717 ( 
.A(n_8700),
.B(n_1977),
.C(n_1949),
.Y(n_8717)
);

BUFx2_ASAP7_75t_L g8718 ( 
.A(n_8686),
.Y(n_8718)
);

NOR3x1_ASAP7_75t_L g8719 ( 
.A(n_8689),
.B(n_718),
.C(n_719),
.Y(n_8719)
);

INVx1_ASAP7_75t_L g8720 ( 
.A(n_8684),
.Y(n_8720)
);

AOI21xp5_ASAP7_75t_L g8721 ( 
.A1(n_8696),
.A2(n_720),
.B(n_721),
.Y(n_8721)
);

NAND2xp5_ASAP7_75t_L g8722 ( 
.A(n_8697),
.B(n_720),
.Y(n_8722)
);

NOR2x1p5_ASAP7_75t_SL g8723 ( 
.A(n_8687),
.B(n_721),
.Y(n_8723)
);

INVx1_ASAP7_75t_L g8724 ( 
.A(n_8694),
.Y(n_8724)
);

NAND3xp33_ASAP7_75t_L g8725 ( 
.A(n_8683),
.B(n_8693),
.C(n_8701),
.Y(n_8725)
);

NAND4xp25_ASAP7_75t_L g8726 ( 
.A(n_8702),
.B(n_722),
.C(n_724),
.D(n_725),
.Y(n_8726)
);

NAND2xp5_ASAP7_75t_L g8727 ( 
.A(n_8703),
.B(n_724),
.Y(n_8727)
);

NOR3xp33_ASAP7_75t_L g8728 ( 
.A(n_8680),
.B(n_726),
.C(n_727),
.Y(n_8728)
);

NAND4xp25_ASAP7_75t_L g8729 ( 
.A(n_8679),
.B(n_726),
.C(n_728),
.D(n_732),
.Y(n_8729)
);

NAND2xp5_ASAP7_75t_L g8730 ( 
.A(n_8699),
.B(n_732),
.Y(n_8730)
);

NOR2xp67_ASAP7_75t_L g8731 ( 
.A(n_8726),
.B(n_733),
.Y(n_8731)
);

NOR2xp33_ASAP7_75t_L g8732 ( 
.A(n_8711),
.B(n_733),
.Y(n_8732)
);

NOR3x1_ASAP7_75t_L g8733 ( 
.A(n_8722),
.B(n_734),
.C(n_735),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_8723),
.Y(n_8734)
);

NAND3xp33_ASAP7_75t_L g8735 ( 
.A(n_8720),
.B(n_1977),
.C(n_2666),
.Y(n_8735)
);

NOR3xp33_ASAP7_75t_SL g8736 ( 
.A(n_8729),
.B(n_734),
.C(n_736),
.Y(n_8736)
);

AOI21xp5_ASAP7_75t_L g8737 ( 
.A1(n_8730),
.A2(n_1977),
.B(n_737),
.Y(n_8737)
);

INVx1_ASAP7_75t_L g8738 ( 
.A(n_8713),
.Y(n_8738)
);

NAND3xp33_ASAP7_75t_L g8739 ( 
.A(n_8724),
.B(n_2666),
.C(n_738),
.Y(n_8739)
);

OR2x2_ASAP7_75t_L g8740 ( 
.A(n_8714),
.B(n_736),
.Y(n_8740)
);

NAND4xp25_ASAP7_75t_L g8741 ( 
.A(n_8719),
.B(n_738),
.C(n_739),
.D(n_740),
.Y(n_8741)
);

NAND4xp25_ASAP7_75t_L g8742 ( 
.A(n_8712),
.B(n_739),
.C(n_740),
.D(n_741),
.Y(n_8742)
);

NAND2xp5_ASAP7_75t_L g8743 ( 
.A(n_8709),
.B(n_742),
.Y(n_8743)
);

NAND2xp5_ASAP7_75t_L g8744 ( 
.A(n_8708),
.B(n_743),
.Y(n_8744)
);

NAND4xp75_ASAP7_75t_L g8745 ( 
.A(n_8721),
.B(n_743),
.C(n_744),
.D(n_745),
.Y(n_8745)
);

NAND3xp33_ASAP7_75t_L g8746 ( 
.A(n_8715),
.B(n_2666),
.C(n_745),
.Y(n_8746)
);

NAND3xp33_ASAP7_75t_L g8747 ( 
.A(n_8718),
.B(n_2666),
.C(n_746),
.Y(n_8747)
);

OAI22xp5_ASAP7_75t_SL g8748 ( 
.A1(n_8727),
.A2(n_744),
.B1(n_746),
.B2(n_747),
.Y(n_8748)
);

HB1xp67_ASAP7_75t_L g8749 ( 
.A(n_8725),
.Y(n_8749)
);

NAND4xp25_ASAP7_75t_L g8750 ( 
.A(n_8707),
.B(n_748),
.C(n_751),
.D(n_752),
.Y(n_8750)
);

AOI211xp5_ASAP7_75t_L g8751 ( 
.A1(n_8706),
.A2(n_748),
.B(n_751),
.C(n_752),
.Y(n_8751)
);

NOR3xp33_ASAP7_75t_L g8752 ( 
.A(n_8710),
.B(n_753),
.C(n_754),
.Y(n_8752)
);

NOR2xp67_ASAP7_75t_L g8753 ( 
.A(n_8717),
.B(n_754),
.Y(n_8753)
);

NOR2xp67_ASAP7_75t_L g8754 ( 
.A(n_8716),
.B(n_755),
.Y(n_8754)
);

NAND4xp75_ASAP7_75t_L g8755 ( 
.A(n_8728),
.B(n_755),
.C(n_756),
.D(n_757),
.Y(n_8755)
);

NAND2xp5_ASAP7_75t_L g8756 ( 
.A(n_8711),
.B(n_756),
.Y(n_8756)
);

INVx1_ASAP7_75t_L g8757 ( 
.A(n_8723),
.Y(n_8757)
);

NOR2x1_ASAP7_75t_L g8758 ( 
.A(n_8711),
.B(n_757),
.Y(n_8758)
);

NOR2x1p5_ASAP7_75t_SL g8759 ( 
.A(n_8714),
.B(n_758),
.Y(n_8759)
);

NOR3xp33_ASAP7_75t_L g8760 ( 
.A(n_8738),
.B(n_759),
.C(n_760),
.Y(n_8760)
);

AND2x2_ASAP7_75t_SL g8761 ( 
.A(n_8749),
.B(n_759),
.Y(n_8761)
);

INVx1_ASAP7_75t_L g8762 ( 
.A(n_8759),
.Y(n_8762)
);

INVx1_ASAP7_75t_L g8763 ( 
.A(n_8734),
.Y(n_8763)
);

INVxp67_ASAP7_75t_L g8764 ( 
.A(n_8757),
.Y(n_8764)
);

INVx1_ASAP7_75t_L g8765 ( 
.A(n_8758),
.Y(n_8765)
);

INVx3_ASAP7_75t_SL g8766 ( 
.A(n_8740),
.Y(n_8766)
);

INVxp67_ASAP7_75t_SL g8767 ( 
.A(n_8756),
.Y(n_8767)
);

NAND2xp5_ASAP7_75t_L g8768 ( 
.A(n_8731),
.B(n_761),
.Y(n_8768)
);

NAND2xp5_ASAP7_75t_L g8769 ( 
.A(n_8733),
.B(n_761),
.Y(n_8769)
);

HB1xp67_ASAP7_75t_L g8770 ( 
.A(n_8744),
.Y(n_8770)
);

NAND2xp33_ASAP7_75t_SL g8771 ( 
.A(n_8748),
.B(n_762),
.Y(n_8771)
);

NAND2xp5_ASAP7_75t_L g8772 ( 
.A(n_8754),
.B(n_763),
.Y(n_8772)
);

INVx1_ASAP7_75t_L g8773 ( 
.A(n_8743),
.Y(n_8773)
);

INVx1_ASAP7_75t_L g8774 ( 
.A(n_8732),
.Y(n_8774)
);

INVx1_ASAP7_75t_L g8775 ( 
.A(n_8742),
.Y(n_8775)
);

OR2x2_ASAP7_75t_L g8776 ( 
.A(n_8741),
.B(n_764),
.Y(n_8776)
);

NAND2xp5_ASAP7_75t_L g8777 ( 
.A(n_8736),
.B(n_764),
.Y(n_8777)
);

NAND2xp5_ASAP7_75t_SL g8778 ( 
.A(n_8751),
.B(n_765),
.Y(n_8778)
);

NAND2xp5_ASAP7_75t_SL g8779 ( 
.A(n_8753),
.B(n_765),
.Y(n_8779)
);

AOI21xp33_ASAP7_75t_L g8780 ( 
.A1(n_8747),
.A2(n_766),
.B(n_767),
.Y(n_8780)
);

NAND2xp5_ASAP7_75t_L g8781 ( 
.A(n_8737),
.B(n_766),
.Y(n_8781)
);

NAND2xp5_ASAP7_75t_L g8782 ( 
.A(n_8745),
.B(n_768),
.Y(n_8782)
);

OR2x2_ASAP7_75t_L g8783 ( 
.A(n_8750),
.B(n_770),
.Y(n_8783)
);

NOR2xp67_ASAP7_75t_L g8784 ( 
.A(n_8739),
.B(n_770),
.Y(n_8784)
);

HB1xp67_ASAP7_75t_L g8785 ( 
.A(n_8762),
.Y(n_8785)
);

NOR3xp33_ASAP7_75t_L g8786 ( 
.A(n_8764),
.B(n_8755),
.C(n_8746),
.Y(n_8786)
);

NAND3xp33_ASAP7_75t_L g8787 ( 
.A(n_8765),
.B(n_8763),
.C(n_8770),
.Y(n_8787)
);

AOI211x1_ASAP7_75t_L g8788 ( 
.A1(n_8769),
.A2(n_8735),
.B(n_8752),
.C(n_773),
.Y(n_8788)
);

NAND2xp5_ASAP7_75t_L g8789 ( 
.A(n_8766),
.B(n_771),
.Y(n_8789)
);

AOI211xp5_ASAP7_75t_L g8790 ( 
.A1(n_8768),
.A2(n_8767),
.B(n_8772),
.C(n_8774),
.Y(n_8790)
);

AND2x2_ASAP7_75t_L g8791 ( 
.A(n_8761),
.B(n_772),
.Y(n_8791)
);

INVx1_ASAP7_75t_L g8792 ( 
.A(n_8777),
.Y(n_8792)
);

INVx1_ASAP7_75t_L g8793 ( 
.A(n_8779),
.Y(n_8793)
);

NAND3xp33_ASAP7_75t_SL g8794 ( 
.A(n_8773),
.B(n_772),
.C(n_774),
.Y(n_8794)
);

NOR2xp67_ASAP7_75t_L g8795 ( 
.A(n_8776),
.B(n_774),
.Y(n_8795)
);

OR2x2_ASAP7_75t_L g8796 ( 
.A(n_8783),
.B(n_775),
.Y(n_8796)
);

NAND2xp5_ASAP7_75t_L g8797 ( 
.A(n_8784),
.B(n_775),
.Y(n_8797)
);

NAND4xp75_ASAP7_75t_L g8798 ( 
.A(n_8775),
.B(n_776),
.C(n_777),
.D(n_778),
.Y(n_8798)
);

NAND3xp33_ASAP7_75t_SL g8799 ( 
.A(n_8760),
.B(n_777),
.C(n_779),
.Y(n_8799)
);

NOR2x1_ASAP7_75t_L g8800 ( 
.A(n_8782),
.B(n_781),
.Y(n_8800)
);

NOR3xp33_ASAP7_75t_L g8801 ( 
.A(n_8771),
.B(n_781),
.C(n_783),
.Y(n_8801)
);

NAND4xp25_ASAP7_75t_L g8802 ( 
.A(n_8781),
.B(n_785),
.C(n_787),
.D(n_789),
.Y(n_8802)
);

AOI22xp5_ASAP7_75t_L g8803 ( 
.A1(n_8787),
.A2(n_8778),
.B1(n_8780),
.B2(n_793),
.Y(n_8803)
);

AND2x2_ASAP7_75t_L g8804 ( 
.A(n_8785),
.B(n_790),
.Y(n_8804)
);

INVx1_ASAP7_75t_L g8805 ( 
.A(n_8791),
.Y(n_8805)
);

AOI22xp5_ASAP7_75t_L g8806 ( 
.A1(n_8795),
.A2(n_790),
.B1(n_791),
.B2(n_794),
.Y(n_8806)
);

NAND2xp5_ASAP7_75t_SL g8807 ( 
.A(n_8790),
.B(n_791),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_8797),
.Y(n_8808)
);

INVx1_ASAP7_75t_L g8809 ( 
.A(n_8789),
.Y(n_8809)
);

NAND2xp33_ASAP7_75t_SL g8810 ( 
.A(n_8804),
.B(n_8796),
.Y(n_8810)
);

INVx1_ASAP7_75t_L g8811 ( 
.A(n_8805),
.Y(n_8811)
);

AOI211xp5_ASAP7_75t_L g8812 ( 
.A1(n_8808),
.A2(n_8793),
.B(n_8786),
.C(n_8792),
.Y(n_8812)
);

NOR3xp33_ASAP7_75t_SL g8813 ( 
.A(n_8809),
.B(n_8799),
.C(n_8794),
.Y(n_8813)
);

AND2x2_ASAP7_75t_L g8814 ( 
.A(n_8806),
.B(n_8800),
.Y(n_8814)
);

OA211x2_ASAP7_75t_L g8815 ( 
.A1(n_8810),
.A2(n_8807),
.B(n_8801),
.C(n_8802),
.Y(n_8815)
);

OAI211xp5_ASAP7_75t_SL g8816 ( 
.A1(n_8812),
.A2(n_8803),
.B(n_8788),
.C(n_8798),
.Y(n_8816)
);

AOI22xp33_ASAP7_75t_L g8817 ( 
.A1(n_8811),
.A2(n_795),
.B1(n_796),
.B2(n_797),
.Y(n_8817)
);

AOI21xp5_ASAP7_75t_L g8818 ( 
.A1(n_8814),
.A2(n_2666),
.B(n_798),
.Y(n_8818)
);

AND4x1_ASAP7_75t_L g8819 ( 
.A(n_8813),
.B(n_796),
.C(n_798),
.D(n_799),
.Y(n_8819)
);

NAND2xp5_ASAP7_75t_L g8820 ( 
.A(n_8811),
.B(n_800),
.Y(n_8820)
);

NAND3x1_ASAP7_75t_SL g8821 ( 
.A(n_8814),
.B(n_800),
.C(n_801),
.Y(n_8821)
);

NOR2x1_ASAP7_75t_L g8822 ( 
.A(n_8811),
.B(n_801),
.Y(n_8822)
);

AOI222xp33_ASAP7_75t_L g8823 ( 
.A1(n_8811),
.A2(n_802),
.B1(n_804),
.B2(n_805),
.C1(n_806),
.C2(n_807),
.Y(n_8823)
);

OR2x2_ASAP7_75t_L g8824 ( 
.A(n_8811),
.B(n_802),
.Y(n_8824)
);

INVx2_ASAP7_75t_L g8825 ( 
.A(n_8824),
.Y(n_8825)
);

INVx3_ASAP7_75t_L g8826 ( 
.A(n_8819),
.Y(n_8826)
);

NAND2xp5_ASAP7_75t_L g8827 ( 
.A(n_8822),
.B(n_8820),
.Y(n_8827)
);

INVx3_ASAP7_75t_L g8828 ( 
.A(n_8816),
.Y(n_8828)
);

INVx2_ASAP7_75t_L g8829 ( 
.A(n_8815),
.Y(n_8829)
);

NAND3x1_ASAP7_75t_L g8830 ( 
.A(n_8818),
.B(n_805),
.C(n_806),
.Y(n_8830)
);

NOR2x1_ASAP7_75t_L g8831 ( 
.A(n_8821),
.B(n_807),
.Y(n_8831)
);

NOR3xp33_ASAP7_75t_L g8832 ( 
.A(n_8823),
.B(n_809),
.C(n_810),
.Y(n_8832)
);

INVx1_ASAP7_75t_L g8833 ( 
.A(n_8817),
.Y(n_8833)
);

INVx1_ASAP7_75t_L g8834 ( 
.A(n_8822),
.Y(n_8834)
);

INVx2_ASAP7_75t_L g8835 ( 
.A(n_8824),
.Y(n_8835)
);

INVxp67_ASAP7_75t_SL g8836 ( 
.A(n_8822),
.Y(n_8836)
);

BUFx3_ASAP7_75t_L g8837 ( 
.A(n_8824),
.Y(n_8837)
);

INVx2_ASAP7_75t_L g8838 ( 
.A(n_8824),
.Y(n_8838)
);

NAND3xp33_ASAP7_75t_L g8839 ( 
.A(n_8829),
.B(n_2439),
.C(n_811),
.Y(n_8839)
);

OAI22xp33_ASAP7_75t_L g8840 ( 
.A1(n_8828),
.A2(n_809),
.B1(n_811),
.B2(n_813),
.Y(n_8840)
);

NOR3xp33_ASAP7_75t_L g8841 ( 
.A(n_8836),
.B(n_813),
.C(n_814),
.Y(n_8841)
);

AOI322xp5_ASAP7_75t_L g8842 ( 
.A1(n_8834),
.A2(n_8831),
.A3(n_8838),
.B1(n_8835),
.B2(n_8825),
.C1(n_8827),
.C2(n_8832),
.Y(n_8842)
);

NAND2xp5_ASAP7_75t_L g8843 ( 
.A(n_8837),
.B(n_814),
.Y(n_8843)
);

AOI22xp5_ASAP7_75t_L g8844 ( 
.A1(n_8826),
.A2(n_2678),
.B1(n_2590),
.B2(n_2584),
.Y(n_8844)
);

INVx1_ASAP7_75t_L g8845 ( 
.A(n_8843),
.Y(n_8845)
);

OAI31xp33_ASAP7_75t_L g8846 ( 
.A1(n_8840),
.A2(n_8833),
.A3(n_8830),
.B(n_817),
.Y(n_8846)
);

INVx1_ASAP7_75t_L g8847 ( 
.A(n_8841),
.Y(n_8847)
);

INVx1_ASAP7_75t_L g8848 ( 
.A(n_8839),
.Y(n_8848)
);

INVx1_ASAP7_75t_L g8849 ( 
.A(n_8842),
.Y(n_8849)
);

OAI22xp5_ASAP7_75t_SL g8850 ( 
.A1(n_8849),
.A2(n_8844),
.B1(n_816),
.B2(n_817),
.Y(n_8850)
);

XNOR2xp5_ASAP7_75t_SL g8851 ( 
.A(n_8847),
.B(n_815),
.Y(n_8851)
);

INVx1_ASAP7_75t_L g8852 ( 
.A(n_8845),
.Y(n_8852)
);

XNOR2x1_ASAP7_75t_L g8853 ( 
.A(n_8848),
.B(n_8846),
.Y(n_8853)
);

NOR2xp33_ASAP7_75t_L g8854 ( 
.A(n_8849),
.B(n_815),
.Y(n_8854)
);

INVx2_ASAP7_75t_L g8855 ( 
.A(n_8849),
.Y(n_8855)
);

OAI22xp5_ASAP7_75t_L g8856 ( 
.A1(n_8849),
.A2(n_2678),
.B1(n_2590),
.B2(n_2584),
.Y(n_8856)
);

INVx2_ASAP7_75t_L g8857 ( 
.A(n_8849),
.Y(n_8857)
);

INVx3_ASAP7_75t_SL g8858 ( 
.A(n_8849),
.Y(n_8858)
);

AOI22xp5_ASAP7_75t_L g8859 ( 
.A1(n_8849),
.A2(n_2678),
.B1(n_2590),
.B2(n_2584),
.Y(n_8859)
);

XOR2xp5_ASAP7_75t_L g8860 ( 
.A(n_8849),
.B(n_818),
.Y(n_8860)
);

OAI22xp5_ASAP7_75t_L g8861 ( 
.A1(n_8849),
.A2(n_2678),
.B1(n_2590),
.B2(n_2705),
.Y(n_8861)
);

INVx2_ASAP7_75t_SL g8862 ( 
.A(n_8849),
.Y(n_8862)
);

INVx1_ASAP7_75t_L g8863 ( 
.A(n_8849),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_8855),
.Y(n_8864)
);

NAND3xp33_ASAP7_75t_L g8865 ( 
.A(n_8863),
.B(n_818),
.C(n_819),
.Y(n_8865)
);

AOI22xp33_ASAP7_75t_L g8866 ( 
.A1(n_8862),
.A2(n_820),
.B1(n_821),
.B2(n_822),
.Y(n_8866)
);

OAI22xp5_ASAP7_75t_L g8867 ( 
.A1(n_8857),
.A2(n_2705),
.B1(n_825),
.B2(n_826),
.Y(n_8867)
);

OAI21xp5_ASAP7_75t_L g8868 ( 
.A1(n_8852),
.A2(n_824),
.B(n_825),
.Y(n_8868)
);

AOI21xp5_ASAP7_75t_L g8869 ( 
.A1(n_8853),
.A2(n_826),
.B(n_827),
.Y(n_8869)
);

INVx2_ASAP7_75t_L g8870 ( 
.A(n_8858),
.Y(n_8870)
);

OAI31xp33_ASAP7_75t_L g8871 ( 
.A1(n_8860),
.A2(n_827),
.A3(n_828),
.B(n_829),
.Y(n_8871)
);

AOI21x1_ASAP7_75t_L g8872 ( 
.A1(n_8851),
.A2(n_8854),
.B(n_8850),
.Y(n_8872)
);

CKINVDCx20_ASAP7_75t_R g8873 ( 
.A(n_8870),
.Y(n_8873)
);

OAI221xp5_ASAP7_75t_L g8874 ( 
.A1(n_8864),
.A2(n_8859),
.B1(n_8861),
.B2(n_8856),
.C(n_833),
.Y(n_8874)
);

INVx2_ASAP7_75t_L g8875 ( 
.A(n_8872),
.Y(n_8875)
);

OR2x2_ASAP7_75t_L g8876 ( 
.A(n_8865),
.B(n_828),
.Y(n_8876)
);

AOI22xp5_ASAP7_75t_L g8877 ( 
.A1(n_8868),
.A2(n_2705),
.B1(n_832),
.B2(n_835),
.Y(n_8877)
);

BUFx2_ASAP7_75t_SL g8878 ( 
.A(n_8869),
.Y(n_8878)
);

INVx1_ASAP7_75t_L g8879 ( 
.A(n_8866),
.Y(n_8879)
);

AOI21xp5_ASAP7_75t_L g8880 ( 
.A1(n_8873),
.A2(n_8871),
.B(n_8867),
.Y(n_8880)
);

AOI21xp33_ASAP7_75t_L g8881 ( 
.A1(n_8875),
.A2(n_829),
.B(n_832),
.Y(n_8881)
);

INVx1_ASAP7_75t_L g8882 ( 
.A(n_8878),
.Y(n_8882)
);

NAND2xp5_ASAP7_75t_L g8883 ( 
.A(n_8879),
.B(n_836),
.Y(n_8883)
);

AOI21xp5_ASAP7_75t_L g8884 ( 
.A1(n_8874),
.A2(n_836),
.B(n_837),
.Y(n_8884)
);

INVx1_ASAP7_75t_L g8885 ( 
.A(n_8882),
.Y(n_8885)
);

INVxp67_ASAP7_75t_L g8886 ( 
.A(n_8880),
.Y(n_8886)
);

AOI22xp5_ASAP7_75t_L g8887 ( 
.A1(n_8883),
.A2(n_8876),
.B1(n_8877),
.B2(n_2705),
.Y(n_8887)
);

XNOR2xp5_ASAP7_75t_L g8888 ( 
.A(n_8885),
.B(n_8884),
.Y(n_8888)
);

OA21x2_ASAP7_75t_L g8889 ( 
.A1(n_8886),
.A2(n_8881),
.B(n_839),
.Y(n_8889)
);

OAI22xp33_ASAP7_75t_SL g8890 ( 
.A1(n_8887),
.A2(n_838),
.B1(n_839),
.B2(n_840),
.Y(n_8890)
);

OAI22xp5_ASAP7_75t_L g8891 ( 
.A1(n_8888),
.A2(n_838),
.B1(n_840),
.B2(n_841),
.Y(n_8891)
);

OAI22xp5_ASAP7_75t_L g8892 ( 
.A1(n_8889),
.A2(n_842),
.B1(n_843),
.B2(n_844),
.Y(n_8892)
);

AOI31xp33_ASAP7_75t_L g8893 ( 
.A1(n_8890),
.A2(n_843),
.A3(n_845),
.B(n_846),
.Y(n_8893)
);

OAI21xp5_ASAP7_75t_L g8894 ( 
.A1(n_8892),
.A2(n_845),
.B(n_846),
.Y(n_8894)
);

OAI22xp5_ASAP7_75t_L g8895 ( 
.A1(n_8893),
.A2(n_847),
.B1(n_2439),
.B2(n_3358),
.Y(n_8895)
);

INVx1_ASAP7_75t_L g8896 ( 
.A(n_8891),
.Y(n_8896)
);

OAI21xp5_ASAP7_75t_L g8897 ( 
.A1(n_8892),
.A2(n_847),
.B(n_1530),
.Y(n_8897)
);

XNOR2xp5_ASAP7_75t_L g8898 ( 
.A(n_8896),
.B(n_1608),
.Y(n_8898)
);

INVx2_ASAP7_75t_L g8899 ( 
.A(n_8897),
.Y(n_8899)
);

INVx1_ASAP7_75t_L g8900 ( 
.A(n_8894),
.Y(n_8900)
);

NAND2xp5_ASAP7_75t_L g8901 ( 
.A(n_8898),
.B(n_8899),
.Y(n_8901)
);

OA21x2_ASAP7_75t_L g8902 ( 
.A1(n_8900),
.A2(n_8895),
.B(n_1612),
.Y(n_8902)
);

OR2x6_ASAP7_75t_L g8903 ( 
.A(n_8899),
.B(n_2439),
.Y(n_8903)
);

OAI22xp5_ASAP7_75t_SL g8904 ( 
.A1(n_8901),
.A2(n_8902),
.B1(n_8903),
.B2(n_1651),
.Y(n_8904)
);

AOI22xp33_ASAP7_75t_L g8905 ( 
.A1(n_8904),
.A2(n_1724),
.B1(n_2439),
.B2(n_3358),
.Y(n_8905)
);

AOI211xp5_ASAP7_75t_L g8906 ( 
.A1(n_8905),
.A2(n_3358),
.B(n_3345),
.C(n_3335),
.Y(n_8906)
);


endmodule