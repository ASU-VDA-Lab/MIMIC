module real_aes_1823_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_0), .B(n_497), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_1), .A2(n_499), .B(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_2), .B(n_798), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g105 ( .A1(n_3), .A2(n_4), .B1(n_106), .B2(n_107), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_3), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_4), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_5), .B(n_208), .Y(n_534) );
INVx1_ASAP7_75t_L g140 ( .A(n_6), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_7), .B(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_8), .B(n_208), .Y(n_583) );
INVx1_ASAP7_75t_L g178 ( .A(n_9), .Y(n_178) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_10), .A2(n_104), .B1(n_105), .B2(n_108), .C1(n_785), .C2(n_789), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g798 ( .A(n_11), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_12), .Y(n_146) );
NAND2xp33_ASAP7_75t_L g575 ( .A(n_13), .B(n_205), .Y(n_575) );
INVx2_ASAP7_75t_L g122 ( .A(n_14), .Y(n_122) );
AOI221x1_ASAP7_75t_L g519 ( .A1(n_15), .A2(n_28), .B1(n_497), .B2(n_499), .C(n_520), .Y(n_519) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_16), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_17), .B(n_497), .Y(n_571) );
INVx1_ASAP7_75t_L g206 ( .A(n_18), .Y(n_206) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_19), .A2(n_175), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_20), .B(n_170), .Y(n_523) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_21), .A2(n_101), .B1(n_791), .B2(n_802), .C1(n_813), .C2(n_815), .Y(n_100) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_21), .A2(n_80), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_21), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_22), .B(n_208), .Y(n_508) );
AO21x1_ASAP7_75t_L g529 ( .A1(n_23), .A2(n_497), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g484 ( .A(n_24), .Y(n_484) );
INVx1_ASAP7_75t_L g203 ( .A(n_25), .Y(n_203) );
INVx1_ASAP7_75t_SL g190 ( .A(n_26), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_27), .B(n_133), .Y(n_248) );
AOI33xp33_ASAP7_75t_L g228 ( .A1(n_29), .A2(n_54), .A3(n_126), .B1(n_151), .B2(n_229), .B3(n_230), .Y(n_228) );
NAND2x1_ASAP7_75t_L g550 ( .A(n_30), .B(n_208), .Y(n_550) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_31), .B(n_205), .Y(n_582) );
INVx1_ASAP7_75t_L g131 ( .A(n_32), .Y(n_131) );
OA21x2_ASAP7_75t_L g121 ( .A1(n_33), .A2(n_87), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g172 ( .A(n_33), .B(n_87), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_34), .B(n_155), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_35), .B(n_205), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_36), .B(n_208), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_37), .B(n_205), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_38), .A2(n_499), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g139 ( .A(n_39), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g150 ( .A(n_39), .Y(n_150) );
AND2x2_ASAP7_75t_L g159 ( .A(n_39), .B(n_129), .Y(n_159) );
OR2x6_ASAP7_75t_L g482 ( .A(n_40), .B(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_41), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_42), .B(n_497), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_43), .B(n_155), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g241 ( .A1(n_44), .A2(n_120), .B1(n_197), .B2(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_45), .B(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_46), .B(n_133), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_47), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_48), .B(n_205), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_49), .B(n_175), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_50), .B(n_133), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_51), .A2(n_499), .B(n_581), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_52), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_53), .B(n_205), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_55), .B(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g127 ( .A(n_56), .Y(n_127) );
INVx1_ASAP7_75t_L g135 ( .A(n_56), .Y(n_135) );
AND2x2_ASAP7_75t_L g169 ( .A(n_57), .B(n_170), .Y(n_169) );
AOI221xp5_ASAP7_75t_L g176 ( .A1(n_58), .A2(n_75), .B1(n_148), .B2(n_155), .C(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_59), .B(n_155), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_60), .B(n_208), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_61), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_62), .B(n_120), .Y(n_153) );
AOI21xp5_ASAP7_75t_SL g215 ( .A1(n_63), .A2(n_148), .B(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_64), .A2(n_499), .B(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g200 ( .A(n_65), .Y(n_200) );
AO21x1_ASAP7_75t_L g531 ( .A1(n_66), .A2(n_499), .B(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_67), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g166 ( .A(n_68), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_69), .B(n_497), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_70), .A2(n_148), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g544 ( .A(n_71), .B(n_171), .Y(n_544) );
INVx1_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
INVx1_ASAP7_75t_L g137 ( .A(n_72), .Y(n_137) );
AND2x2_ASAP7_75t_L g585 ( .A(n_73), .B(n_119), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_74), .B(n_155), .Y(n_231) );
AND2x2_ASAP7_75t_L g192 ( .A(n_76), .B(n_119), .Y(n_192) );
INVx1_ASAP7_75t_L g201 ( .A(n_77), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_78), .A2(n_148), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_79), .A2(n_148), .B(n_223), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g807 ( .A(n_80), .Y(n_807) );
INVx1_ASAP7_75t_L g485 ( .A(n_81), .Y(n_485) );
AND2x2_ASAP7_75t_L g494 ( .A(n_82), .B(n_119), .Y(n_494) );
AND2x2_ASAP7_75t_SL g213 ( .A(n_83), .B(n_119), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_84), .B(n_497), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_85), .A2(n_148), .B1(n_226), .B2(n_227), .Y(n_225) );
AND2x2_ASAP7_75t_L g530 ( .A(n_86), .B(n_197), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_88), .B(n_205), .Y(n_509) );
AND2x2_ASAP7_75t_L g553 ( .A(n_89), .B(n_119), .Y(n_553) );
INVx1_ASAP7_75t_L g217 ( .A(n_90), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_91), .B(n_208), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_92), .A2(n_499), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_93), .B(n_205), .Y(n_521) );
AND2x2_ASAP7_75t_L g232 ( .A(n_94), .B(n_119), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_95), .B(n_208), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_96), .A2(n_124), .B(n_130), .C(n_138), .Y(n_123) );
BUFx2_ASAP7_75t_L g799 ( .A(n_97), .Y(n_799) );
BUFx2_ASAP7_75t_SL g819 ( .A(n_97), .Y(n_819) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_98), .A2(n_499), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_99), .B(n_133), .Y(n_218) );
INVxp67_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_477), .B1(n_486), .B2(n_781), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g785 ( .A1(n_110), .A2(n_786), .B1(n_787), .B2(n_788), .Y(n_785) );
NAND3x1_ASAP7_75t_L g110 ( .A(n_111), .B(n_356), .C(n_423), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_316), .Y(n_111) );
NOR3x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_267), .C(n_296), .Y(n_112) );
OAI221xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_181), .B1(n_220), .B2(n_235), .C(n_252), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_SL g430 ( .A1(n_114), .A2(n_194), .B(n_431), .C(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_115), .A2(n_402), .B1(n_405), .B2(n_407), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_115), .B(n_221), .Y(n_476) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_160), .Y(n_115) );
BUFx2_ASAP7_75t_L g395 ( .A(n_116), .Y(n_395) );
INVx1_ASAP7_75t_SL g408 ( .A(n_116), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_116), .B(n_263), .Y(n_450) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g233 ( .A(n_117), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g278 ( .A(n_117), .B(n_174), .Y(n_278) );
INVx1_ASAP7_75t_L g289 ( .A(n_117), .Y(n_289) );
INVx2_ASAP7_75t_L g293 ( .A(n_117), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_117), .B(n_264), .Y(n_420) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_143), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B1(n_141), .B2(n_142), .Y(n_118) );
INVx3_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
INVx4_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_120), .B(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_121), .Y(n_175) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_122), .B(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g197 ( .A(n_122), .B(n_172), .Y(n_197) );
INVxp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_125), .A2(n_166), .B(n_167), .C(n_168), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_125), .A2(n_168), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g189 ( .A1(n_125), .A2(n_168), .B(n_190), .C(n_191), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_125), .A2(n_132), .B1(n_200), .B2(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_125), .A2(n_168), .B(n_217), .C(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g250 ( .A(n_125), .Y(n_250) );
OR2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_128), .Y(n_125) );
AND2x2_ASAP7_75t_L g156 ( .A(n_126), .B(n_157), .Y(n_156) );
INVxp33_ASAP7_75t_L g229 ( .A(n_126), .Y(n_229) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g152 ( .A(n_127), .B(n_140), .Y(n_152) );
AND2x4_ASAP7_75t_L g208 ( .A(n_127), .B(n_136), .Y(n_208) );
INVx3_ASAP7_75t_L g151 ( .A(n_128), .Y(n_151) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x6_ASAP7_75t_L g205 ( .A(n_129), .B(n_134), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g497 ( .A(n_133), .B(n_139), .Y(n_497) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_140), .Y(n_157) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_142), .A2(n_162), .B(n_169), .Y(n_161) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_142), .A2(n_162), .B(n_169), .Y(n_264) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_142), .A2(n_538), .B(n_544), .Y(n_537) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_142), .A2(n_547), .B(n_553), .Y(n_546) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_142), .A2(n_547), .B(n_553), .Y(n_559) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_142), .A2(n_538), .B(n_544), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_147), .B1(n_153), .B2(n_154), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVxp67_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_152), .Y(n_148) );
NOR2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx1_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
AND2x6_ASAP7_75t_L g499 ( .A(n_152), .B(n_159), .Y(n_499) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
INVx1_ASAP7_75t_L g243 ( .A(n_156), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_158), .Y(n_244) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g369 ( .A(n_160), .B(n_370), .Y(n_369) );
NOR2x1_ASAP7_75t_L g160 ( .A(n_161), .B(n_173), .Y(n_160) );
INVx2_ASAP7_75t_L g272 ( .A(n_161), .Y(n_272) );
AND2x2_ASAP7_75t_L g292 ( .A(n_161), .B(n_293), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g417 ( .A(n_161), .B(n_293), .Y(n_417) );
AND2x2_ASAP7_75t_L g442 ( .A(n_161), .B(n_285), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_168), .B(n_197), .Y(n_209) );
INVx1_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_168), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_168), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_168), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_168), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_168), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_168), .A2(n_541), .B(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_168), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_168), .A2(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_168), .A2(n_582), .B(n_583), .Y(n_581) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_170), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_170), .A2(n_496), .B(n_498), .Y(n_495) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_170), .A2(n_519), .B(n_523), .Y(n_518) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_170), .A2(n_519), .B(n_523), .Y(n_589) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g234 ( .A(n_174), .Y(n_234) );
INVx1_ASAP7_75t_L g256 ( .A(n_174), .Y(n_256) );
INVxp67_ASAP7_75t_L g295 ( .A(n_174), .Y(n_295) );
AND2x4_ASAP7_75t_L g335 ( .A(n_174), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_174), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_174), .B(n_286), .Y(n_421) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_180), .Y(n_174) );
INVx2_ASAP7_75t_SL g223 ( .A(n_175), .Y(n_223) );
INVx1_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_193), .Y(n_182) );
AND2x2_ASAP7_75t_L g309 ( .A(n_183), .B(n_281), .Y(n_309) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_184), .Y(n_237) );
AND2x2_ASAP7_75t_L g265 ( .A(n_184), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g276 ( .A(n_184), .Y(n_276) );
INVx1_ASAP7_75t_L g300 ( .A(n_184), .Y(n_300) );
AND2x2_ASAP7_75t_L g303 ( .A(n_184), .B(n_195), .Y(n_303) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_184), .Y(n_325) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_192), .Y(n_184) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_185), .A2(n_579), .B(n_585), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
NOR2x1_ASAP7_75t_L g193 ( .A(n_194), .B(n_210), .Y(n_193) );
AND2x2_ASAP7_75t_L g290 ( .A(n_194), .B(n_212), .Y(n_290) );
NAND2x1_ASAP7_75t_L g323 ( .A(n_194), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g426 ( .A(n_194), .Y(n_426) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx3_ASAP7_75t_L g266 ( .A(n_195), .Y(n_266) );
AND2x2_ASAP7_75t_L g281 ( .A(n_195), .B(n_240), .Y(n_281) );
NOR2x1_ASAP7_75t_SL g350 ( .A(n_195), .B(n_212), .Y(n_350) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_198), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_197), .A2(n_215), .B(n_219), .Y(n_214) );
INVx1_ASAP7_75t_SL g504 ( .A(n_197), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_197), .B(n_536), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_197), .A2(n_571), .B(n_572), .Y(n_570) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_202), .B(n_209), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B1(n_206), .B2(n_207), .Y(n_202) );
INVxp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVxp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_210), .B(n_374), .Y(n_387) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g312 ( .A(n_211), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx4_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
AND2x4_ASAP7_75t_L g258 ( .A(n_212), .B(n_259), .Y(n_258) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_212), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_212), .B(n_275), .Y(n_375) );
AND2x2_ASAP7_75t_L g403 ( .A(n_212), .B(n_240), .Y(n_403) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
NAND2x1_ASAP7_75t_SL g220 ( .A(n_221), .B(n_233), .Y(n_220) );
OR2x2_ASAP7_75t_L g431 ( .A(n_221), .B(n_343), .Y(n_431) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x4_ASAP7_75t_L g271 ( .A(n_222), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g336 ( .A(n_222), .Y(n_336) );
AND2x2_ASAP7_75t_L g370 ( .A(n_222), .B(n_293), .Y(n_370) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_232), .Y(n_222) );
AO21x2_ASAP7_75t_L g286 ( .A1(n_223), .A2(n_224), .B(n_232), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_231), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g343 ( .A(n_233), .Y(n_343) );
AND2x2_ASAP7_75t_L g351 ( .A(n_233), .B(n_284), .Y(n_351) );
AND2x2_ASAP7_75t_L g468 ( .A(n_233), .B(n_271), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g422 ( .A(n_237), .B(n_363), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_237), .B(n_262), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_238), .A2(n_299), .B(n_302), .Y(n_298) );
AND2x2_ASAP7_75t_L g368 ( .A(n_238), .B(n_274), .Y(n_368) );
INVx2_ASAP7_75t_SL g455 ( .A(n_238), .Y(n_455) );
AND2x4_ASAP7_75t_SL g238 ( .A(n_239), .B(n_251), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
INVx2_ASAP7_75t_L g306 ( .A(n_240), .Y(n_306) );
AND2x4_ASAP7_75t_L g313 ( .A(n_240), .B(n_266), .Y(n_313) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_246), .Y(n_240) );
NOR3xp33_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .C(n_245), .Y(n_242) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_251), .Y(n_269) );
AND2x4_ASAP7_75t_L g345 ( .A(n_251), .B(n_259), .Y(n_345) );
OR2x2_ASAP7_75t_L g471 ( .A(n_251), .B(n_472), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g252 ( .A(n_253), .B(n_257), .C(n_260), .D(n_265), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g318 ( .A(n_254), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g415 ( .A(n_254), .Y(n_415) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_255), .B(n_263), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_255), .B(n_320), .Y(n_449) );
BUFx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_258), .B(n_274), .Y(n_327) );
INVx2_ASAP7_75t_L g429 ( .A(n_258), .Y(n_429) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_258), .B(n_299), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_258), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g331 ( .A(n_262), .B(n_278), .Y(n_331) );
AND2x2_ASAP7_75t_L g399 ( .A(n_262), .B(n_335), .Y(n_399) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g284 ( .A(n_263), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_264), .Y(n_338) );
AND2x2_ASAP7_75t_L g389 ( .A(n_264), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_264), .B(n_286), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_265), .B(n_429), .Y(n_436) );
INVx1_ASAP7_75t_SL g472 ( .A(n_265), .Y(n_472) );
INVx1_ASAP7_75t_L g301 ( .A(n_266), .Y(n_301) );
AND2x2_ASAP7_75t_L g363 ( .A(n_266), .B(n_306), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_277), .B(n_279), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
AND2x2_ASAP7_75t_L g329 ( .A(n_271), .B(n_278), .Y(n_329) );
AND2x2_ASAP7_75t_L g437 ( .A(n_271), .B(n_288), .Y(n_437) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g311 ( .A(n_274), .Y(n_311) );
AND2x2_ASAP7_75t_L g344 ( .A(n_274), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g349 ( .A(n_274), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_274), .B(n_313), .Y(n_398) );
NOR3xp33_ASAP7_75t_L g448 ( .A(n_274), .B(n_449), .C(n_450), .Y(n_448) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_283), .B1(n_290), .B2(n_291), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx2_ASAP7_75t_L g374 ( .A(n_281), .Y(n_374) );
AND2x2_ASAP7_75t_L g308 ( .A(n_282), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g330 ( .A(n_282), .B(n_303), .Y(n_330) );
AND2x2_ASAP7_75t_SL g362 ( .A(n_282), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
INVx1_ASAP7_75t_L g341 ( .A(n_284), .Y(n_341) );
AND2x2_ASAP7_75t_L g294 ( .A(n_285), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g383 ( .A(n_289), .B(n_335), .Y(n_383) );
INVx1_ASAP7_75t_L g441 ( .A(n_289), .Y(n_441) );
INVx1_ASAP7_75t_L g297 ( .A(n_291), .Y(n_297) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_292), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g428 ( .A(n_292), .B(n_335), .Y(n_428) );
AND2x2_ASAP7_75t_L g394 ( .A(n_294), .B(n_395), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_294), .B(n_463), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_307), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_299), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g355 ( .A(n_299), .B(n_304), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_299), .B(n_345), .Y(n_406) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_300), .B(n_363), .Y(n_393) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_300), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_302), .A2(n_329), .B1(n_330), .B2(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_SL g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_303), .B(n_345), .Y(n_364) );
INVx1_ASAP7_75t_L g465 ( .A(n_303), .Y(n_465) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_310), .B(n_314), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_309), .B(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g446 ( .A(n_312), .Y(n_446) );
INVx4_ASAP7_75t_L g348 ( .A(n_313), .Y(n_348) );
INVxp33_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g376 ( .A(n_315), .B(n_377), .Y(n_376) );
NOR2x1_ASAP7_75t_L g316 ( .A(n_317), .B(n_332), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_328), .Y(n_317) );
INVx1_ASAP7_75t_L g366 ( .A(n_319), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g371 ( .A(n_323), .Y(n_371) );
INVx1_ASAP7_75t_L g404 ( .A(n_324), .Y(n_404) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g367 ( .A1(n_329), .A2(n_368), .B1(n_369), .B2(n_371), .Y(n_367) );
INVx1_ASAP7_75t_L g381 ( .A(n_330), .Y(n_381) );
NAND4xp25_ASAP7_75t_SL g332 ( .A(n_333), .B(n_339), .C(n_346), .D(n_352), .Y(n_332) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g354 ( .A(n_335), .Y(n_354) );
AND2x2_ASAP7_75t_L g466 ( .A(n_335), .B(n_463), .Y(n_466) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_344), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g473 ( .A(n_343), .B(n_410), .Y(n_473) );
INVx1_ASAP7_75t_L g470 ( .A(n_344), .Y(n_470) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_345), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B(n_351), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_384), .Y(n_356) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_372), .C(n_380), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_365), .B(n_367), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_364), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_394), .B1(n_397), .B2(n_399), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_365), .A2(n_373), .B1(n_376), .B2(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g377 ( .A(n_370), .Y(n_377) );
AND2x4_ASAP7_75t_L g388 ( .A(n_370), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_375), .Y(n_475) );
AOI31xp33_ASAP7_75t_L g474 ( .A1(n_378), .A2(n_451), .A3(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_400), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_396), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_391), .B2(n_394), .Y(n_386) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_390), .Y(n_454) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_411), .Y(n_400) );
AND2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AND2x2_ASAP7_75t_L g412 ( .A(n_403), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_403), .A2(n_461), .B1(n_464), .B2(n_466), .Y(n_460) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_408), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_414), .B1(n_418), .B2(n_422), .Y(n_411) );
NOR2xp33_ASAP7_75t_SL g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx2_ASAP7_75t_SL g463 ( .A(n_420), .Y(n_463) );
INVx2_ASAP7_75t_L g444 ( .A(n_421), .Y(n_444) );
AND2x2_ASAP7_75t_L g423 ( .A(n_424), .B(n_458), .Y(n_423) );
AOI211xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_430), .B(n_433), .C(n_447), .Y(n_424) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B(n_429), .Y(n_425) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_429), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_434), .B(n_438), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_443), .B2(n_445), .Y(n_438) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
AND2x2_ASAP7_75t_L g443 ( .A(n_441), .B(n_444), .Y(n_443) );
AO22x1_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B1(n_452), .B2(n_456), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .C(n_474), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_460), .B(n_467), .Y(n_459) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI21xp33_ASAP7_75t_R g469 ( .A1(n_470), .A2(n_471), .B(n_473), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_478), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
OR2x6_ASAP7_75t_SL g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AND2x6_ASAP7_75t_SL g784 ( .A(n_480), .B(n_482), .Y(n_784) );
OR2x2_ASAP7_75t_L g790 ( .A(n_480), .B(n_482), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_480), .B(n_481), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g787 ( .A(n_487), .Y(n_787) );
NOR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_668), .Y(n_487) );
AO211x2_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_513), .B(n_563), .C(n_636), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND3x2_ASAP7_75t_L g717 ( .A(n_491), .B(n_598), .C(n_614), .Y(n_717) );
AND2x4_ASAP7_75t_L g720 ( .A(n_491), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g576 ( .A(n_492), .B(n_577), .Y(n_576) );
INVx4_ASAP7_75t_L g629 ( .A(n_492), .Y(n_629) );
AND2x2_ASAP7_75t_SL g714 ( .A(n_492), .B(n_623), .Y(n_714) );
AND2x2_ASAP7_75t_L g757 ( .A(n_492), .B(n_578), .Y(n_757) );
INVx5_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
AND2x2_ASAP7_75t_L g625 ( .A(n_493), .B(n_569), .Y(n_625) );
AND2x2_ASAP7_75t_L g643 ( .A(n_493), .B(n_578), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_493), .B(n_577), .Y(n_703) );
NOR2x1_ASAP7_75t_SL g730 ( .A(n_493), .B(n_503), .Y(n_730) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_503), .B(n_569), .Y(n_568) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B(n_511), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_504), .B(n_512), .Y(n_511) );
AO21x2_ASAP7_75t_L g602 ( .A1(n_504), .A2(n_505), .B(n_511), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .Y(n_505) );
AO21x1_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_545), .B(n_554), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OAI22xp33_ASAP7_75t_L g611 ( .A1(n_515), .A2(n_612), .B1(n_616), .B2(n_617), .Y(n_611) );
OR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
AND2x2_ASAP7_75t_L g672 ( .A(n_516), .B(n_560), .Y(n_672) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g605 ( .A(n_517), .B(n_588), .Y(n_605) );
AND2x2_ASAP7_75t_L g677 ( .A(n_517), .B(n_562), .Y(n_677) );
AND2x2_ASAP7_75t_L g696 ( .A(n_517), .B(n_662), .Y(n_696) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g555 ( .A(n_518), .Y(n_555) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_518), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_524), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g656 ( .A(n_525), .B(n_557), .Y(n_656) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
AND2x2_ASAP7_75t_L g560 ( .A(n_526), .B(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g593 ( .A(n_526), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_SL g653 ( .A(n_526), .B(n_589), .Y(n_653) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx2_ASAP7_75t_L g746 ( .A(n_527), .Y(n_746) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g588 ( .A(n_528), .Y(n_588) );
OAI21x1_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_531), .B(n_535), .Y(n_528) );
INVx1_ASAP7_75t_L g536 ( .A(n_530), .Y(n_536) );
INVx2_ASAP7_75t_L g594 ( .A(n_537), .Y(n_594) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_537), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_539), .B(n_543), .Y(n_538) );
INVx2_ASAP7_75t_L g590 ( .A(n_545), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_545), .B(n_722), .Y(n_748) );
AND2x2_ASAP7_75t_L g767 ( .A(n_545), .B(n_757), .Y(n_767) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_SL g635 ( .A(n_546), .B(n_594), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x2_ASAP7_75t_L g634 ( .A(n_555), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_555), .B(n_604), .Y(n_639) );
INVx1_ASAP7_75t_SL g766 ( .A(n_555), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_556), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
INVx1_ASAP7_75t_L g592 ( .A(n_557), .Y(n_592) );
AND2x2_ASAP7_75t_L g778 ( .A(n_557), .B(n_779), .Y(n_778) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g654 ( .A(n_558), .B(n_561), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_558), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g708 ( .A(n_558), .B(n_562), .Y(n_708) );
AND2x2_ASAP7_75t_L g739 ( .A(n_558), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g604 ( .A(n_559), .B(n_562), .Y(n_604) );
INVxp67_ASAP7_75t_L g621 ( .A(n_559), .Y(n_621) );
BUFx3_ASAP7_75t_L g662 ( .A(n_559), .Y(n_662) );
AND2x2_ASAP7_75t_L g682 ( .A(n_560), .B(n_683), .Y(n_682) );
NAND2xp33_ASAP7_75t_L g695 ( .A(n_560), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_561), .B(n_588), .Y(n_651) );
AND2x2_ASAP7_75t_L g740 ( .A(n_561), .B(n_589), .Y(n_740) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g667 ( .A(n_562), .B(n_589), .Y(n_667) );
OR3x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_611), .C(n_626), .Y(n_563) );
OAI321xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_576), .A3(n_586), .B1(n_591), .B2(n_595), .C(n_603), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_568), .Y(n_642) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_568), .Y(n_660) );
OR2x2_ASAP7_75t_L g664 ( .A(n_568), .B(n_576), .Y(n_664) );
BUFx3_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
AND2x2_ASAP7_75t_L g615 ( .A(n_569), .B(n_601), .Y(n_615) );
INVx1_ASAP7_75t_L g632 ( .A(n_569), .Y(n_632) );
INVx2_ASAP7_75t_L g648 ( .A(n_569), .Y(n_648) );
OR2x2_ASAP7_75t_L g687 ( .A(n_569), .B(n_577), .Y(n_687) );
INVx2_ASAP7_75t_L g675 ( .A(n_576), .Y(n_675) );
AND2x2_ASAP7_75t_L g599 ( .A(n_577), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g614 ( .A(n_577), .Y(n_614) );
AND2x4_ASAP7_75t_L g623 ( .A(n_577), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_577), .B(n_600), .Y(n_646) );
AND2x2_ASAP7_75t_L g753 ( .A(n_577), .B(n_648), .Y(n_753) );
INVx4_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_578), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_584), .Y(n_579) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_587), .B(n_590), .Y(n_586) );
AND2x2_ASAP7_75t_L g727 ( .A(n_587), .B(n_654), .Y(n_727) );
INVx1_ASAP7_75t_SL g744 ( .A(n_587), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_587), .B(n_720), .Y(n_773) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
OR2x2_ASAP7_75t_L g616 ( .A(n_588), .B(n_589), .Y(n_616) );
AND2x2_ASAP7_75t_L g709 ( .A(n_590), .B(n_605), .Y(n_709) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_594), .B(n_605), .Y(n_732) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_596), .A2(n_745), .B1(n_750), .B2(n_752), .Y(n_749) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g674 ( .A(n_597), .B(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g769 ( .A(n_597), .B(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g725 ( .A(n_598), .B(n_643), .Y(n_725) );
AND2x4_ASAP7_75t_L g679 ( .A(n_599), .B(n_625), .Y(n_679) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_601), .Y(n_777) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g610 ( .A(n_602), .Y(n_610) );
INVx1_ASAP7_75t_L g624 ( .A(n_602), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .C(n_606), .D(n_607), .Y(n_603) );
AND2x2_ASAP7_75t_L g761 ( .A(n_604), .B(n_746), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_604), .B(n_772), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_605), .B(n_681), .Y(n_680) );
OAI322xp33_ASAP7_75t_L g688 ( .A1(n_605), .A2(n_689), .A3(n_693), .B1(n_695), .B2(n_697), .C1(n_699), .C2(n_704), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_605), .B(n_654), .Y(n_704) );
INVx1_ASAP7_75t_L g772 ( .A(n_605), .Y(n_772) );
INVx2_ASAP7_75t_L g618 ( .A(n_606), .Y(n_618) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_609), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_610), .B(n_629), .Y(n_686) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_613), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g659 ( .A(n_614), .Y(n_659) );
AND2x2_ASAP7_75t_L g731 ( .A(n_614), .B(n_642), .Y(n_731) );
AOI31xp33_ASAP7_75t_L g617 ( .A1(n_615), .A2(n_618), .A3(n_619), .B(n_622), .Y(n_617) );
AND2x2_ASAP7_75t_L g628 ( .A(n_615), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g756 ( .A(n_615), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_SL g763 ( .A(n_615), .B(n_643), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_615), .Y(n_764) );
INVx1_ASAP7_75t_SL g722 ( .A(n_616), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g750 ( .A(n_616), .B(n_744), .C(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g650 ( .A(n_621), .B(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g631 ( .A(n_623), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g692 ( .A(n_623), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g774 ( .A1(n_623), .A2(n_653), .A3(n_656), .B1(n_775), .B2(n_776), .C1(n_778), .C2(n_780), .Y(n_774) );
AND2x2_ASAP7_75t_L g780 ( .A(n_623), .B(n_629), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_630), .B(n_633), .Y(n_626) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_629), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g775 ( .A(n_629), .B(n_662), .Y(n_775) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g701 ( .A(n_632), .Y(n_701) );
AND2x2_ASAP7_75t_L g729 ( .A(n_632), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g776 ( .A(n_632), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g681 ( .A(n_635), .Y(n_681) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
O2A1O1Ixp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_641), .C(n_644), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND2x2_ASAP7_75t_L g698 ( .A(n_643), .B(n_648), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B(n_655), .C(n_657), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_645), .A2(n_671), .B1(n_673), .B2(n_676), .C(n_678), .Y(n_670) );
OR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g690 ( .A(n_647), .Y(n_690) );
OR2x2_ASAP7_75t_L g710 ( .A(n_647), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g755 ( .A(n_650), .Y(n_755) );
INVx1_ASAP7_75t_L g779 ( .A(n_651), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_653), .B(n_654), .Y(n_652) );
AND2x2_ASAP7_75t_L g661 ( .A(n_653), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_653), .B(n_723), .Y(n_735) );
INVx1_ASAP7_75t_L g715 ( .A(n_654), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_663), .B2(n_665), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_SL g723 ( .A(n_662), .Y(n_723) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND4xp75_ASAP7_75t_L g668 ( .A(n_669), .B(n_705), .C(n_733), .D(n_758), .Y(n_668) );
NOR2xp67_ASAP7_75t_L g669 ( .A(n_670), .B(n_688), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_SL g745 ( .A(n_677), .B(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_684), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_681), .B(n_744), .Y(n_743) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_L g721 ( .A(n_687), .Y(n_721) );
OR2x2_ASAP7_75t_L g736 ( .A(n_687), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g751 ( .A(n_696), .Y(n_751) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_698), .A2(n_743), .B(n_745), .Y(n_742) );
INVxp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_718), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_710), .B1(n_713), .B2(n_715), .C(n_716), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g754 ( .A1(n_708), .A2(n_755), .B(n_756), .Y(n_754) );
INVx3_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
OAI322xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .A3(n_723), .B1(n_724), .B2(n_726), .C1(n_728), .C2(n_732), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
NOR2x1_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx1_ASAP7_75t_L g741 ( .A(n_729), .Y(n_741) );
INVx1_ASAP7_75t_L g737 ( .A(n_730), .Y(n_737) );
AND2x2_ASAP7_75t_L g752 ( .A(n_730), .B(n_753), .Y(n_752) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_747), .Y(n_733) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_738), .B2(n_741), .C(n_742), .Y(n_734) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
OAI211xp5_ASAP7_75t_SL g747 ( .A1(n_741), .A2(n_748), .B(n_749), .C(n_754), .Y(n_747) );
INVx2_ASAP7_75t_SL g770 ( .A(n_757), .Y(n_770) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_759), .B(n_768), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_762), .B1(n_764), .B2(n_765), .Y(n_759) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
OAI211xp5_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_771), .B(n_773), .C(n_774), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx3_ASAP7_75t_SL g782 ( .A(n_783), .Y(n_782) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_784), .Y(n_788) );
XOR2x2_ASAP7_75t_L g804 ( .A(n_787), .B(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_SL g792 ( .A(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_800), .Y(n_793) );
INVxp67_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_SL g795 ( .A(n_796), .B(n_799), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
OR2x2_ASAP7_75t_SL g814 ( .A(n_797), .B(n_799), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_797), .A2(n_817), .B(n_820), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_800), .B(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
BUFx2_ASAP7_75t_R g810 ( .A(n_801), .Y(n_810) );
BUFx2_ASAP7_75t_L g821 ( .A(n_801), .Y(n_821) );
INVxp33_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_808), .B(n_811), .Y(n_803) );
INVx1_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
CKINVDCx11_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
CKINVDCx8_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
endmodule