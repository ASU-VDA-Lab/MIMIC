module fake_ariane_1139_n_1208 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1208);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1208;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_1174;
wire n_640;
wire n_197;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_176;
wire n_404;
wire n_172;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_183;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_1169;
wire n_789;
wire n_788;
wire n_908;
wire n_850;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_1029;
wire n_341;
wire n_205;
wire n_985;
wire n_421;
wire n_245;
wire n_1167;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_906;
wire n_690;
wire n_416;
wire n_1180;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_1154;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_1138;
wire n_1149;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_1196;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_1181;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_162;
wire n_1131;
wire n_765;
wire n_1187;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_1177;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_1170;
wire n_1151;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_905;
wire n_279;
wire n_958;
wire n_702;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_207;
wire n_363;
wire n_720;
wire n_1067;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_1163;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_186;
wire n_801;
wire n_1184;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_1173;
wire n_311;
wire n_239;
wire n_402;
wire n_1068;
wire n_1052;
wire n_272;
wire n_829;
wire n_1198;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_167;
wire n_422;
wire n_1106;
wire n_784;
wire n_648;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_158;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_1201;
wire n_1107;
wire n_173;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_331;
wire n_309;
wire n_559;
wire n_1134;
wire n_1185;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_1141;
wire n_350;
wire n_291;
wire n_822;
wire n_1143;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_721;
wire n_600;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_1099;
wire n_1153;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_1145;
wire n_971;
wire n_240;
wire n_369;
wire n_1192;
wire n_224;
wire n_894;
wire n_787;
wire n_1105;
wire n_547;
wire n_1195;
wire n_420;
wire n_562;
wire n_518;
wire n_677;
wire n_604;
wire n_614;
wire n_439;
wire n_1172;
wire n_222;
wire n_478;
wire n_703;
wire n_1207;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_868;
wire n_256;
wire n_831;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_1160;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_1085;
wire n_1152;
wire n_432;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_1197;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_1165;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_192;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_1205;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_163;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_1156;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_1202;
wire n_627;
wire n_1039;
wire n_1188;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_1150;
wire n_233;
wire n_728;
wire n_957;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_685;
wire n_459;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_1142;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_1194;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_1159;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_847;
wire n_939;
wire n_1135;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_178;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_1038;
wire n_201;
wire n_572;
wire n_343;
wire n_1199;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_1193;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_947;
wire n_171;
wire n_409;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_1179;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_1081;
wire n_1166;
wire n_182;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_1158;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_774;
wire n_407;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_1168;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_1157;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_1182;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_179;
wire n_1126;
wire n_395;
wire n_621;
wire n_1178;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_213;
wire n_862;
wire n_895;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_626;
wire n_430;
wire n_493;
wire n_722;
wire n_1206;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1146;
wire n_1100;
wire n_1171;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_1203;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_999;
wire n_1083;
wire n_998;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_174;
wire n_275;
wire n_704;
wire n_1060;
wire n_1175;
wire n_1044;
wire n_1148;
wire n_751;
wire n_1027;
wire n_615;
wire n_1070;
wire n_204;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1139;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_159;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1189;
wire n_1124;
wire n_250;
wire n_932;
wire n_1183;
wire n_773;
wire n_165;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_1110;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_944;
wire n_749;
wire n_1204;
wire n_994;
wire n_289;
wire n_548;
wire n_815;
wire n_542;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_782;
wire n_650;
wire n_856;
wire n_425;
wire n_1161;
wire n_431;
wire n_1176;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1155;
wire n_1191;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_1164;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_191;
wire n_797;
wire n_489;
wire n_480;
wire n_1011;
wire n_642;
wire n_211;
wire n_978;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_1147;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_30),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_37),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_1),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_17),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_153),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_28),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_111),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_71),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_66),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_26),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_54),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_5),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_47),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_59),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_65),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_106),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_56),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_3),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_97),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_137),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_101),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_17),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_126),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_41),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_94),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_77),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_151),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_108),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_99),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_20),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_92),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_157),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_4),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_67),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_93),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_16),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_170),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_187),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_181),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_161),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_159),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_168),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_164),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_202),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_167),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_169),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_238),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_242),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_232),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_234),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_234),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_237),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_243),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_224),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_230),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_227),
.B(n_203),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_228),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_236),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_236),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_216),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_217),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_217),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_217),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_217),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_217),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_217),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_267),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_267),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_289),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_290),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_288),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_274),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_288),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_247),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_248),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_294),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

INVxp67_ASAP7_75t_SL g321 ( 
.A(n_256),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_295),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_296),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_251),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

INVxp33_ASAP7_75t_SL g332 ( 
.A(n_296),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_297),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_297),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_265),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_271),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_268),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_273),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_268),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_250),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_347),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_298),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_347),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_261),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_300),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_300),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_307),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_307),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_299),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_323),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_262),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_310),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_311),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_306),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_311),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_319),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_319),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_326),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_339),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_313),
.B(n_315),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_340),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_333),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_333),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_301),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_R g384 ( 
.A(n_324),
.B(n_277),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_302),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_344),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_317),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_305),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_280),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_349),
.B(n_312),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_362),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_377),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_384),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_353),
.A2(n_334),
.B1(n_252),
.B2(n_250),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_370),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_371),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_375),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_252),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_283),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_383),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_382),
.B(n_330),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_386),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_389),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_320),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_390),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_351),
.Y(n_414)
);

OAI21x1_ASAP7_75t_L g415 ( 
.A1(n_376),
.A2(n_308),
.B(n_328),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_345),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_352),
.B(n_318),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_391),
.Y(n_421)
);

AND2x6_ASAP7_75t_L g422 ( 
.A(n_350),
.B(n_345),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_354),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_368),
.B(n_321),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_360),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_366),
.B(n_335),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_369),
.B(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_373),
.B(n_162),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_378),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_325),
.Y(n_436)
);

BUFx12f_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_388),
.B(n_337),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_367),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_367),
.B(n_276),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_361),
.B(n_279),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_357),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_349),
.B(n_281),
.Y(n_447)
);

CKINVDCx8_ASAP7_75t_R g448 ( 
.A(n_352),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_383),
.B(n_304),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_374),
.B(n_342),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_357),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_364),
.A2(n_282),
.B1(n_212),
.B2(n_278),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_349),
.B(n_284),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_364),
.A2(n_308),
.B1(n_331),
.B2(n_329),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_364),
.B(n_328),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_364),
.B(n_329),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_357),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_357),
.Y(n_463)
);

BUFx8_ASAP7_75t_SL g464 ( 
.A(n_351),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_364),
.B(n_331),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_351),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_413),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_444),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_447),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_413),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_393),
.B(n_285),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_395),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_392),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_464),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_403),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_393),
.B(n_285),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_402),
.B(n_309),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_443),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_405),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_412),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_442),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_450),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_410),
.B(n_322),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_416),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_419),
.B(n_163),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_446),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_449),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_452),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_464),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_457),
.Y(n_501)
);

AND3x1_ASAP7_75t_L g502 ( 
.A(n_400),
.B(n_272),
.C(n_336),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_402),
.B(n_272),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_414),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_462),
.Y(n_507)
);

INVx5_ASAP7_75t_L g508 ( 
.A(n_453),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_419),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_411),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_428),
.B(n_191),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_463),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_437),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_410),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_410),
.B(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_397),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_428),
.B(n_426),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_432),
.B(n_184),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_453),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_510),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_510),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_478),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_474),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_478),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_470),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_500),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_500),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_431),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_513),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_506),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_476),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_506),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_495),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_R g535 ( 
.A(n_470),
.B(n_448),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_495),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_425),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_475),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_492),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_484),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_477),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_508),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_473),
.B(n_426),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_489),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_503),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_471),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_501),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_518),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_479),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_481),
.B(n_418),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_515),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_518),
.Y(n_556)
);

BUFx10_ASAP7_75t_L g557 ( 
.A(n_468),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_538),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_508),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_525),
.B(n_549),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_545),
.A2(n_502),
.B1(n_461),
.B2(n_465),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_557),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_541),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_553),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_523),
.Y(n_565)
);

AO21x2_ASAP7_75t_L g566 ( 
.A1(n_523),
.A2(n_460),
.B(n_415),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_530),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_537),
.B(n_508),
.Y(n_568)
);

BUFx10_ASAP7_75t_L g569 ( 
.A(n_522),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_525),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_544),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_532),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_511),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_539),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_550),
.A2(n_440),
.B1(n_398),
.B2(n_515),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_555),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_535),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_544),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_555),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_542),
.Y(n_584)
);

BUFx10_ASAP7_75t_L g585 ( 
.A(n_522),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_542),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_557),
.Y(n_587)
);

NAND3xp33_ASAP7_75t_L g588 ( 
.A(n_540),
.B(n_456),
.C(n_461),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_552),
.A2(n_465),
.B1(n_407),
.B2(n_480),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_552),
.A2(n_431),
.B1(n_438),
.B2(n_407),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_550),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_557),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_548),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_534),
.Y(n_594)
);

INVx4_ASAP7_75t_L g595 ( 
.A(n_521),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_551),
.B(n_441),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

NAND2xp33_ASAP7_75t_SL g598 ( 
.A(n_543),
.B(n_467),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_543),
.B(n_485),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_524),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_543),
.B(n_467),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_529),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_546),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_546),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_526),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_531),
.B(n_421),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_533),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_527),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_545),
.B(n_490),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_538),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_538),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_538),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_521),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_538),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_538),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_550),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_525),
.B(n_485),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_525),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_538),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_521),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_525),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_544),
.B(n_490),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

INVx8_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_535),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_545),
.B(n_490),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_538),
.Y(n_630)
);

AO21x2_ASAP7_75t_L g631 ( 
.A1(n_523),
.A2(n_458),
.B(n_491),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_538),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_525),
.B(n_491),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_525),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_525),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_538),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_538),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_525),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_538),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_538),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_538),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_560),
.B(n_441),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_564),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_615),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_558),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_622),
.Y(n_647)
);

AO21x2_ASAP7_75t_L g648 ( 
.A1(n_566),
.A2(n_417),
.B(n_516),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_561),
.B(n_494),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_634),
.B(n_519),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_567),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_630),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_616),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_580),
.B(n_438),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_582),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_636),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_574),
.B(n_486),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_621),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_571),
.B(n_519),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_619),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_574),
.B(n_487),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_563),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_613),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_583),
.B(n_438),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_571),
.B(n_497),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_561),
.B(n_440),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_621),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_635),
.B(n_498),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_635),
.B(n_499),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_576),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_576),
.Y(n_672)
);

INVx4_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_627),
.Y(n_674)
);

OAI22x1_ASAP7_75t_L g675 ( 
.A1(n_579),
.A2(n_588),
.B1(n_577),
.B2(n_601),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_589),
.B(n_494),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_637),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_620),
.B(n_505),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_620),
.B(n_507),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_582),
.B(n_519),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_627),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_639),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_621),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_624),
.B(n_638),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_641),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_614),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_617),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_624),
.B(n_494),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_589),
.A2(n_493),
.B1(n_514),
.B2(n_422),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_618),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_588),
.A2(n_590),
.B1(n_575),
.B2(n_493),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_619),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_624),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_638),
.B(n_494),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_626),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_632),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_597),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_616),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_640),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_638),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_565),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_628),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_592),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_625),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_633),
.B(n_512),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_612),
.B(n_469),
.Y(n_706)
);

OAI21xp33_ASAP7_75t_L g707 ( 
.A1(n_590),
.A2(n_406),
.B(n_429),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_578),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_592),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_584),
.B(n_504),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_562),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_625),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_612),
.B(n_472),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_599),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_570),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_573),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_586),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_631),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_599),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_562),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_572),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_631),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_629),
.B(n_483),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_655),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_643),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_684),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_658),
.B(n_629),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_684),
.B(n_572),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_712),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_645),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_667),
.A2(n_581),
.B1(n_591),
.B2(n_594),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_647),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_718),
.Y(n_734)
);

BUFx6f_ASAP7_75t_SL g735 ( 
.A(n_653),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_646),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_698),
.B(n_595),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_708),
.B(n_609),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_671),
.B(n_572),
.Y(n_739)
);

AOI22x1_ASAP7_75t_L g740 ( 
.A1(n_673),
.A2(n_595),
.B1(n_623),
.B2(n_425),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_652),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_671),
.B(n_572),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_657),
.Y(n_743)
);

OR2x2_ASAP7_75t_SL g744 ( 
.A(n_658),
.B(n_607),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_677),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_672),
.B(n_607),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_662),
.B(n_596),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_722),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_704),
.B(n_605),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_662),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_683),
.B(n_604),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_693),
.B(n_642),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_667),
.A2(n_466),
.B1(n_607),
.B2(n_623),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_697),
.B(n_610),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_663),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_702),
.B(n_423),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_722),
.Y(n_758)
);

NOR2x1p5_ASAP7_75t_L g759 ( 
.A(n_672),
.B(n_437),
.Y(n_759)
);

BUFx4f_ASAP7_75t_L g760 ( 
.A(n_722),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_722),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_715),
.B(n_659),
.Y(n_762)
);

NAND2xp33_ASAP7_75t_L g763 ( 
.A(n_707),
.B(n_422),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_702),
.B(n_423),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_685),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_661),
.A2(n_466),
.B1(n_603),
.B2(n_608),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_644),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_687),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_690),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_644),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_653),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_695),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_659),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_664),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_715),
.B(n_587),
.Y(n_776)
);

NAND2x1p5_ASAP7_75t_L g777 ( 
.A(n_673),
.B(n_568),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_691),
.A2(n_596),
.B1(n_397),
.B2(n_399),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_696),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_654),
.B(n_593),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_699),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_668),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_668),
.B(n_606),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_665),
.B(n_611),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_700),
.B(n_569),
.Y(n_785)
);

AO22x2_ASAP7_75t_L g786 ( 
.A1(n_723),
.A2(n_651),
.B1(n_720),
.B2(n_719),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_700),
.B(n_569),
.Y(n_787)
);

INVx2_ASAP7_75t_SL g788 ( 
.A(n_674),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_709),
.B(n_568),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_666),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_709),
.B(n_602),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_651),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_689),
.A2(n_422),
.B1(n_496),
.B2(n_435),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_666),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_678),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_669),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_669),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_674),
.B(n_585),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_670),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_794),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_750),
.B(n_670),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_747),
.B(n_676),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_732),
.B(n_675),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_795),
.B(n_676),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_754),
.B(n_649),
.C(n_712),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_795),
.B(n_678),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_737),
.B(n_772),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_792),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_797),
.B(n_679),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_789),
.B(n_681),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_728),
.B(n_679),
.Y(n_811)
);

OAI221xp5_ASAP7_75t_L g812 ( 
.A1(n_763),
.A2(n_649),
.B1(n_689),
.B2(n_705),
.C(n_691),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_738),
.B(n_692),
.Y(n_813)
);

INVx8_ASAP7_75t_L g814 ( 
.A(n_735),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_790),
.B(n_705),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_735),
.B(n_681),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_755),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_796),
.B(n_799),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_778),
.A2(n_713),
.B1(n_704),
.B2(n_459),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_725),
.B(n_710),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_726),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_776),
.Y(n_822)
);

OAI221xp5_ASAP7_75t_L g823 ( 
.A1(n_793),
.A2(n_433),
.B1(n_427),
.B2(n_430),
.C(n_459),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_776),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_734),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_784),
.A2(n_422),
.B1(n_713),
.B2(n_704),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_762),
.B(n_710),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_766),
.B(n_585),
.Y(n_828)
);

AOI221xp5_ASAP7_75t_L g829 ( 
.A1(n_731),
.A2(n_200),
.B1(n_199),
.B2(n_203),
.C(n_436),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_798),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_762),
.B(n_724),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_730),
.A2(n_721),
.B(n_703),
.C(n_660),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_757),
.B(n_600),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_753),
.B(n_733),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_706),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_789),
.B(n_704),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_736),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_785),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_788),
.B(n_713),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_740),
.B(n_423),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_756),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_729),
.B(n_713),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_743),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_745),
.B(n_706),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_752),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_764),
.B(n_600),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_780),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_765),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_739),
.A2(n_742),
.B1(n_777),
.B2(n_714),
.Y(n_849)
);

AND2x6_ASAP7_75t_SL g850 ( 
.A(n_787),
.B(n_411),
.Y(n_850)
);

NAND2x1_ASAP7_75t_L g851 ( 
.A(n_730),
.B(n_721),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_746),
.B(n_423),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_767),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_L g854 ( 
.A(n_740),
.B(n_434),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_727),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_774),
.Y(n_856)
);

NOR2x1_ASAP7_75t_L g857 ( 
.A(n_759),
.B(n_703),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_782),
.B(n_714),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_769),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_751),
.B(n_660),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_770),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_773),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_749),
.A2(n_422),
.B1(n_496),
.B2(n_493),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_779),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_751),
.B(n_688),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_775),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_781),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_783),
.Y(n_868)
);

OR2x6_ASAP7_75t_L g869 ( 
.A(n_729),
.B(n_650),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_786),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_786),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_791),
.B(n_688),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_791),
.B(n_694),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_749),
.A2(n_404),
.B1(n_717),
.B2(n_399),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_768),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_744),
.A2(n_650),
.B1(n_656),
.B2(n_644),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_748),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_783),
.B(n_694),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_748),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_822),
.B(n_771),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_870),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_821),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_824),
.B(n_771),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_803),
.A2(n_433),
.B(n_760),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_871),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_802),
.B(n_768),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_855),
.B(n_768),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_808),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_869),
.B(n_749),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_832),
.B(n_748),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_825),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_807),
.B(n_434),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_817),
.B(n_758),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_800),
.B(n_758),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_843),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_811),
.B(n_758),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_814),
.B(n_434),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_804),
.B(n_801),
.Y(n_898)
);

BUFx4f_ASAP7_75t_L g899 ( 
.A(n_814),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_835),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_838),
.B(n_761),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_851),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_806),
.B(n_761),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_868),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_844),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_853),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_827),
.B(n_856),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_820),
.B(n_761),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_859),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_845),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_848),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_861),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_809),
.B(n_749),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_R g914 ( 
.A(n_814),
.B(n_424),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_879),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_862),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_865),
.B(n_760),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_869),
.B(n_644),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_816),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_869),
.B(n_656),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_858),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_805),
.A2(n_424),
.B(n_496),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_830),
.B(n_656),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_L g924 ( 
.A1(n_831),
.A2(n_404),
.B(n_421),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_828),
.B(n_434),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_834),
.Y(n_926)
);

OR2x2_ASAP7_75t_SL g927 ( 
.A(n_860),
.B(n_439),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_847),
.B(n_648),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_815),
.B(n_711),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_842),
.B(n_711),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_864),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_876),
.B(n_701),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_818),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_813),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_833),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_876),
.B(n_439),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_902),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_933),
.B(n_900),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_884),
.A2(n_935),
.B1(n_926),
.B2(n_927),
.Y(n_939)
);

AND2x2_ASAP7_75t_SL g940 ( 
.A(n_899),
.B(n_840),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_935),
.B(n_849),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_905),
.B(n_872),
.Y(n_942)
);

A2O1A1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_922),
.A2(n_823),
.B(n_812),
.C(n_829),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_936),
.A2(n_854),
.B(n_810),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_L g945 ( 
.A1(n_913),
.A2(n_826),
.B1(n_863),
.B2(n_873),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_924),
.A2(n_863),
.B(n_852),
.C(n_826),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_927),
.A2(n_857),
.B1(n_874),
.B2(n_846),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_936),
.A2(n_836),
.B(n_839),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_921),
.B(n_850),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_882),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_898),
.B(n_850),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_889),
.B(n_879),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_914),
.B(n_879),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_890),
.A2(n_878),
.B(n_877),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_890),
.A2(n_877),
.B(n_875),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_902),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_906),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_882),
.B(n_866),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_895),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_899),
.A2(n_875),
.B(n_598),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_895),
.B(n_867),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_906),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_928),
.A2(n_819),
.B(n_837),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_909),
.B(n_841),
.Y(n_964)
);

NOR3xp33_ASAP7_75t_L g965 ( 
.A(n_925),
.B(n_602),
.C(n_451),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_919),
.B(n_439),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_919),
.B(n_439),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_889),
.B(n_648),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_899),
.A2(n_598),
.B(n_559),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_889),
.B(n_716),
.Y(n_970)
);

BUFx4f_ASAP7_75t_L g971 ( 
.A(n_918),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_904),
.A2(n_177),
.B(n_179),
.C(n_163),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_912),
.B(n_680),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_915),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_SL g975 ( 
.A1(n_932),
.A2(n_482),
.B(n_468),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_912),
.B(n_680),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_916),
.B(n_680),
.Y(n_977)
);

OR2x2_ASAP7_75t_SL g978 ( 
.A(n_934),
.B(n_468),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_932),
.A2(n_214),
.B(n_177),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_928),
.A2(n_194),
.B(n_454),
.C(n_420),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_916),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_932),
.A2(n_454),
.B(n_504),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_902),
.B(n_504),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_918),
.B(n_504),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_931),
.B(n_680),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_897),
.A2(n_173),
.B(n_175),
.C(n_172),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_929),
.A2(n_930),
.B1(n_881),
.B2(n_885),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_892),
.B(n_0),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_880),
.B(n_0),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_910),
.B(n_680),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_918),
.B(n_504),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_920),
.A2(n_896),
.B1(n_915),
.B2(n_886),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_915),
.A2(n_509),
.B(n_482),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_911),
.Y(n_994)
);

INVxp67_ASAP7_75t_L g995 ( 
.A(n_887),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_920),
.B(n_509),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_930),
.A2(n_176),
.B(n_178),
.C(n_180),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_891),
.Y(n_998)
);

AO22x1_ASAP7_75t_L g999 ( 
.A1(n_949),
.A2(n_893),
.B1(n_885),
.B2(n_881),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_995),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_941),
.A2(n_894),
.B(n_903),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_938),
.B(n_907),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_943),
.A2(n_940),
.B(n_953),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_994),
.B(n_907),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_951),
.B(n_880),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_939),
.A2(n_893),
.B(n_883),
.Y(n_1006)
);

NOR3xp33_ASAP7_75t_L g1007 ( 
.A(n_966),
.B(n_883),
.C(n_887),
.Y(n_1007)
);

CKINVDCx10_ASAP7_75t_R g1008 ( 
.A(n_967),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_974),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_SL g1010 ( 
.A(n_989),
.B(n_920),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_963),
.A2(n_930),
.B1(n_891),
.B2(n_888),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_971),
.B(n_917),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_955),
.A2(n_908),
.B(n_901),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_944),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_957),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_967),
.B(n_917),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_954),
.A2(n_923),
.B(n_901),
.C(n_908),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_971),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_1008),
.B(n_988),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1014),
.B(n_950),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_1003),
.B(n_972),
.C(n_997),
.Y(n_1021)
);

HAxp5_ASAP7_75t_L g1022 ( 
.A(n_1000),
.B(n_1013),
.CON(n_1022),
.SN(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_1018),
.A2(n_980),
.B(n_979),
.C(n_965),
.Y(n_1023)
);

BUFx12f_ASAP7_75t_L g1024 ( 
.A(n_1009),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_1018),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1002),
.B(n_959),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_1010),
.B(n_937),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1012),
.A2(n_975),
.B(n_947),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_1005),
.A2(n_956),
.B(n_937),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_999),
.A2(n_952),
.B(n_992),
.Y(n_1030)
);

AOI21x1_ASAP7_75t_L g1031 ( 
.A1(n_1006),
.A2(n_962),
.B(n_981),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1009),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_SL g1033 ( 
.A1(n_1007),
.A2(n_956),
.B(n_960),
.C(n_948),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_1009),
.B(n_974),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1016),
.B(n_923),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1004),
.B(n_1001),
.Y(n_1036)
);

INVx5_ASAP7_75t_L g1037 ( 
.A(n_1016),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1015),
.B(n_942),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_1017),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1011),
.B(n_958),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_1003),
.A2(n_961),
.B(n_945),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_1003),
.A2(n_983),
.B(n_969),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1004),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_1037),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1020),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1035),
.B(n_974),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1039),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_1025),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_1041),
.B(n_987),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1036),
.B(n_1043),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_1032),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1045),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1047),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1049),
.A2(n_1033),
.B(n_1042),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_1053),
.Y(n_1055)
);

HB1xp67_ASAP7_75t_L g1056 ( 
.A(n_1052),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_1031),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_1055),
.A2(n_1048),
.B(n_1050),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

AO21x2_ASAP7_75t_L g1060 ( 
.A1(n_1058),
.A2(n_1051),
.B(n_1021),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1060),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1060),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_1061),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1062),
.B(n_1044),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1063),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1064),
.B(n_1046),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1066),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1065),
.Y(n_1068)
);

AOI22x1_ASAP7_75t_L g1069 ( 
.A1(n_1066),
.A2(n_1059),
.B1(n_1024),
.B2(n_1051),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_1068),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1067),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_1019),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_1070),
.B(n_1037),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1071),
.B(n_1072),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_1073),
.B(n_1037),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_1073),
.B(n_1074),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_1040),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1076),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1078),
.A2(n_1022),
.B(n_1034),
.C(n_1030),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1077),
.B(n_1038),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1080),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1079),
.B(n_1029),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1081),
.B(n_1029),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_1082),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1084),
.B(n_1028),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1083),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1083),
.Y(n_1087)
);

NAND4xp75_ASAP7_75t_SL g1088 ( 
.A(n_1086),
.B(n_3),
.C(n_1),
.D(n_2),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1087),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1085),
.B(n_2),
.Y(n_1090)
);

O2A1O1Ixp33_ASAP7_75t_SL g1091 ( 
.A1(n_1090),
.A2(n_1027),
.B(n_1026),
.C(n_986),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1089),
.A2(n_1023),
.B(n_409),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1092),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1091),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1094),
.B(n_1088),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1093),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1096),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1095),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_1097),
.B(n_1098),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1097),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1100),
.B(n_182),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_L g1103 ( 
.A(n_1101),
.B(n_1102),
.C(n_185),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1101),
.A2(n_186),
.B(n_183),
.Y(n_1104)
);

OAI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1101),
.A2(n_188),
.B1(n_189),
.B2(n_193),
.C(n_195),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1103),
.A2(n_198),
.B(n_197),
.Y(n_1106)
);

AOI21xp33_ASAP7_75t_L g1107 ( 
.A1(n_1104),
.A2(n_204),
.B(n_201),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1105),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_1106),
.Y(n_1109)
);

INVx1_ASAP7_75t_SL g1110 ( 
.A(n_1107),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1109),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1110),
.B(n_5),
.Y(n_1112)
);

NOR2x1p5_ASAP7_75t_SL g1113 ( 
.A(n_1111),
.B(n_205),
.Y(n_1113)
);

AOI221x1_ASAP7_75t_L g1114 ( 
.A1(n_1112),
.A2(n_207),
.B1(n_208),
.B2(n_210),
.C(n_211),
.Y(n_1114)
);

AOI211x1_ASAP7_75t_L g1115 ( 
.A1(n_1114),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_1115)
);

NOR3xp33_ASAP7_75t_L g1116 ( 
.A(n_1113),
.B(n_213),
.C(n_6),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1116),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1115),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1118),
.B(n_7),
.Y(n_1119)
);

BUFx2_ASAP7_75t_L g1120 ( 
.A(n_1117),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_9),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_L g1123 ( 
.A(n_1120),
.B(n_409),
.C(n_10),
.Y(n_1123)
);

NAND3x1_ASAP7_75t_L g1124 ( 
.A(n_1122),
.B(n_11),
.C(n_12),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1123),
.A2(n_409),
.B(n_13),
.C(n_14),
.Y(n_1125)
);

OAI221xp5_ASAP7_75t_L g1126 ( 
.A1(n_1121),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_1126)
);

NAND3xp33_ASAP7_75t_L g1127 ( 
.A(n_1126),
.B(n_15),
.C(n_16),
.Y(n_1127)
);

OAI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_1125),
.A2(n_1124),
.B(n_18),
.Y(n_1128)
);

NOR3x1_ASAP7_75t_L g1129 ( 
.A(n_1127),
.B(n_18),
.C(n_19),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_1128),
.B(n_998),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1129),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_L g1132 ( 
.A(n_1130),
.B(n_993),
.Y(n_1132)
);

NOR3x2_ASAP7_75t_L g1133 ( 
.A(n_1131),
.B(n_19),
.C(n_20),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1132),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_21),
.B(n_22),
.Y(n_1135)
);

AO22x2_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1136),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1135),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1137),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1138),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1137),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1140),
.B(n_1141),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1139),
.Y(n_1143)
);

OAI22x1_ASAP7_75t_L g1144 ( 
.A1(n_1140),
.A2(n_24),
.B1(n_25),
.B2(n_970),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_1142),
.Y(n_1145)
);

CKINVDCx12_ASAP7_75t_R g1146 ( 
.A(n_1143),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_1146),
.Y(n_1147)
);

AO22x2_ASAP7_75t_L g1148 ( 
.A1(n_1145),
.A2(n_1144),
.B1(n_25),
.B2(n_24),
.Y(n_1148)
);

OA22x2_ASAP7_75t_L g1149 ( 
.A1(n_1147),
.A2(n_968),
.B1(n_29),
.B2(n_31),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1148),
.B(n_27),
.Y(n_1150)
);

OAI221xp5_ASAP7_75t_L g1151 ( 
.A1(n_1150),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.C(n_35),
.Y(n_1151)
);

XOR2xp5_ASAP7_75t_L g1152 ( 
.A(n_1149),
.B(n_36),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1151),
.A2(n_1152),
.B(n_991),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1151),
.B(n_968),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1154),
.A2(n_996),
.B1(n_984),
.B2(n_985),
.C(n_977),
.Y(n_1155)
);

XNOR2xp5_ASAP7_75t_L g1156 ( 
.A(n_1153),
.B(n_38),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1156),
.Y(n_1157)
);

AOI21xp33_ASAP7_75t_SL g1158 ( 
.A1(n_1155),
.A2(n_39),
.B(n_40),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1156),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1159),
.A2(n_978),
.B1(n_976),
.B2(n_973),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1157),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1158),
.A2(n_946),
.B(n_990),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1159),
.B(n_42),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1161),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1163),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1162),
.A2(n_46),
.B(n_48),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1165),
.B(n_1160),
.Y(n_1167)
);

OAI22x1_ASAP7_75t_L g1168 ( 
.A1(n_1164),
.A2(n_1166),
.B1(n_50),
.B2(n_51),
.Y(n_1168)
);

OAI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1165),
.A2(n_49),
.B1(n_53),
.B2(n_55),
.C(n_57),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_SL g1170 ( 
.A(n_1167),
.B(n_58),
.C(n_60),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1169),
.A2(n_61),
.B(n_62),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1168),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1167),
.A2(n_70),
.B(n_72),
.C(n_73),
.Y(n_1173)
);

OAI21xp33_ASAP7_75t_L g1174 ( 
.A1(n_1167),
.A2(n_74),
.B(n_75),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1167),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_1175)
);

OAI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1167),
.A2(n_81),
.B(n_82),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1167),
.Y(n_1177)
);

OAI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1167),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_SL g1179 ( 
.A1(n_1167),
.A2(n_87),
.B(n_88),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1167),
.B(n_89),
.Y(n_1180)
);

OA21x2_ASAP7_75t_L g1181 ( 
.A1(n_1167),
.A2(n_90),
.B(n_91),
.Y(n_1181)
);

XNOR2xp5_ASAP7_75t_L g1182 ( 
.A(n_1177),
.B(n_95),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1180),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1176),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1170),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1174),
.B(n_98),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1175),
.Y(n_1187)
);

AOI221xp5_ASAP7_75t_L g1188 ( 
.A1(n_1173),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.C(n_105),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1179),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1172),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1187),
.A2(n_1190),
.B1(n_1184),
.B2(n_1183),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1182),
.A2(n_1181),
.B(n_1178),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1188),
.A2(n_1181),
.B(n_1171),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_R g1194 ( 
.A1(n_1189),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_1194)
);

OAI321xp33_ASAP7_75t_L g1195 ( 
.A1(n_1186),
.A2(n_112),
.A3(n_113),
.B1(n_115),
.B2(n_116),
.C(n_117),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1185),
.Y(n_1196)
);

AOI222xp33_ASAP7_75t_L g1197 ( 
.A1(n_1187),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.C1(n_123),
.C2(n_124),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1191),
.B(n_127),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1196),
.A2(n_1192),
.B(n_1193),
.Y(n_1199)
);

OR2x2_ASAP7_75t_L g1200 ( 
.A(n_1194),
.B(n_128),
.Y(n_1200)
);

AOI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1199),
.A2(n_1197),
.B1(n_1195),
.B2(n_134),
.Y(n_1201)
);

AOI21xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1201),
.A2(n_1200),
.B(n_1198),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1202),
.A2(n_982),
.B(n_132),
.Y(n_1203)
);

OAI221xp5_ASAP7_75t_R g1204 ( 
.A1(n_1203),
.A2(n_129),
.B1(n_135),
.B2(n_138),
.C(n_139),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1204),
.A2(n_964),
.B(n_141),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1205),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_1206)
);

AOI211xp5_ASAP7_75t_L g1207 ( 
.A1(n_1206),
.A2(n_144),
.B(n_145),
.C(n_146),
.Y(n_1207)
);

AOI211xp5_ASAP7_75t_L g1208 ( 
.A1(n_1207),
.A2(n_888),
.B(n_147),
.C(n_148),
.Y(n_1208)
);


endmodule