module fake_jpeg_16278_n_270 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_1),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_33),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_49),
.Y(n_78)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_65),
.Y(n_92)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_31),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_20),
.B1(n_23),
.B2(n_32),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_74),
.B1(n_29),
.B2(n_19),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_23),
.B1(n_20),
.B2(n_28),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_47),
.B1(n_41),
.B2(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_70),
.Y(n_93)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_37),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_44),
.Y(n_108)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_76),
.A2(n_55),
.B1(n_44),
.B2(n_60),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_36),
.B(n_39),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_97),
.B(n_24),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_17),
.B(n_19),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_47),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_95),
.C(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_50),
.B(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_34),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_94),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_56),
.B1(n_75),
.B2(n_72),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_34),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_35),
.C(n_34),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_21),
.B(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_104),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_35),
.C(n_34),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_41),
.B1(n_44),
.B2(n_40),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_70),
.B1(n_49),
.B2(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_21),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_31),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_51),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_105),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_31),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

AOI22x1_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_53),
.B1(n_62),
.B2(n_44),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_114),
.B1(n_116),
.B2(n_127),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_124),
.B(n_130),
.Y(n_151)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_117),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_122),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_125),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_62),
.B1(n_32),
.B2(n_30),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_121),
.A2(n_22),
.B1(n_76),
.B2(n_104),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_77),
.B(n_25),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_1),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_17),
.B(n_30),
.C(n_29),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_1),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_80),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_133),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_93),
.B(n_27),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_134),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_78),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_95),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_86),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_94),
.B1(n_90),
.B2(n_100),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_152),
.B1(n_159),
.B2(n_161),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_86),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_87),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_160),
.B(n_124),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_154),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_100),
.B1(n_83),
.B2(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_101),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_156),
.B1(n_116),
.B2(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_109),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_81),
.B1(n_98),
.B2(n_102),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_109),
.A2(n_82),
.B(n_81),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_129),
.A2(n_82),
.B1(n_79),
.B2(n_85),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_112),
.B(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_79),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_144),
.B(n_162),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_186),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_120),
.B(n_125),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_173),
.B(n_178),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_131),
.B1(n_118),
.B2(n_121),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_174),
.B1(n_150),
.B2(n_160),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_122),
.B(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_177),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_130),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_152),
.Y(n_201)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_35),
.Y(n_186)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

BUFx4f_ASAP7_75t_SL g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_151),
.A2(n_26),
.B(n_3),
.C(n_5),
.D(n_6),
.Y(n_189)
);

AOI221xp5_ASAP7_75t_L g209 ( 
.A1(n_189),
.A2(n_171),
.B1(n_167),
.B2(n_155),
.C(n_138),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_196),
.B1(n_177),
.B2(n_181),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_140),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_203),
.C(n_204),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_157),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_176),
.Y(n_223)
);

OAI321xp33_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_209),
.A3(n_179),
.B1(n_173),
.B2(n_168),
.C(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_147),
.C(n_151),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_161),
.C(n_159),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_180),
.C(n_184),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_150),
.C(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_211),
.B(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_216),
.A2(n_218),
.B1(n_201),
.B2(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_204),
.A2(n_172),
.B1(n_205),
.B2(n_207),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_225),
.B1(n_182),
.B2(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_165),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.C(n_226),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_183),
.C(n_166),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_203),
.C(n_202),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_229),
.C(n_234),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_192),
.C(n_207),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_169),
.B1(n_199),
.B2(n_5),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_210),
.C(n_197),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_196),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_239),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_226),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_218),
.B(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_233),
.A2(n_175),
.B(n_169),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_248),
.Y(n_253)
);

NOR4xp25_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_210),
.C(n_223),
.D(n_189),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_244),
.A2(n_228),
.A3(n_231),
.B1(n_199),
.B2(n_13),
.C1(n_15),
.C2(n_16),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_238),
.C(n_229),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_14),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_239),
.B1(n_235),
.B2(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_246),
.B1(n_245),
.B2(n_7),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_245),
.B1(n_3),
.B2(n_7),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_15),
.A3(n_14),
.B1(n_85),
.B2(n_8),
.C1(n_9),
.C2(n_2),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_261),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_252),
.C(n_254),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_264),
.B(n_265),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_260),
.A2(n_256),
.B(n_250),
.Y(n_264)
);

AOI321xp33_ASAP7_75t_L g266 ( 
.A1(n_263),
.A2(n_252),
.A3(n_3),
.B1(n_8),
.B2(n_10),
.C(n_12),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_267),
.B1(n_2),
.B2(n_8),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_12),
.Y(n_269)
);


endmodule