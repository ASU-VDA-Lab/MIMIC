module real_jpeg_5233_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_1),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_1),
.A2(n_135),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_1),
.A2(n_135),
.B1(n_275),
.B2(n_280),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_1),
.A2(n_135),
.B1(n_378),
.B2(n_380),
.Y(n_377)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_2),
.A2(n_65),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_2),
.A2(n_65),
.B1(n_238),
.B2(n_242),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_3),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_4),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_4),
.A2(n_72),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_153),
.B1(n_199),
.B2(n_214),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_5),
.A2(n_153),
.B1(n_275),
.B2(n_280),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_5),
.A2(n_153),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_6),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_6),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_6),
.A2(n_85),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_9),
.Y(n_307)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_9),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_9),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_10),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_10),
.A2(n_120),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_10),
.A2(n_53),
.B1(n_120),
.B2(n_263),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_10),
.A2(n_120),
.B1(n_284),
.B2(n_288),
.Y(n_283)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_13),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_13),
.A2(n_202),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_13),
.B(n_270),
.C(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_13),
.B(n_110),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_13),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_13),
.B(n_61),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_13),
.B(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_14),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_14),
.Y(n_195)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_16),
.A2(n_53),
.B1(n_56),
.B2(n_59),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_16),
.A2(n_59),
.B1(n_124),
.B2(n_128),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_16),
.A2(n_59),
.B1(n_352),
.B2(n_354),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_248),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_247),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_218),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_21),
.B(n_218),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_159),
.C(n_177),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_22),
.A2(n_23),
.B1(n_159),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_89),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_24),
.B(n_90),
.C(n_158),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_66),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_25),
.B(n_66),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_52),
.B1(n_60),
.B2(n_62),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_26),
.A2(n_257),
.B(n_261),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_26),
.A2(n_60),
.B1(n_292),
.B2(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_26),
.A2(n_261),
.B(n_333),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_27),
.A2(n_61),
.B1(n_63),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_27),
.A2(n_61),
.B1(n_161),
.B2(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_27),
.B(n_262),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_42),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_40),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_31),
.Y(n_226)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_31),
.Y(n_268)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_31),
.Y(n_294)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_32),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_32),
.Y(n_335)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_33),
.Y(n_163)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_33),
.Y(n_340)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_41),
.Y(n_296)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_42),
.A2(n_292),
.B(n_297),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_44),
.Y(n_270)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_47),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_47),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_48),
.Y(n_209)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g353 ( 
.A(n_49),
.Y(n_353)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_52),
.A2(n_60),
.B(n_297),
.Y(n_406)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_58),
.Y(n_228)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_61),
.B(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_77),
.B1(n_82),
.B2(n_87),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_67),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_75),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_76),
.Y(n_279)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_77),
.B(n_283),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_77),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_77),
.A2(n_206),
.B1(n_351),
.B2(n_386),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_83),
.A2(n_167),
.B1(n_168),
.B2(n_171),
.Y(n_166)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_88),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_131),
.B1(n_157),
.B2(n_158),
.Y(n_89)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

AOI22x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_110),
.B1(n_117),
.B2(n_122),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_91),
.A2(n_212),
.B(n_216),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_91),
.A2(n_216),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_91),
.B(n_117),
.Y(n_382)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_92),
.A2(n_123),
.B1(n_217),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_92),
.A2(n_213),
.B1(n_217),
.B2(n_377),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_110),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_102),
.B2(n_107),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_95),
.Y(n_361)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_96),
.Y(n_366)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_100),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_100),
.Y(n_347)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_100),
.Y(n_381)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_110),
.Y(n_217)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_110)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_114),
.Y(n_165)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_116),
.Y(n_259)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_118),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g358 ( 
.A1(n_128),
.A2(n_227),
.A3(n_345),
.B1(n_359),
.B2(n_362),
.Y(n_358)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_137),
.B1(n_145),
.B2(n_151),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_180),
.B(n_182),
.Y(n_179)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_137),
.A2(n_151),
.B(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_138),
.A2(n_402),
.B(n_403),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_145),
.B(n_202),
.Y(n_384)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_190),
.A3(n_194),
.B1(n_196),
.B2(n_201),
.Y(n_189)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_159),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_160),
.B(n_166),
.Y(n_234)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_167),
.A2(n_168),
.B1(n_205),
.B2(n_210),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_167),
.A2(n_171),
.B(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_167),
.A2(n_274),
.B(n_282),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_167),
.A2(n_202),
.B(n_282),
.Y(n_308)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_169),
.B(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_176),
.Y(n_281)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_176),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_177),
.B(n_421),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_188),
.C(n_211),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_178),
.A2(n_179),
.B1(n_211),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_181),
.B(n_183),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_202),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_SL g402 ( 
.A1(n_184),
.A2(n_201),
.B(n_202),
.Y(n_402)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_188),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_203),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_189),
.A2(n_203),
.B1(n_204),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_189),
.Y(n_395)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_200),
.Y(n_379)
);

OAI21xp33_ASAP7_75t_SL g343 ( 
.A1(n_202),
.A2(n_239),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_211),
.Y(n_416)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_217),
.A2(n_377),
.B(n_382),
.Y(n_376)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_218),
.Y(n_431)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_220),
.CI(n_233),
.CON(n_218),
.SN(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_229),
.B2(n_232),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_229),
.Y(n_232)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_246),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_409),
.B(n_428),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_390),
.B(n_408),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_368),
.B(n_389),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_327),
.B(n_367),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_300),
.B(n_326),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_272),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_255),
.B(n_272),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_256),
.A2(n_265),
.B1(n_266),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_260),
.Y(n_264)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_289),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_290),
.C(n_299),
.Y(n_328)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_298),
.B2(n_299),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_293),
.Y(n_363)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_316),
.B(n_325),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_309),
.B(n_315),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_314),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_311),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_350),
.B(n_355),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_323),
.Y(n_325)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_329),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_348),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_341),
.B2(n_342),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_341),
.C(n_348),
.Y(n_369)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx5_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx6_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_358),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_349),
.B(n_358),
.Y(n_374)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_SL g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_369),
.B(n_370),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_372),
.B1(n_375),
.B2(n_388),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_374),
.C(n_388),
.Y(n_391)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_375),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_383),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_376),
.B(n_384),
.C(n_385),
.Y(n_396)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_392),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_391),
.B(n_392),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_399),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_396),
.B1(n_397),
.B2(n_398),
.Y(n_393)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_396),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_396),
.B(n_397),
.C(n_399),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_404),
.B2(n_407),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_400),
.B(n_405),
.C(n_406),
.Y(n_419)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_404),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_423),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_412),
.A2(n_429),
.B(n_430),
.Y(n_428)
);

NOR2x1_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_420),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_420),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.C(n_419),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_414),
.B(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_419),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_425),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_425),
.Y(n_429)
);


endmodule