module fake_netlist_1_2169_n_44 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_44);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_44;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_13;
wire n_25;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_7), .Y(n_11) );
CKINVDCx16_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_11), .B(n_0), .Y(n_20) );
OAI22xp33_ASAP7_75t_L g21 ( .A1(n_12), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_11), .B(n_1), .Y(n_22) );
INVxp33_ASAP7_75t_SL g23 ( .A(n_16), .Y(n_23) );
OAI221xp5_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_22), .B1(n_18), .B2(n_13), .C(n_19), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_18), .B(n_17), .Y(n_25) );
OAI221xp5_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_16), .B1(n_17), .B2(n_15), .C(n_5), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_19), .Y(n_27) );
OAI211xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_22), .B(n_19), .C(n_23), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_21), .B1(n_19), .B2(n_4), .Y(n_29) );
NAND3xp33_ASAP7_75t_L g30 ( .A(n_24), .B(n_2), .C(n_3), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_29), .B(n_25), .Y(n_32) );
INVx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
NOR2x1_ASAP7_75t_L g36 ( .A(n_34), .B(n_28), .Y(n_36) );
OAI22xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_27), .B1(n_25), .B2(n_8), .Y(n_37) );
AOI221xp5_ASAP7_75t_L g38 ( .A1(n_35), .A2(n_27), .B1(n_5), .B2(n_8), .C(n_9), .Y(n_38) );
INVxp67_ASAP7_75t_L g39 ( .A(n_36), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_37), .Y(n_40) );
INVx2_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
AOI22xp33_ASAP7_75t_L g43 ( .A1(n_41), .A2(n_4), .B1(n_33), .B2(n_40), .Y(n_43) );
AOI22xp5_ASAP7_75t_SL g44 ( .A1(n_42), .A2(n_33), .B1(n_41), .B2(n_43), .Y(n_44) );
endmodule