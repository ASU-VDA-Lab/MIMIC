module real_aes_7145_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g553 ( .A1(n_0), .A2(n_160), .B(n_554), .C(n_557), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_1), .B(n_498), .Y(n_558) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
INVx1_ASAP7_75t_L g194 ( .A(n_3), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_4), .B(n_152), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_5), .A2(n_467), .B(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_6), .A2(n_137), .B(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_7), .A2(n_35), .B1(n_146), .B2(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_8), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_9), .B(n_137), .Y(n_163) );
AND2x6_ASAP7_75t_L g161 ( .A(n_10), .B(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_11), .A2(n_161), .B(n_457), .C(n_459), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_12), .B(n_36), .Y(n_117) );
INVx1_ASAP7_75t_L g142 ( .A(n_13), .Y(n_142) );
INVx1_ASAP7_75t_L g187 ( .A(n_14), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_15), .B(n_150), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_16), .B(n_152), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_17), .B(n_138), .Y(n_199) );
AO32x2_ASAP7_75t_L g221 ( .A1(n_18), .A2(n_137), .A3(n_167), .B1(n_178), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_19), .B(n_146), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_20), .B(n_138), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_21), .A2(n_54), .B1(n_146), .B2(n_224), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g246 ( .A1(n_22), .A2(n_82), .B1(n_146), .B2(n_150), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_23), .B(n_146), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_24), .A2(n_178), .B(n_457), .C(n_518), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g485 ( .A1(n_25), .A2(n_178), .B(n_457), .C(n_486), .Y(n_485) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_26), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_27), .B(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_28), .A2(n_467), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_29), .B(n_180), .Y(n_218) );
INVx2_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_31), .A2(n_469), .B(n_477), .C(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_32), .B(n_146), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_33), .B(n_180), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_34), .B(n_232), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_37), .B(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_38), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_39), .A2(n_78), .B1(n_122), .B2(n_123), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_39), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_40), .B(n_152), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_41), .B(n_467), .Y(n_484) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_42), .A2(n_79), .B1(n_440), .B2(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_42), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_43), .A2(n_469), .B(n_471), .C(n_477), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_44), .A2(n_121), .B1(n_124), .B2(n_125), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_44), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_45), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g555 ( .A(n_46), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_47), .A2(n_91), .B1(n_224), .B2(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g472 ( .A(n_48), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_49), .B(n_146), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_50), .B(n_146), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_51), .B(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_51), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_52), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_53), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_SL g203 ( .A1(n_55), .A2(n_59), .B1(n_146), .B2(n_150), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_56), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_57), .B(n_146), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_58), .B(n_146), .Y(n_229) );
INVx1_ASAP7_75t_L g162 ( .A(n_60), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_61), .B(n_467), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_62), .B(n_498), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_63), .A2(n_158), .B(n_190), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_64), .B(n_146), .Y(n_195) );
INVx1_ASAP7_75t_L g141 ( .A(n_65), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_66), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_67), .B(n_152), .Y(n_508) );
AO32x2_ASAP7_75t_L g242 ( .A1(n_68), .A2(n_137), .A3(n_178), .B1(n_243), .B2(n_247), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_69), .B(n_153), .Y(n_460) );
INVx1_ASAP7_75t_L g173 ( .A(n_70), .Y(n_173) );
INVx1_ASAP7_75t_L g213 ( .A(n_71), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_72), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_73), .B(n_474), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_74), .A2(n_457), .B(n_477), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_75), .B(n_150), .Y(n_214) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_76), .Y(n_493) );
INVx1_ASAP7_75t_L g109 ( .A(n_77), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_78), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_79), .A2(n_129), .B1(n_439), .B2(n_440), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_79), .Y(n_440) );
AOI222xp33_ASAP7_75t_SL g103 ( .A1(n_80), .A2(n_104), .B1(n_118), .B2(n_740), .C1(n_745), .C2(n_764), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_80), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_81), .B(n_473), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_83), .B(n_224), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_84), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_85), .B(n_150), .Y(n_217) );
INVx2_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_87), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_88), .B(n_177), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_89), .B(n_150), .Y(n_149) );
OR2x2_ASAP7_75t_L g113 ( .A(n_90), .B(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g443 ( .A(n_90), .B(n_115), .Y(n_443) );
INVx2_ASAP7_75t_L g731 ( .A(n_90), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_92), .A2(n_102), .B1(n_150), .B2(n_151), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_93), .B(n_467), .Y(n_504) );
INVx1_ASAP7_75t_L g507 ( .A(n_94), .Y(n_507) );
INVxp67_ASAP7_75t_L g496 ( .A(n_95), .Y(n_496) );
AOI222xp33_ASAP7_75t_SL g119 ( .A1(n_96), .A2(n_120), .B1(n_126), .B2(n_732), .C1(n_733), .C2(n_737), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_97), .B(n_150), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_98), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g453 ( .A(n_99), .Y(n_453) );
INVx1_ASAP7_75t_L g531 ( .A(n_100), .Y(n_531) );
AND2x2_ASAP7_75t_L g479 ( .A(n_101), .B(n_180), .Y(n_479) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
NOR2xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_110), .Y(n_107) );
INVx1_ASAP7_75t_SL g744 ( .A(n_108), .Y(n_744) );
INVx1_ASAP7_75t_L g743 ( .A(n_110), .Y(n_743) );
OA21x2_ASAP7_75t_L g765 ( .A1(n_110), .A2(n_744), .B(n_762), .Y(n_765) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
AOI211xp5_ASAP7_75t_L g758 ( .A1(n_112), .A2(n_757), .B(n_759), .C(n_760), .Y(n_758) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g756 ( .A(n_113), .Y(n_756) );
BUFx2_ASAP7_75t_L g762 ( .A(n_113), .Y(n_762) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_114), .B(n_731), .Y(n_739) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g730 ( .A(n_115), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
INVxp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g732 ( .A(n_120), .Y(n_732) );
INVx1_ASAP7_75t_L g124 ( .A(n_121), .Y(n_124) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_441), .B1(n_444), .B2(n_728), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g733 ( .A1(n_128), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
INVx2_ASAP7_75t_L g439 ( .A(n_129), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_129), .A2(n_439), .B1(n_750), .B2(n_751), .Y(n_749) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_130), .B(n_363), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_321), .Y(n_130) );
NOR4xp25_ASAP7_75t_L g131 ( .A(n_132), .B(n_261), .C(n_297), .D(n_311), .Y(n_131) );
OAI221xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_205), .B1(n_237), .B2(n_248), .C(n_252), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_133), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_181), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_164), .Y(n_135) );
AND2x2_ASAP7_75t_L g258 ( .A(n_136), .B(n_165), .Y(n_258) );
INVx3_ASAP7_75t_L g266 ( .A(n_136), .Y(n_266) );
AND2x2_ASAP7_75t_L g320 ( .A(n_136), .B(n_184), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_136), .B(n_183), .Y(n_356) );
AND2x2_ASAP7_75t_L g414 ( .A(n_136), .B(n_276), .Y(n_414) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_163), .Y(n_136) );
INVx4_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_137), .A2(n_484), .B(n_485), .Y(n_483) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_137), .Y(n_490) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g167 ( .A(n_138), .Y(n_167) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_139), .B(n_140), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_155), .B(n_161), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B(n_152), .Y(n_144) );
INVx3_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_146), .Y(n_533) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g224 ( .A(n_147), .Y(n_224) );
BUFx3_ASAP7_75t_L g245 ( .A(n_147), .Y(n_245) );
AND2x6_ASAP7_75t_L g457 ( .A(n_147), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx2_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_152), .A2(n_170), .B(n_171), .Y(n_169) );
O2A1O1Ixp5_ASAP7_75t_SL g211 ( .A1(n_152), .A2(n_212), .B(n_213), .C(n_214), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_152), .B(n_496), .Y(n_495) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g243 ( .A1(n_153), .A2(n_177), .B1(n_244), .B2(n_246), .Y(n_243) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
INVx1_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
AND2x2_ASAP7_75t_L g455 ( .A(n_154), .B(n_159), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_154), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .Y(n_155) );
INVx2_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_160), .A2(n_174), .B(n_194), .C(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_160), .A2(n_177), .B1(n_202), .B2(n_203), .Y(n_201) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_160), .A2(n_177), .B1(n_223), .B2(n_225), .Y(n_222) );
BUFx3_ASAP7_75t_L g178 ( .A(n_161), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_161), .A2(n_186), .B(n_193), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_211), .B(n_215), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_161), .A2(n_228), .B(n_233), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g454 ( .A(n_161), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g467 ( .A(n_161), .B(n_455), .Y(n_467) );
INVx4_ASAP7_75t_SL g478 ( .A(n_161), .Y(n_478) );
AND2x2_ASAP7_75t_L g249 ( .A(n_164), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g263 ( .A(n_164), .B(n_184), .Y(n_263) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_165), .B(n_184), .Y(n_278) );
AND2x2_ASAP7_75t_L g290 ( .A(n_165), .B(n_266), .Y(n_290) );
OR2x2_ASAP7_75t_L g292 ( .A(n_165), .B(n_250), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_165), .B(n_250), .Y(n_327) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_165), .Y(n_372) );
INVx1_ASAP7_75t_L g380 ( .A(n_165), .Y(n_380) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_179), .Y(n_165) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_166), .A2(n_185), .B(n_196), .Y(n_184) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_167), .B(n_463), .Y(n_462) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_178), .Y(n_168) );
O2A1O1Ixp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .C(n_176), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_174), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_176), .A2(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g556 ( .A(n_177), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_178), .B(n_201), .C(n_204), .Y(n_200) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_180), .A2(n_210), .B(n_218), .Y(n_209) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_180), .A2(n_227), .B(n_236), .Y(n_226) );
INVx2_ASAP7_75t_L g247 ( .A(n_180), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_180), .A2(n_466), .B(n_468), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_180), .A2(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g524 ( .A(n_180), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g297 ( .A1(n_181), .A2(n_298), .B1(n_302), .B2(n_306), .C(n_307), .Y(n_297) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g257 ( .A(n_182), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_197), .Y(n_182) );
INVx2_ASAP7_75t_L g256 ( .A(n_183), .Y(n_256) );
AND2x2_ASAP7_75t_L g309 ( .A(n_183), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g328 ( .A(n_183), .B(n_266), .Y(n_328) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g391 ( .A(n_184), .B(n_266), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .C(n_190), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_188), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_188), .A2(n_487), .B(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_190), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_191), .A2(n_216), .B(n_217), .Y(n_215) );
INVx4_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g474 ( .A(n_192), .Y(n_474) );
AND2x2_ASAP7_75t_L g313 ( .A(n_197), .B(n_258), .Y(n_313) );
OAI322xp33_ASAP7_75t_L g381 ( .A1(n_197), .A2(n_337), .A3(n_382), .B1(n_384), .B2(n_387), .C1(n_389), .C2(n_393), .Y(n_381) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2x1_ASAP7_75t_L g264 ( .A(n_198), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g277 ( .A(n_198), .Y(n_277) );
AND2x2_ASAP7_75t_L g386 ( .A(n_198), .B(n_266), .Y(n_386) );
AND2x2_ASAP7_75t_L g418 ( .A(n_198), .B(n_290), .Y(n_418) );
OR2x2_ASAP7_75t_L g421 ( .A(n_198), .B(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
INVx1_ASAP7_75t_L g251 ( .A(n_199), .Y(n_251) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_201), .A2(n_204), .B(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g451 ( .A1(n_204), .A2(n_452), .B(n_462), .Y(n_451) );
INVx3_ASAP7_75t_L g498 ( .A(n_204), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_204), .B(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g527 ( .A1(n_204), .A2(n_528), .B(n_535), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_204), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_219), .Y(n_206) );
INVx1_ASAP7_75t_L g434 ( .A(n_207), .Y(n_434) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g239 ( .A(n_208), .B(n_226), .Y(n_239) );
INVx2_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g296 ( .A(n_209), .Y(n_296) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_209), .Y(n_304) );
OR2x2_ASAP7_75t_L g428 ( .A(n_209), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g253 ( .A(n_219), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g293 ( .A(n_219), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g345 ( .A(n_219), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_226), .Y(n_219) );
AND2x2_ASAP7_75t_L g240 ( .A(n_220), .B(n_241), .Y(n_240) );
NOR2xp67_ASAP7_75t_L g300 ( .A(n_220), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g354 ( .A(n_220), .B(n_242), .Y(n_354) );
OR2x2_ASAP7_75t_L g362 ( .A(n_220), .B(n_296), .Y(n_362) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
BUFx2_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
AND2x2_ASAP7_75t_L g281 ( .A(n_221), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g305 ( .A(n_221), .B(n_226), .Y(n_305) );
AND2x2_ASAP7_75t_L g369 ( .A(n_221), .B(n_242), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_226), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_226), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g282 ( .A(n_226), .Y(n_282) );
INVx1_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
AND2x2_ASAP7_75t_L g299 ( .A(n_226), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_226), .Y(n_377) );
INVx1_ASAP7_75t_L g429 ( .A(n_226), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_240), .Y(n_237) );
AND2x2_ASAP7_75t_L g406 ( .A(n_238), .B(n_315), .Y(n_406) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g333 ( .A(n_240), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g432 ( .A(n_240), .B(n_367), .Y(n_432) );
INVx1_ASAP7_75t_L g254 ( .A(n_241), .Y(n_254) );
AND2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_274), .Y(n_280) );
BUFx2_ASAP7_75t_L g339 ( .A(n_241), .Y(n_339) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_242), .Y(n_260) );
INVx1_ASAP7_75t_L g270 ( .A(n_242), .Y(n_270) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_245), .Y(n_476) );
INVx2_ASAP7_75t_L g557 ( .A(n_245), .Y(n_557) );
INVx1_ASAP7_75t_L g521 ( .A(n_247), .Y(n_521) );
NOR2xp67_ASAP7_75t_L g408 ( .A(n_248), .B(n_255), .Y(n_408) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI32xp33_ASAP7_75t_L g252 ( .A1(n_249), .A2(n_253), .A3(n_255), .B1(n_257), .B2(n_259), .Y(n_252) );
AND2x2_ASAP7_75t_L g392 ( .A(n_249), .B(n_265), .Y(n_392) );
AND2x2_ASAP7_75t_L g430 ( .A(n_249), .B(n_328), .Y(n_430) );
INVx1_ASAP7_75t_L g310 ( .A(n_250), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_254), .B(n_316), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_255), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_255), .B(n_258), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_255), .B(n_327), .Y(n_409) );
OR2x2_ASAP7_75t_L g423 ( .A(n_255), .B(n_292), .Y(n_423) );
INVx3_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g350 ( .A(n_256), .B(n_258), .Y(n_350) );
OR2x2_ASAP7_75t_L g359 ( .A(n_256), .B(n_346), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_258), .B(n_309), .Y(n_331) );
INVx2_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
OR2x2_ASAP7_75t_L g361 ( .A(n_260), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g376 ( .A(n_260), .B(n_377), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_260), .A2(n_353), .B(n_434), .C(n_435), .Y(n_433) );
OAI321xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_267), .A3(n_272), .B1(n_275), .B2(n_279), .C(n_283), .Y(n_261) );
INVx1_ASAP7_75t_L g374 ( .A(n_262), .Y(n_374) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
AND2x2_ASAP7_75t_L g385 ( .A(n_263), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g337 ( .A(n_265), .Y(n_337) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_266), .B(n_380), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_267), .A2(n_405), .B1(n_407), .B2(n_409), .C(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g342 ( .A(n_269), .B(n_316), .Y(n_342) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_270), .B(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_272), .A2(n_313), .B(n_358), .C(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g324 ( .A(n_274), .B(n_281), .Y(n_324) );
BUFx2_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
INVx1_ASAP7_75t_L g349 ( .A(n_274), .Y(n_349) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OR2x2_ASAP7_75t_L g355 ( .A(n_277), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g438 ( .A(n_277), .Y(n_438) );
INVx1_ASAP7_75t_L g431 ( .A(n_278), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AND2x2_ASAP7_75t_L g284 ( .A(n_280), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g388 ( .A(n_280), .B(n_305), .Y(n_388) );
INVx1_ASAP7_75t_L g317 ( .A(n_281), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B1(n_291), .B2(n_293), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_285), .B(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g353 ( .A(n_286), .B(n_354), .Y(n_353) );
BUFx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_SL g316 ( .A(n_287), .B(n_296), .Y(n_316) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g308 ( .A(n_290), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g318 ( .A(n_292), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_295), .A2(n_413), .B1(n_415), .B2(n_416), .C(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g301 ( .A(n_296), .Y(n_301) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_296), .Y(n_367) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_299), .B(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_300), .A2(n_305), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_303), .B(n_313), .Y(n_410) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g379 ( .A(n_304), .Y(n_379) );
AND2x2_ASAP7_75t_L g338 ( .A(n_305), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g427 ( .A(n_305), .Y(n_427) );
INVx1_ASAP7_75t_L g343 ( .A(n_308), .Y(n_343) );
INVx1_ASAP7_75t_L g398 ( .A(n_309), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B1(n_317), .B2(n_318), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_315), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g383 ( .A(n_316), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_316), .B(n_354), .Y(n_420) );
OR2x2_ASAP7_75t_L g393 ( .A(n_317), .B(n_346), .Y(n_393) );
INVx1_ASAP7_75t_L g332 ( .A(n_318), .Y(n_332) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_320), .B(n_371), .Y(n_370) );
NOR3xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_340), .C(n_351), .Y(n_321) );
OAI211xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_325), .B(n_329), .C(n_335), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_324), .A2(n_395), .B1(n_399), .B2(n_402), .C(n_404), .Y(n_394) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g336 ( .A(n_327), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_391), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_328), .A2(n_376), .B(n_378), .C(n_380), .Y(n_375) );
INVx2_ASAP7_75t_L g422 ( .A(n_328), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_332), .B(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g401 ( .A(n_334), .B(n_354), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
OAI21xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_343), .B(n_344), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI21xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_347), .B(n_350), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_345), .B(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_350), .B(n_437), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_355), .B(n_357), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g378 ( .A(n_354), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND4x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_394), .C(n_411), .D(n_433), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_381), .Y(n_364) );
OAI211xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_370), .B(n_373), .C(n_375), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_369), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_380), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVx1_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
INVx2_ASAP7_75t_SL g403 ( .A(n_391), .Y(n_403) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g416 ( .A(n_401), .Y(n_416) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_419), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OAI221xp5_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_421), .B1(n_423), .B2(n_424), .C(n_425), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B1(n_431), .B2(n_432), .Y(n_425) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g734 ( .A(n_442), .Y(n_734) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g735 ( .A(n_444), .Y(n_735) );
OR3x1_ASAP7_75t_L g444 ( .A(n_445), .B(n_626), .C(n_691), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g445 ( .A(n_446), .B(n_567), .C(n_593), .D(n_616), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_499), .B1(n_537), .B2(n_544), .C(n_559), .Y(n_446) );
CKINVDCx14_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_448), .A2(n_560), .B1(n_584), .B2(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_480), .Y(n_448) );
INVx1_ASAP7_75t_SL g620 ( .A(n_449), .Y(n_620) );
OR2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_464), .Y(n_449) );
OR2x2_ASAP7_75t_L g542 ( .A(n_450), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g562 ( .A(n_450), .B(n_481), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_450), .B(n_489), .Y(n_575) );
AND2x2_ASAP7_75t_L g592 ( .A(n_450), .B(n_464), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_450), .B(n_540), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_450), .B(n_591), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_450), .B(n_480), .Y(n_713) );
AOI211xp5_ASAP7_75t_SL g724 ( .A1(n_450), .A2(n_630), .B(n_725), .C(n_726), .Y(n_724) );
INVx5_ASAP7_75t_SL g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_451), .B(n_481), .Y(n_596) );
AND2x2_ASAP7_75t_L g599 ( .A(n_451), .B(n_482), .Y(n_599) );
OR2x2_ASAP7_75t_L g644 ( .A(n_451), .B(n_481), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_451), .B(n_489), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B(n_456), .Y(n_452) );
INVx5_ASAP7_75t_L g470 ( .A(n_457), .Y(n_470) );
INVx5_ASAP7_75t_SL g543 ( .A(n_464), .Y(n_543) );
AND2x2_ASAP7_75t_L g561 ( .A(n_464), .B(n_562), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_464), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g647 ( .A(n_464), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g679 ( .A(n_464), .B(n_489), .Y(n_679) );
OR2x2_ASAP7_75t_L g685 ( .A(n_464), .B(n_575), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_464), .B(n_635), .Y(n_694) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_479), .Y(n_464) );
BUFx2_ASAP7_75t_L g516 ( .A(n_467), .Y(n_516) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_470), .A2(n_478), .B(n_493), .C(n_494), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_SL g551 ( .A1(n_470), .A2(n_478), .B(n_552), .C(n_553), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_475), .C(n_476), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g506 ( .A1(n_473), .A2(n_476), .B(n_507), .C(n_508), .Y(n_506) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
AND2x2_ASAP7_75t_L g576 ( .A(n_481), .B(n_543), .Y(n_576) );
INVx1_ASAP7_75t_SL g589 ( .A(n_481), .Y(n_589) );
OR2x2_ASAP7_75t_L g624 ( .A(n_481), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g630 ( .A(n_481), .B(n_489), .Y(n_630) );
AND2x2_ASAP7_75t_L g688 ( .A(n_481), .B(n_540), .Y(n_688) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_482), .B(n_543), .Y(n_615) );
INVx3_ASAP7_75t_L g540 ( .A(n_489), .Y(n_540) );
OR2x2_ASAP7_75t_L g581 ( .A(n_489), .B(n_543), .Y(n_581) );
AND2x2_ASAP7_75t_L g591 ( .A(n_489), .B(n_589), .Y(n_591) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_489), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_489), .B(n_562), .Y(n_648) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_497), .Y(n_489) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_498), .A2(n_550), .B(n_558), .Y(n_549) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_499), .A2(n_665), .B1(n_667), .B2(n_669), .C(n_672), .Y(n_664) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_511), .Y(n_500) );
AND2x2_ASAP7_75t_L g638 ( .A(n_501), .B(n_619), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_501), .B(n_697), .Y(n_701) );
OR2x2_ASAP7_75t_L g722 ( .A(n_501), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_501), .B(n_727), .Y(n_726) );
BUFx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx5_ASAP7_75t_L g569 ( .A(n_502), .Y(n_569) );
AND2x2_ASAP7_75t_L g646 ( .A(n_502), .B(n_513), .Y(n_646) );
AND2x2_ASAP7_75t_L g707 ( .A(n_502), .B(n_586), .Y(n_707) );
AND2x2_ASAP7_75t_L g720 ( .A(n_502), .B(n_540), .Y(n_720) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_509), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_512), .B(n_525), .Y(n_511) );
AND2x4_ASAP7_75t_L g547 ( .A(n_512), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g565 ( .A(n_512), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g572 ( .A(n_512), .Y(n_572) );
AND2x2_ASAP7_75t_L g641 ( .A(n_512), .B(n_619), .Y(n_641) );
AND2x2_ASAP7_75t_L g651 ( .A(n_512), .B(n_569), .Y(n_651) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_512), .Y(n_659) );
AND2x2_ASAP7_75t_L g671 ( .A(n_512), .B(n_549), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_512), .B(n_603), .Y(n_675) );
AND2x2_ASAP7_75t_L g712 ( .A(n_512), .B(n_707), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_512), .B(n_586), .Y(n_723) );
OR2x2_ASAP7_75t_L g725 ( .A(n_512), .B(n_661), .Y(n_725) );
INVx5_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g611 ( .A(n_513), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g621 ( .A(n_513), .B(n_566), .Y(n_621) );
AND2x2_ASAP7_75t_L g633 ( .A(n_513), .B(n_549), .Y(n_633) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_513), .Y(n_663) );
AND2x4_ASAP7_75t_L g697 ( .A(n_513), .B(n_548), .Y(n_697) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_522), .Y(n_513) );
AOI21xp5_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_517), .B(n_521), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
BUFx2_ASAP7_75t_L g546 ( .A(n_525), .Y(n_546) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g586 ( .A(n_526), .Y(n_586) );
AND2x2_ASAP7_75t_L g619 ( .A(n_526), .B(n_549), .Y(n_619) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g566 ( .A(n_527), .B(n_549), .Y(n_566) );
BUFx2_ASAP7_75t_L g612 ( .A(n_527), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_534), .Y(n_528) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_539), .B(n_620), .Y(n_699) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_540), .B(n_562), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_540), .B(n_543), .Y(n_601) );
AND2x2_ASAP7_75t_L g656 ( .A(n_540), .B(n_592), .Y(n_656) );
AOI221xp5_ASAP7_75t_SL g593 ( .A1(n_541), .A2(n_594), .B1(n_602), .B2(n_604), .C(n_608), .Y(n_593) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g588 ( .A(n_542), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g629 ( .A(n_542), .B(n_630), .Y(n_629) );
OAI321xp33_ASAP7_75t_L g636 ( .A1(n_542), .A2(n_595), .A3(n_637), .B1(n_639), .B2(n_640), .C(n_642), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_543), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_546), .B(n_697), .Y(n_715) );
AND2x2_ASAP7_75t_L g602 ( .A(n_547), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_547), .B(n_606), .Y(n_605) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_548), .Y(n_578) );
AND2x2_ASAP7_75t_L g585 ( .A(n_548), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_548), .B(n_660), .Y(n_690) );
INVx1_ASAP7_75t_L g727 ( .A(n_548), .Y(n_727) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .B(n_564), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_561), .A2(n_671), .B(n_720), .C(n_721), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_562), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_562), .B(n_600), .Y(n_666) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g609 ( .A(n_566), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_566), .B(n_569), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_566), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_566), .B(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B1(n_582), .B2(n_587), .Y(n_567) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g583 ( .A(n_569), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g606 ( .A(n_569), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g618 ( .A(n_569), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_569), .B(n_612), .Y(n_654) );
OR2x2_ASAP7_75t_L g661 ( .A(n_569), .B(n_586), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_569), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g711 ( .A(n_569), .B(n_697), .Y(n_711) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_573), .B1(n_577), .B2(n_579), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g617 ( .A(n_572), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_575), .A2(n_590), .B1(n_658), .B2(n_662), .Y(n_657) );
INVx1_ASAP7_75t_L g705 ( .A(n_576), .Y(n_705) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_580), .A2(n_617), .B1(n_620), .B2(n_621), .C(n_622), .Y(n_616) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g595 ( .A(n_581), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_585), .B(n_651), .Y(n_683) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_586), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_586), .Y(n_607) );
NAND2xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g625 ( .A(n_592), .Y(n_625) );
AND2x2_ASAP7_75t_L g634 ( .A(n_592), .B(n_635), .Y(n_634) );
NAND2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_597), .Y(n_594) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
AND2x2_ASAP7_75t_L g678 ( .A(n_599), .B(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_602), .A2(n_628), .B1(n_631), .B2(n_634), .C(n_636), .Y(n_627) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_606), .B(n_663), .Y(n_662) );
AOI21xp33_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B(n_613), .Y(n_608) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_613), .Y(n_710) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OR2x2_ASAP7_75t_L g652 ( .A(n_615), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g673 ( .A(n_618), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_618), .B(n_678), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_621), .B(n_643), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_627), .B(n_645), .C(n_664), .D(n_677), .Y(n_626) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g635 ( .A(n_630), .Y(n_635) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g668 ( .A(n_639), .B(n_644), .Y(n_668) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI211xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_649), .C(n_657), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g716 ( .A1(n_647), .A2(n_689), .B(n_717), .C(n_724), .Y(n_716) );
INVx1_ASAP7_75t_SL g676 ( .A(n_648), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_654), .B2(n_655), .Y(n_649) );
INVx1_ASAP7_75t_L g680 ( .A(n_654), .Y(n_680) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_660), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_660), .B(n_671), .Y(n_704) );
INVx2_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g681 ( .A(n_671), .Y(n_681) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_676), .Y(n_672) );
INVxp33_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_680), .A3(n_681), .B1(n_682), .B2(n_684), .C1(n_686), .C2(n_689), .Y(n_677) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_709), .C(n_716), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .B1(n_698), .B2(n_700), .C(n_702), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_SL g708 ( .A(n_697), .Y(n_708) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_709) );
NAND2xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g736 ( .A(n_729), .Y(n_736) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVxp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI211xp5_ASAP7_75t_SL g746 ( .A1(n_747), .A2(n_757), .B(n_758), .C(n_761), .Y(n_746) );
NOR3xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_753), .C(n_756), .Y(n_747) );
INVxp67_ASAP7_75t_L g759 ( .A(n_748), .Y(n_759) );
INVx1_ASAP7_75t_L g755 ( .A(n_749), .Y(n_755) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_L g760 ( .A(n_753), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
NOR2xp33_ASAP7_75t_SL g761 ( .A(n_762), .B(n_763), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
endmodule