module fake_jpeg_1459_n_387 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_387);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_387;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_62),
.Y(n_103)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_47),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_49),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_15),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_9),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_56),
.B(n_59),
.Y(n_118)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_9),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_74),
.Y(n_113)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_8),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_68),
.B(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_1),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_1),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_73),
.A2(n_99),
.B(n_49),
.Y(n_145)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_21),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_77),
.A2(n_20),
.B1(n_43),
.B2(n_35),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_83),
.Y(n_121)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_81),
.B(n_86),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_40),
.B(n_8),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_88),
.B(n_91),
.Y(n_148)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_41),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_93),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_41),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_29),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_98),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_95),
.B(n_3),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_28),
.B(n_10),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_20),
.B(n_27),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_36),
.B1(n_25),
.B2(n_45),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_52),
.A2(n_27),
.B1(n_44),
.B2(n_43),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_108),
.A2(n_122),
.B1(n_139),
.B2(n_142),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_36),
.B1(n_45),
.B2(n_30),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_123),
.B1(n_129),
.B2(n_134),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_69),
.A2(n_44),
.B1(n_35),
.B2(n_32),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_119),
.A2(n_135),
.B1(n_150),
.B2(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_31),
.B1(n_30),
.B2(n_22),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_61),
.A2(n_32),
.B1(n_31),
.B2(n_22),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_73),
.B(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_11),
.C(n_12),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_133),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_12),
.B1(n_14),
.B2(n_5),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_71),
.A2(n_4),
.B1(n_6),
.B2(n_14),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_4),
.B1(n_6),
.B2(n_91),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_73),
.A2(n_4),
.B1(n_79),
.B2(n_88),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_70),
.A2(n_80),
.B1(n_48),
.B2(n_76),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_85),
.A2(n_65),
.B1(n_63),
.B2(n_66),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_156),
.B1(n_152),
.B2(n_101),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_131),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_61),
.A2(n_89),
.B1(n_47),
.B2(n_82),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_126),
.B1(n_102),
.B2(n_156),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_54),
.A2(n_95),
.B1(n_50),
.B2(n_57),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_54),
.B(n_75),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_120),
.B(n_92),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_51),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_161),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_98),
.B(n_99),
.C(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_159),
.B(n_170),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_98),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_99),
.B1(n_148),
.B2(n_146),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_164),
.A2(n_174),
.B1(n_196),
.B2(n_106),
.Y(n_224)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_103),
.B(n_127),
.C(n_121),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_178),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_125),
.B(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_173),
.B(n_183),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_128),
.B1(n_115),
.B2(n_112),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_112),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_136),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_100),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_184),
.B(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_185),
.B(n_191),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_116),
.B(n_126),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_110),
.Y(n_227)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_130),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_110),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_152),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_190),
.B(n_175),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_101),
.B(n_114),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_198),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_114),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_109),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_200),
.Y(n_226)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_109),
.B(n_140),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_201),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_144),
.C(n_140),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_229),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_212),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_167),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_230),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_224),
.A2(n_195),
.B1(n_182),
.B2(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_200),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_168),
.C(n_159),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_190),
.A2(n_175),
.B(n_195),
.C(n_161),
.Y(n_231)
);

AO21x1_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_181),
.B(n_187),
.Y(n_255)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_168),
.A2(n_164),
.A3(n_170),
.B1(n_165),
.B2(n_172),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_186),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_165),
.B1(n_163),
.B2(n_158),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_234),
.A2(n_243),
.B1(n_225),
.B2(n_219),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_208),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_251),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_183),
.B(n_168),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_252),
.B(n_256),
.Y(n_259)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_160),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_258),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_202),
.A2(n_196),
.B1(n_179),
.B2(n_195),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_224),
.B1(n_213),
.B2(n_202),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_198),
.B1(n_176),
.B2(n_180),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_255),
.B1(n_223),
.B2(n_231),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_246),
.Y(n_270)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

BUFx8_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_162),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_257),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_209),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_192),
.B(n_181),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_181),
.C(n_169),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_235),
.C(n_252),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_193),
.B(n_166),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_177),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_217),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_251),
.B(n_210),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_266),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_210),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_269),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_215),
.B1(n_233),
.B2(n_212),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_280),
.B1(n_245),
.B2(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_219),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_260),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_215),
.C(n_205),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_276),
.C(n_226),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_221),
.C(n_213),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_223),
.B(n_209),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_281),
.B(n_249),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_242),
.B(n_223),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_234),
.B1(n_280),
.B2(n_265),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_287),
.B1(n_289),
.B2(n_294),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_285),
.A2(n_262),
.B(n_279),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_293),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_243),
.B1(n_255),
.B2(n_258),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_264),
.B(n_254),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_290),
.B(n_217),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_291),
.Y(n_317)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_261),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_255),
.A3(n_257),
.B1(n_226),
.B2(n_239),
.C1(n_247),
.C2(n_253),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_268),
.A2(n_259),
.B1(n_273),
.B2(n_271),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_302),
.C(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_238),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_300),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_236),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_269),
.A2(n_214),
.B1(n_207),
.B2(n_216),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_267),
.B1(n_277),
.B2(n_274),
.Y(n_311)
);

INVxp33_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

BUFx12f_ASAP7_75t_SL g301 ( 
.A(n_278),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_287),
.A2(n_259),
.B1(n_281),
.B2(n_264),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_307),
.C(n_309),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_275),
.C(n_276),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_290),
.B(n_263),
.CI(n_277),
.CON(n_308),
.SN(n_308)
);

XOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_308),
.B(n_291),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_267),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_311),
.A2(n_292),
.B1(n_286),
.B2(n_297),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_274),
.C(n_216),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_313),
.B(n_284),
.C(n_299),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_282),
.A2(n_262),
.B1(n_279),
.B2(n_248),
.Y(n_314)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_301),
.B(n_291),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_319),
.B(n_284),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_227),
.Y(n_320)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_320),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_294),
.A2(n_248),
.B1(n_207),
.B2(n_227),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_304),
.B(n_282),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_323),
.B(n_328),
.Y(n_350)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_288),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_322),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_336),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_313),
.B(n_321),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_334),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_306),
.B(n_284),
.C(n_203),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_335),
.B(n_317),
.Y(n_341)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_309),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_307),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_305),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_315),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_341),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

INVxp33_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_345),
.B(n_346),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_326),
.A2(n_310),
.B(n_317),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_334),
.A2(n_318),
.B(n_315),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_348),
.B(n_327),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_349),
.A2(n_325),
.B(n_332),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g366 ( 
.A1(n_352),
.A2(n_319),
.B(n_349),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_353),
.A2(n_346),
.B(n_340),
.Y(n_361)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_350),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_356),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_344),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_327),
.C(n_335),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_358),
.B(n_359),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_338),
.C(n_333),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_342),
.B(n_324),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_360),
.B(n_339),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_364),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_331),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_365),
.B(n_355),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_366),
.A2(n_367),
.B(n_308),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_357),
.A2(n_311),
.B(n_320),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_308),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_368),
.B(n_204),
.C(n_203),
.Y(n_375)
);

OAI21xp33_ASAP7_75t_L g377 ( 
.A1(n_371),
.A2(n_373),
.B(n_375),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_207),
.Y(n_372)
);

NOR2x1_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_232),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_363),
.A2(n_248),
.B(n_204),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_361),
.C(n_368),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_380),
.B(n_189),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_188),
.Y(n_382)
);

O2A1O1Ixp33_ASAP7_75t_SL g380 ( 
.A1(n_370),
.A2(n_228),
.B(n_188),
.C(n_232),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_370),
.C(n_232),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_382),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_377),
.B(n_228),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_188),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_386),
.B(n_385),
.Y(n_387)
);


endmodule