module fake_netlist_1_10177_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_4), .B(n_2), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_3), .B(n_2), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_11), .B(n_0), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_11), .B(n_0), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_10), .B(n_1), .Y(n_18) );
INVxp67_ASAP7_75t_SL g19 ( .A(n_14), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_19), .B(n_18), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_22), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AO21x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_16), .B(n_13), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_24), .B(n_21), .Y(n_27) );
AOI21xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_17), .B(n_18), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_25), .B(n_17), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_30), .B(n_15), .Y(n_32) );
NOR2xp33_ASAP7_75t_L g33 ( .A(n_28), .B(n_13), .Y(n_33) );
AOI22xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_12), .B1(n_3), .B2(n_1), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_31), .Y(n_35) );
AND3x4_ASAP7_75t_L g36 ( .A(n_34), .B(n_33), .C(n_5), .Y(n_36) );
NAND2xp5_ASAP7_75t_L g37 ( .A(n_36), .B(n_35), .Y(n_37) );
endmodule