module fake_jpeg_5887_n_251 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_251);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_28),
.Y(n_35)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_23),
.B(n_22),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_45),
.B(n_31),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_14),
.B1(n_21),
.B2(n_17),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_21),
.B1(n_25),
.B2(n_19),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_14),
.B1(n_17),
.B2(n_23),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_43),
.B1(n_21),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_14),
.B1(n_17),
.B2(n_22),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_34),
.B(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_62),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_23),
.B1(n_31),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_18),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_29),
.B1(n_34),
.B2(n_23),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_42),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_53),
.A2(n_36),
.B1(n_45),
.B2(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_40),
.B1(n_46),
.B2(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_75),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_38),
.B(n_46),
.C(n_18),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_62),
.Y(n_82)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_46),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_46),
.B1(n_40),
.B2(n_26),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_13),
.C(n_19),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_60),
.A3(n_58),
.B1(n_51),
.B2(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_86),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_84),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_70),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_91),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_40),
.B(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_99),
.B1(n_73),
.B2(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_95),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_42),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_67),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_19),
.B(n_47),
.Y(n_99)
);

NOR2xp67_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_81),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_104),
.B(n_94),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_89),
.B1(n_95),
.B2(n_97),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_79),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_94),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_67),
.C(n_65),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_114),
.C(n_82),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_76),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_64),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_117),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_18),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_99),
.B(n_93),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_126),
.Y(n_152)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_128),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_101),
.B1(n_26),
.B2(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_99),
.B(n_89),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_137),
.C(n_101),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_134),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_66),
.B1(n_16),
.B2(n_20),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_86),
.Y(n_136)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_91),
.C(n_92),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_104),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_146),
.C(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_115),
.B1(n_114),
.B2(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_140),
.A2(n_148),
.B1(n_123),
.B2(n_137),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_134),
.B1(n_136),
.B2(n_121),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_76),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_131),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_22),
.B1(n_66),
.B2(n_75),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_121),
.Y(n_162)
);

INVx13_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_32),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_153),
.A2(n_128),
.B(n_132),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_42),
.B1(n_44),
.B2(n_24),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_32),
.C(n_30),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_168),
.CI(n_152),
.CON(n_180),
.SN(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_163),
.B(n_169),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_124),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_120),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_153),
.A2(n_132),
.B(n_135),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_30),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_44),
.B1(n_16),
.B2(n_42),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_142),
.B1(n_149),
.B2(n_156),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_32),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_176),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_30),
.C(n_16),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_24),
.C(n_20),
.Y(n_187)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_152),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_184),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_180),
.B(n_172),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_147),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_164),
.B(n_140),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_151),
.B(n_154),
.C(n_16),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_174),
.C(n_171),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_24),
.B1(n_20),
.B2(n_2),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_24),
.B1(n_20),
.B2(n_2),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_192),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_195),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_203),
.C(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_205),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_170),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_159),
.C(n_161),
.Y(n_205)
);

AO221x1_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_167),
.B1(n_169),
.B2(n_162),
.C(n_3),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_212),
.B(n_216),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_208),
.A2(n_193),
.B(n_180),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_200),
.A2(n_191),
.B1(n_186),
.B2(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_198),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_215),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_187),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_197),
.B(n_186),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_6),
.B(n_11),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_208),
.B1(n_186),
.B2(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_7),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_224),
.B(n_6),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_6),
.B1(n_11),
.B2(n_10),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_9),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_12),
.C(n_4),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_4),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_213),
.B1(n_217),
.B2(n_8),
.Y(n_232)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_227),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_235),
.B(n_228),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_238),
.B(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_12),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_221),
.B(n_226),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_242),
.B(n_243),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_244),
.B(n_8),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_8),
.C(n_9),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_3),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_0),
.B(n_1),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_1),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_247),
.Y(n_251)
);


endmodule