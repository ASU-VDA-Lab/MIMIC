module fake_ariane_1388_n_1084 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1084);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1084;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_528;
wire n_584;
wire n_424;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_945;
wire n_702;
wire n_958;
wire n_905;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_989;
wire n_242;
wire n_645;
wire n_858;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_600;
wire n_481;
wire n_721;
wire n_840;
wire n_1053;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_617;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_583;
wire n_509;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_931;
wire n_827;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_976;
wire n_909;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_SL g199 ( 
.A(n_152),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_50),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_97),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_0),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_121),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_20),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_14),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_183),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_70),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_14),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_164),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_82),
.Y(n_219)
);

BUFx10_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_23),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_125),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_167),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_42),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_33),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_68),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_61),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_51),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_99),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_177),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_171),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_92),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_16),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_31),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_191),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_48),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_163),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_43),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_63),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g247 ( 
.A(n_157),
.B(n_60),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_69),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_169),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_129),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_62),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_90),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_85),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_182),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_16),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_84),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_57),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_24),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_3),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_78),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_66),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_103),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_179),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_9),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_156),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_176),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_30),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_139),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_220),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

BUFx2_ASAP7_75t_SL g280 ( 
.A(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_200),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_210),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_223),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_205),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_227),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_229),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_222),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_236),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_251),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_232),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_212),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_245),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_226),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_260),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_238),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_202),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_199),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_231),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_250),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_278),
.A2(n_247),
.B1(n_271),
.B2(n_270),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_304),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_250),
.Y(n_328)
);

NAND2xp33_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_250),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_280),
.B(n_259),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_314),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_204),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_314),
.Y(n_333)
);

BUFx8_ASAP7_75t_L g334 ( 
.A(n_318),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_259),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_283),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

OAI22x1_ASAP7_75t_SL g338 ( 
.A1(n_317),
.A2(n_320),
.B1(n_276),
.B2(n_274),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_316),
.A2(n_208),
.B(n_207),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_259),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_L g341 ( 
.A1(n_276),
.A2(n_272),
.B1(n_267),
.B2(n_213),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_313),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_214),
.Y(n_344)
);

OA21x2_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_217),
.B(n_216),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_288),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_259),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_277),
.B(n_218),
.Y(n_350)
);

OA21x2_ASAP7_75t_L g351 ( 
.A1(n_292),
.A2(n_224),
.B(n_219),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_293),
.B(n_225),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_275),
.A2(n_256),
.B1(n_255),
.B2(n_254),
.Y(n_354)
);

NOR2x1_ASAP7_75t_L g355 ( 
.A(n_279),
.B(n_230),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_282),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_282),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_233),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_303),
.Y(n_369)
);

BUFx8_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_306),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_273),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_307),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_309),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_358),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_310),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_341),
.B(n_295),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_327),
.B(n_343),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_312),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_361),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_344),
.B(n_315),
.Y(n_391)
);

INVx8_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_322),
.Y(n_393)
);

BUFx10_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_322),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_337),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_376),
.B(n_234),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_337),
.Y(n_402)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_336),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_336),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_317),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

AND3x2_ASAP7_75t_L g407 ( 
.A(n_325),
.B(n_0),
.C(n_1),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_342),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_342),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_239),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_350),
.B(n_240),
.Y(n_412)
);

AO21x2_ASAP7_75t_L g413 ( 
.A1(n_332),
.A2(n_244),
.B(n_243),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_375),
.B(n_355),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_343),
.B(n_248),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

INVxp33_ASAP7_75t_SL g419 ( 
.A(n_326),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_357),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_356),
.Y(n_421)
);

AO21x2_ASAP7_75t_L g422 ( 
.A1(n_354),
.A2(n_348),
.B(n_340),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_324),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_347),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_347),
.Y(n_426)
);

BUFx10_ASAP7_75t_L g427 ( 
.A(n_324),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_353),
.A2(n_253),
.B1(n_249),
.B2(n_3),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_347),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_353),
.B(n_1),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_347),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_373),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_363),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_363),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_340),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_2),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_346),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_324),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_349),
.B(n_2),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_324),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_L g447 ( 
.A(n_355),
.B(n_4),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_349),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_335),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_L g450 ( 
.A(n_364),
.B(n_4),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_397),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_419),
.B(n_323),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_394),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_323),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_395),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

AND2x6_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_335),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_394),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_408),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_393),
.B(n_362),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

AOI21x1_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_345),
.B(n_339),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_403),
.B(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_436),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_378),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_381),
.B(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_379),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_405),
.B(n_372),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

XNOR2x2_ASAP7_75t_L g475 ( 
.A(n_428),
.B(n_333),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_394),
.B(n_403),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_404),
.B(n_352),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_391),
.B(n_333),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_414),
.B(n_348),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_392),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_404),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_377),
.B(n_374),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_365),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_384),
.B(n_338),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_417),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_380),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_392),
.B(n_365),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_386),
.B(n_352),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_388),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_435),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_434),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_366),
.Y(n_496)
);

NAND2x1p5_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_444),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_445),
.B(n_366),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_439),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_444),
.B(n_367),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_434),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_437),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_431),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_439),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_441),
.B(n_338),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_401),
.B(n_334),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_367),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_423),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_392),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_392),
.B(n_334),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_437),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_334),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_442),
.B(n_368),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_411),
.B(n_329),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_442),
.B(n_368),
.Y(n_518)
);

AO21x1_ASAP7_75t_L g519 ( 
.A1(n_450),
.A2(n_335),
.B(n_351),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_443),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_423),
.B(n_335),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_400),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_443),
.Y(n_523)
);

CKINVDCx11_ASAP7_75t_R g524 ( 
.A(n_427),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_398),
.B(n_370),
.Y(n_525)
);

INVx4_ASAP7_75t_SL g526 ( 
.A(n_446),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_400),
.Y(n_527)
);

INVx4_ASAP7_75t_SL g528 ( 
.A(n_446),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_413),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_402),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_478),
.A2(n_450),
.B1(n_412),
.B2(n_447),
.Y(n_535)
);

AND2x6_ASAP7_75t_SL g536 ( 
.A(n_477),
.B(n_370),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_422),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_482),
.B(n_383),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_479),
.B(n_498),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_422),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_422),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_488),
.B(n_427),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_482),
.B(n_383),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_504),
.B(n_413),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_500),
.B(n_413),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_529),
.A2(n_351),
.B1(n_339),
.B2(n_345),
.Y(n_546)
);

NOR3xp33_ASAP7_75t_L g547 ( 
.A(n_453),
.B(n_447),
.C(n_421),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_500),
.B(n_383),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_455),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_455),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_473),
.B(n_370),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_503),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_475),
.A2(n_351),
.B1(n_339),
.B2(n_345),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_514),
.B(n_421),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_457),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_534),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_515),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_476),
.B(n_534),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_517),
.A2(n_425),
.B(n_421),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_451),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_518),
.B(n_425),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_484),
.B(n_425),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_534),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_532),
.A2(n_351),
.B1(n_339),
.B2(n_345),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_516),
.A2(n_410),
.B1(n_409),
.B2(n_415),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_513),
.B(n_382),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_533),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_491),
.B(n_382),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_514),
.B(n_410),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_513),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_458),
.B(n_415),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_461),
.B(n_416),
.Y(n_574)
);

INVxp67_ASAP7_75t_SL g575 ( 
.A(n_512),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_469),
.B(n_390),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_462),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_466),
.A2(n_485),
.B1(n_521),
.B2(n_459),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_494),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_494),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_502),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_477),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_467),
.Y(n_584)
);

INVx8_ASAP7_75t_L g585 ( 
.A(n_459),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_502),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_466),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_485),
.B(n_416),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_483),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_452),
.B(n_418),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_460),
.B(n_390),
.Y(n_591)
);

NOR2x1p5_ASAP7_75t_L g592 ( 
.A(n_487),
.B(n_407),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_459),
.B(n_396),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_508),
.B(n_418),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_456),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_459),
.A2(n_396),
.B1(n_399),
.B2(n_420),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_521),
.B(n_420),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_507),
.B(n_399),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_499),
.B(n_402),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_454),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_524),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_579),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_580),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_537),
.B(n_505),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_539),
.B(n_509),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_581),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_586),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_539),
.B(n_511),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_577),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_560),
.A2(n_496),
.B(n_490),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_551),
.B(n_486),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_563),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_585),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_556),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_569),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_600),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_520),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_590),
.A2(n_506),
.B1(n_544),
.B2(n_587),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_549),
.B(n_523),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_570),
.B(n_535),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_576),
.B(n_497),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_585),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_584),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_550),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_552),
.B(n_510),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_554),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_585),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_545),
.B(n_519),
.Y(n_629)
);

OR2x2_ASAP7_75t_SL g630 ( 
.A(n_536),
.B(n_525),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_540),
.B(n_468),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_540),
.B(n_470),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_568),
.B(n_526),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_568),
.B(n_526),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_557),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_599),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_599),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_594),
.B(n_471),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_557),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_561),
.B(n_472),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_568),
.B(n_474),
.Y(n_641)
);

NOR3xp33_ASAP7_75t_SL g642 ( 
.A(n_601),
.B(n_481),
.C(n_480),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_557),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_541),
.B(n_489),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_565),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_571),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_598),
.A2(n_495),
.B1(n_501),
.B2(n_492),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_573),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_565),
.B(n_493),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_573),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_589),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_571),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_572),
.B(n_528),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_595),
.B(n_542),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_574),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_541),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_564),
.B(n_528),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_565),
.B(n_522),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_527),
.Y(n_660)
);

BUFx8_ASAP7_75t_SL g661 ( 
.A(n_583),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_621),
.A2(n_555),
.B(n_593),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_610),
.A2(n_465),
.B(n_567),
.Y(n_663)
);

OAI21x1_ASAP7_75t_L g664 ( 
.A1(n_629),
.A2(n_567),
.B(n_555),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_631),
.A2(n_548),
.B(n_543),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_605),
.B(n_547),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_661),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_644),
.A2(n_538),
.B(n_591),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_629),
.A2(n_546),
.B(n_566),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_611),
.B(n_559),
.C(n_575),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_656),
.A2(n_538),
.B(n_588),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_623),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_622),
.A2(n_553),
.B(n_596),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_623),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_614),
.B(n_558),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_608),
.A2(n_597),
.B(n_592),
.C(n_531),
.Y(n_676)
);

INVx3_ASAP7_75t_SL g677 ( 
.A(n_630),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_SL g678 ( 
.A1(n_632),
.A2(n_389),
.B(n_424),
.Y(n_678)
);

AO31x2_ASAP7_75t_L g679 ( 
.A1(n_657),
.A2(n_432),
.A3(n_430),
.B(n_429),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_656),
.A2(n_426),
.B(n_424),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_640),
.B(n_426),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_646),
.A2(n_430),
.B(n_429),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_658),
.A2(n_432),
.B(n_389),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_646),
.A2(n_389),
.B(n_26),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_626),
.A2(n_389),
.B(n_27),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_633),
.B(n_389),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_652),
.A2(n_28),
.B(n_25),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_635),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_638),
.A2(n_650),
.B(n_648),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_655),
.A2(n_32),
.B(n_29),
.Y(n_690)
);

OAI21xp33_ASAP7_75t_SL g691 ( 
.A1(n_638),
.A2(n_5),
.B(n_6),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_604),
.B(n_6),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_632),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_604),
.B(n_7),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_652),
.A2(n_35),
.B(n_34),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_627),
.B(n_8),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_660),
.A2(n_10),
.B(n_11),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_627),
.B(n_10),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_635),
.B(n_11),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_623),
.Y(n_700)
);

AO21x2_ASAP7_75t_L g701 ( 
.A1(n_636),
.A2(n_37),
.B(n_36),
.Y(n_701)
);

CKINVDCx6p67_ASAP7_75t_R g702 ( 
.A(n_639),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_636),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_637),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_602),
.Y(n_705)
);

AO31x2_ASAP7_75t_L g706 ( 
.A1(n_637),
.A2(n_119),
.A3(n_196),
.B(n_195),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_628),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_628),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_649),
.A2(n_117),
.B(n_194),
.Y(n_709)
);

NOR2x1_ASAP7_75t_L g710 ( 
.A(n_639),
.B(n_39),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_619),
.B(n_12),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_649),
.A2(n_118),
.B(n_193),
.Y(n_712)
);

AO31x2_ASAP7_75t_L g713 ( 
.A1(n_603),
.A2(n_116),
.A3(n_192),
.B(n_189),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_620),
.A2(n_625),
.B(n_641),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_651),
.B(n_12),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_635),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_603),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_702),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_711),
.A2(n_654),
.B1(n_641),
.B2(n_634),
.Y(n_719)
);

BUFx5_ASAP7_75t_L g720 ( 
.A(n_703),
.Y(n_720)
);

NOR2x1_ASAP7_75t_SL g721 ( 
.A(n_666),
.B(n_641),
.Y(n_721)
);

OAI21x1_ASAP7_75t_L g722 ( 
.A1(n_663),
.A2(n_649),
.B(n_607),
.Y(n_722)
);

AO32x2_ASAP7_75t_L g723 ( 
.A1(n_693),
.A2(n_643),
.A3(n_679),
.B1(n_714),
.B2(n_691),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_675),
.B(n_661),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_668),
.A2(n_662),
.B(n_678),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_697),
.A2(n_642),
.B(n_618),
.C(n_624),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_689),
.A2(n_676),
.B(n_692),
.C(n_694),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_703),
.B(n_609),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_SL g729 ( 
.A1(n_699),
.A2(n_696),
.B(n_698),
.C(n_707),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_715),
.B(n_617),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_717),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_677),
.B(n_620),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_667),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_670),
.A2(n_641),
.B1(n_633),
.B2(n_634),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_685),
.A2(n_660),
.B(n_618),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_SL g736 ( 
.A(n_686),
.B(n_633),
.Y(n_736)
);

OAI21x1_ASAP7_75t_L g737 ( 
.A1(n_683),
.A2(n_607),
.B(n_606),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_665),
.A2(n_612),
.B(n_606),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_681),
.B(n_672),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_688),
.Y(n_740)
);

AO31x2_ASAP7_75t_L g741 ( 
.A1(n_704),
.A2(n_612),
.A3(n_615),
.B(n_616),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_717),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_704),
.B(n_615),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_673),
.A2(n_690),
.B(n_671),
.C(n_664),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_688),
.Y(n_745)
);

AOI221x1_ASAP7_75t_L g746 ( 
.A1(n_680),
.A2(n_616),
.B1(n_634),
.B2(n_659),
.C(n_645),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_672),
.A2(n_635),
.B(n_645),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_674),
.B(n_643),
.C(n_653),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_686),
.B(n_613),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_684),
.A2(n_628),
.B(n_647),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_705),
.B(n_653),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_679),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_679),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_674),
.A2(n_645),
.B(n_635),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_688),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_716),
.B(n_653),
.Y(n_756)
);

AO21x1_ASAP7_75t_L g757 ( 
.A1(n_687),
.A2(n_659),
.B(n_645),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_700),
.A2(n_613),
.B1(n_630),
.B2(n_645),
.Y(n_758)
);

NAND2x1_ASAP7_75t_L g759 ( 
.A(n_700),
.B(n_659),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_707),
.A2(n_13),
.B(n_15),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_R g761 ( 
.A(n_716),
.B(n_40),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_716),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_669),
.A2(n_13),
.B(n_15),
.C(n_17),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_710),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_701),
.A2(n_123),
.A3(n_188),
.B(n_187),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_708),
.B(n_18),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_682),
.A2(n_122),
.B(n_186),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_708),
.A2(n_701),
.B(n_712),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_709),
.A2(n_19),
.B(n_20),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_695),
.A2(n_21),
.B(n_22),
.Y(n_770)
);

AO31x2_ASAP7_75t_L g771 ( 
.A1(n_706),
.A2(n_124),
.A3(n_185),
.B(n_184),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_706),
.A2(n_21),
.B(n_22),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_706),
.A2(n_23),
.B(n_198),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_SL g774 ( 
.A1(n_713),
.A2(n_41),
.B(n_44),
.C(n_45),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_713),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_SL g776 ( 
.A1(n_713),
.A2(n_46),
.B(n_47),
.C(n_49),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_675),
.B(n_52),
.Y(n_777)
);

OA21x2_ASAP7_75t_L g778 ( 
.A1(n_663),
.A2(n_53),
.B(n_54),
.Y(n_778)
);

AOI211xp5_ASAP7_75t_L g779 ( 
.A1(n_697),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_779)
);

OA21x2_ASAP7_75t_L g780 ( 
.A1(n_663),
.A2(n_59),
.B(n_64),
.Y(n_780)
);

AOI21x1_ASAP7_75t_L g781 ( 
.A1(n_683),
.A2(n_65),
.B(n_67),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_731),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_732),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_730),
.B(n_74),
.Y(n_784)
);

NOR2x1_ASAP7_75t_L g785 ( 
.A(n_755),
.B(n_75),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_719),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_734),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_733),
.Y(n_788)
);

BUFx12f_ASAP7_75t_L g789 ( 
.A(n_718),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_742),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_740),
.Y(n_792)
);

INVx6_ASAP7_75t_L g793 ( 
.A(n_745),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_770),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_794)
);

CKINVDCx6p67_ASAP7_75t_R g795 ( 
.A(n_749),
.Y(n_795)
);

CKINVDCx8_ASAP7_75t_R g796 ( 
.A(n_724),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_726),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_741),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_751),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_741),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_777),
.A2(n_101),
.B1(n_102),
.B2(n_104),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_728),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_762),
.Y(n_803)
);

INVx6_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_756),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_720),
.B(n_105),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_720),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_761),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_758),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_743),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_772),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_720),
.Y(n_812)
);

CKINVDCx11_ASAP7_75t_R g813 ( 
.A(n_752),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_SL g814 ( 
.A1(n_721),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_759),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_739),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_748),
.B(n_727),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_735),
.A2(n_114),
.B1(n_115),
.B2(n_126),
.Y(n_818)
);

CKINVDCx20_ASAP7_75t_R g819 ( 
.A(n_766),
.Y(n_819)
);

CKINVDCx11_ASAP7_75t_R g820 ( 
.A(n_753),
.Y(n_820)
);

BUFx2_ASAP7_75t_SL g821 ( 
.A(n_757),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_769),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_722),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_775),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_773),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_737),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_778),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_750),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_SL g829 ( 
.A1(n_779),
.A2(n_137),
.B1(n_138),
.B2(n_140),
.Y(n_829)
);

INVx6_ASAP7_75t_L g830 ( 
.A(n_736),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_764),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_723),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_746),
.Y(n_833)
);

BUFx8_ASAP7_75t_SL g834 ( 
.A(n_781),
.Y(n_834)
);

BUFx8_ASAP7_75t_SL g835 ( 
.A(n_767),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_763),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_798),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_782),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_804),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_790),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_789),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_800),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_791),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_810),
.Y(n_844)
);

BUFx3_ASAP7_75t_L g845 ( 
.A(n_792),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_804),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_826),
.A2(n_725),
.B(n_768),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_832),
.B(n_723),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_802),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_824),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_797),
.A2(n_817),
.B(n_836),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_812),
.Y(n_852)
);

OA21x2_ASAP7_75t_L g853 ( 
.A1(n_827),
.A2(n_744),
.B(n_738),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_828),
.Y(n_854)
);

OAI21x1_ASAP7_75t_L g855 ( 
.A1(n_806),
.A2(n_780),
.B(n_747),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_823),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_827),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_806),
.A2(n_754),
.B(n_760),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_821),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_816),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_833),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_815),
.A2(n_797),
.B(n_836),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_788),
.B(n_729),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_804),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_807),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_815),
.A2(n_776),
.B(n_774),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_816),
.Y(n_868)
);

AND2x4_ASAP7_75t_L g869 ( 
.A(n_803),
.B(n_771),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_813),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_805),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_820),
.Y(n_872)
);

OAI22xp33_ASAP7_75t_L g873 ( 
.A1(n_831),
.A2(n_771),
.B1(n_765),
.B2(n_150),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_835),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_834),
.Y(n_875)
);

INVx4_ASAP7_75t_SL g876 ( 
.A(n_830),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_809),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_838),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_838),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_839),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_860),
.Y(n_881)
);

BUFx12f_ASAP7_75t_L g882 ( 
.A(n_841),
.Y(n_882)
);

AO21x2_ASAP7_75t_L g883 ( 
.A1(n_861),
.A2(n_787),
.B(n_784),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_843),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_843),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_837),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_868),
.B(n_795),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_844),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_848),
.B(n_819),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_861),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_850),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_845),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_844),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_848),
.B(n_790),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_850),
.B(n_790),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_857),
.B(n_808),
.Y(n_896)
);

AO21x2_ASAP7_75t_L g897 ( 
.A1(n_851),
.A2(n_765),
.B(n_825),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_857),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_839),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_845),
.B(n_856),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_842),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_856),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_871),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_842),
.Y(n_904)
);

OA21x2_ASAP7_75t_L g905 ( 
.A1(n_847),
.A2(n_818),
.B(n_794),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_890),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_891),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_886),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_886),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_878),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_881),
.B(n_859),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_889),
.B(n_870),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_878),
.Y(n_913)
);

AOI21xp33_ASAP7_75t_L g914 ( 
.A1(n_897),
.A2(n_859),
.B(n_863),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_886),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_880),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_879),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_879),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_889),
.B(n_870),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_882),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_884),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_903),
.B(n_877),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_884),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_885),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_900),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_902),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_900),
.B(n_872),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_908),
.Y(n_928)
);

OR2x2_ASAP7_75t_SL g929 ( 
.A(n_920),
.B(n_872),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_912),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_925),
.B(n_892),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_925),
.B(n_892),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_906),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_916),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_916),
.B(n_897),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_926),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_910),
.Y(n_937)
);

AND3x1_ASAP7_75t_L g938 ( 
.A(n_912),
.B(n_874),
.C(n_875),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_916),
.B(n_897),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_927),
.B(n_903),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_920),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_911),
.Y(n_942)
);

AOI221xp5_ASAP7_75t_L g943 ( 
.A1(n_914),
.A2(n_873),
.B1(n_874),
.B2(n_875),
.C(n_898),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_938),
.B(n_927),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_938),
.B(n_919),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_937),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_930),
.B(n_933),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_930),
.B(n_919),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_940),
.B(n_922),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_942),
.B(n_913),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_941),
.B(n_920),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_940),
.B(n_922),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_931),
.B(n_907),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_931),
.B(n_920),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_946),
.B(n_933),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_947),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_945),
.B(n_941),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_949),
.B(n_936),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_948),
.B(n_950),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_951),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_951),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_954),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_960),
.B(n_955),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_961),
.B(n_948),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_963),
.B(n_948),
.Y(n_966)
);

OAI22xp33_ASAP7_75t_L g967 ( 
.A1(n_959),
.A2(n_943),
.B1(n_944),
.B2(n_952),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_958),
.B(n_941),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_956),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_969),
.B(n_950),
.Y(n_970)
);

NOR4xp25_ASAP7_75t_SL g971 ( 
.A(n_964),
.B(n_962),
.C(n_957),
.D(n_841),
.Y(n_971)
);

OAI21xp33_ASAP7_75t_SL g972 ( 
.A1(n_968),
.A2(n_956),
.B(n_952),
.Y(n_972)
);

NAND2x1p5_ASAP7_75t_L g973 ( 
.A(n_965),
.B(n_887),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_966),
.B(n_953),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_967),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_965),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_969),
.B(n_935),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_967),
.A2(n_929),
.B1(n_952),
.B2(n_935),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_965),
.Y(n_979)
);

OAI22xp33_ASAP7_75t_L g980 ( 
.A1(n_978),
.A2(n_929),
.B1(n_935),
.B2(n_939),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_971),
.A2(n_939),
.B1(n_935),
.B2(n_911),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_979),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_970),
.B(n_882),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_972),
.Y(n_984)
);

AOI221xp5_ASAP7_75t_L g985 ( 
.A1(n_975),
.A2(n_939),
.B1(n_883),
.B2(n_869),
.C(n_928),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_979),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_976),
.B(n_939),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_982),
.A2(n_974),
.B(n_973),
.Y(n_988)
);

NAND3xp33_ASAP7_75t_L g989 ( 
.A(n_986),
.B(n_977),
.C(n_825),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_987),
.Y(n_990)
);

AOI222xp33_ASAP7_75t_L g991 ( 
.A1(n_985),
.A2(n_829),
.B1(n_928),
.B2(n_898),
.C1(n_869),
.C2(n_822),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_983),
.B(n_932),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_984),
.B(n_932),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_980),
.A2(n_883),
.B1(n_887),
.B2(n_896),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_981),
.B(n_934),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_990),
.Y(n_996)
);

OAI222xp33_ASAP7_75t_L g997 ( 
.A1(n_994),
.A2(n_896),
.B1(n_796),
.B2(n_894),
.C1(n_785),
.C2(n_895),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_993),
.A2(n_934),
.B(n_883),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_988),
.B(n_934),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_992),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_989),
.A2(n_995),
.B(n_991),
.C(n_862),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_1000),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_996),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_999),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_997),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1001),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_998),
.Y(n_1007)
);

INVxp33_ASAP7_75t_SL g1008 ( 
.A(n_1000),
.Y(n_1008)
);

NOR2x1_ASAP7_75t_L g1009 ( 
.A(n_996),
.B(n_895),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_L g1010 ( 
.A(n_1002),
.B(n_917),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_1003),
.B(n_814),
.C(n_894),
.Y(n_1011)
);

NOR3x1_ASAP7_75t_L g1012 ( 
.A(n_1004),
.B(n_862),
.C(n_923),
.Y(n_1012)
);

AND4x1_ASAP7_75t_L g1013 ( 
.A(n_1008),
.B(n_783),
.C(n_801),
.D(n_786),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1008),
.B(n_918),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_L g1015 ( 
.A(n_1006),
.B(n_811),
.C(n_799),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_1009),
.B(n_880),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1005),
.B(n_921),
.Y(n_1017)
);

NAND5xp2_ASAP7_75t_SL g1018 ( 
.A(n_1017),
.B(n_1007),
.C(n_793),
.D(n_840),
.E(n_899),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1014),
.Y(n_1019)
);

NOR2xp67_ASAP7_75t_L g1020 ( 
.A(n_1016),
.B(n_924),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_1015),
.A2(n_869),
.B1(n_905),
.B2(n_854),
.Y(n_1021)
);

NOR2x1_ASAP7_75t_L g1022 ( 
.A(n_1010),
.B(n_880),
.Y(n_1022)
);

NOR5xp2_ASAP7_75t_L g1023 ( 
.A(n_1019),
.B(n_1012),
.C(n_1011),
.D(n_1013),
.E(n_888),
.Y(n_1023)
);

NOR2x1p5_ASAP7_75t_L g1024 ( 
.A(n_1018),
.B(n_880),
.Y(n_1024)
);

AOI221xp5_ASAP7_75t_L g1025 ( 
.A1(n_1021),
.A2(n_888),
.B1(n_893),
.B2(n_885),
.C(n_852),
.Y(n_1025)
);

AOI221xp5_ASAP7_75t_SL g1026 ( 
.A1(n_1020),
.A2(n_852),
.B1(n_865),
.B2(n_867),
.C(n_893),
.Y(n_1026)
);

OAI211xp5_ASAP7_75t_L g1027 ( 
.A1(n_1022),
.A2(n_899),
.B(n_867),
.C(n_865),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_1019),
.B(n_899),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_1019),
.B(n_905),
.C(n_864),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_1019),
.Y(n_1030)
);

NOR2x1_ASAP7_75t_L g1031 ( 
.A(n_1019),
.B(n_899),
.Y(n_1031)
);

NAND3xp33_ASAP7_75t_L g1032 ( 
.A(n_1030),
.B(n_1023),
.C(n_1028),
.Y(n_1032)
);

AOI211xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_869),
.B(n_866),
.C(n_855),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_1024),
.Y(n_1034)
);

NOR2x1_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_839),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_1029),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1025),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1026),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_R g1039 ( 
.A(n_1030),
.B(n_793),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1030),
.B(n_915),
.Y(n_1040)
);

NAND3x1_ASAP7_75t_L g1041 ( 
.A(n_1028),
.B(n_846),
.C(n_864),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_1032),
.B(n_148),
.C(n_149),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1040),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_1039),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_1034),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1041),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_1038),
.B(n_846),
.Y(n_1047)
);

NOR2x1p5_ASAP7_75t_L g1048 ( 
.A(n_1037),
.B(n_846),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_SL g1049 ( 
.A1(n_1036),
.A2(n_905),
.B1(n_793),
.B2(n_908),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_1035),
.B(n_876),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_1033),
.B(n_866),
.C(n_153),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_L g1052 ( 
.A(n_1032),
.B(n_151),
.C(n_154),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1036),
.B(n_915),
.Y(n_1053)
);

NOR4xp25_ASAP7_75t_L g1054 ( 
.A(n_1032),
.B(n_909),
.C(n_854),
.D(n_849),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1045),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1042),
.B(n_909),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1043),
.Y(n_1057)
);

OR2x6_ASAP7_75t_L g1058 ( 
.A(n_1044),
.B(n_830),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_1050),
.Y(n_1059)
);

OAI22xp33_ASAP7_75t_SL g1060 ( 
.A1(n_1046),
.A2(n_830),
.B1(n_849),
.B2(n_901),
.Y(n_1060)
);

AOI211xp5_ASAP7_75t_L g1061 ( 
.A1(n_1052),
.A2(n_855),
.B(n_858),
.C(n_847),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1054),
.B(n_905),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_1053),
.B(n_1047),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1055),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1057),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_1059),
.A2(n_1048),
.B1(n_1051),
.B2(n_1049),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1056),
.Y(n_1067)
);

AO22x2_ASAP7_75t_L g1068 ( 
.A1(n_1062),
.A2(n_1063),
.B1(n_1058),
.B2(n_1060),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1061),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_1055),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1055),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_1070),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1064),
.A2(n_853),
.B1(n_904),
.B2(n_901),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1065),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1072),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1075),
.Y(n_1076)
);

XNOR2xp5_ASAP7_75t_L g1077 ( 
.A(n_1076),
.B(n_1071),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_1074),
.B1(n_1069),
.B2(n_1067),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_1077),
.A2(n_1066),
.B1(n_1068),
.B2(n_1073),
.Y(n_1079)
);

OA21x2_ASAP7_75t_L g1080 ( 
.A1(n_1079),
.A2(n_158),
.B(n_159),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1078),
.B(n_162),
.Y(n_1081)
);

AO21x2_ASAP7_75t_L g1082 ( 
.A1(n_1081),
.A2(n_1080),
.B(n_165),
.Y(n_1082)
);

A2O1A1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_1082),
.A2(n_168),
.B(n_170),
.C(n_172),
.Y(n_1083)
);

AOI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1083),
.A2(n_173),
.B(n_174),
.C(n_175),
.Y(n_1084)
);


endmodule