module real_jpeg_32296_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_1),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_3),
.B(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_3),
.B(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

AOI222xp33_ASAP7_75t_SL g36 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.C1(n_41),
.C2(n_45),
.Y(n_36)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_13),
.B1(n_29),
.B2(n_32),
.C(n_36),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_11),
.B(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_12),
.B(n_19),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_19),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_22),
.B(n_26),
.Y(n_13)
);

AO21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B(n_20),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_21),
.Y(n_20)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_23),
.Y(n_27)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);


endmodule