module real_jpeg_24761_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx6_ASAP7_75t_L g80 ( 
.A(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_83),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_5),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_6),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_57),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_7),
.A2(n_27),
.B1(n_61),
.B2(n_62),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_7),
.A2(n_27),
.B1(n_34),
.B2(n_35),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_7),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_9),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_11),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_99)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_15),
.B(n_61),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_15),
.B(n_69),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_15),
.B(n_35),
.C(n_37),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_71),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_15),
.B(n_40),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_15),
.A2(n_34),
.B1(n_35),
.B2(n_71),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_48),
.C(n_52),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_15),
.A2(n_79),
.B(n_166),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_101),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_91),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_21),
.A2(n_22),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_25),
.B(n_43),
.C(n_58),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_26),
.Y(n_93)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_30),
.B1(n_64),
.B2(n_65),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_28),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_28),
.B(n_131),
.Y(n_130)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g89 ( 
.A1(n_30),
.A2(n_62),
.A3(n_65),
.B1(n_73),
.B2(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_32),
.A2(n_106),
.B(n_107),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_32),
.A2(n_107),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_33),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_35),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_35),
.B(n_173),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_40),
.B(n_95),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_41),
.Y(n_106)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_53),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_45),
.A2(n_47),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_47),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_47),
.A2(n_53),
.B(n_138),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_47),
.B(n_71),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_49),
.B(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_54),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_56),
.B(n_140),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_70),
.B(n_74),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_68),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_71),
.B(n_192),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_76),
.B(n_91),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_89),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_89),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_84),
.B2(n_87),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_78),
.A2(n_177),
.B1(n_179),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_82),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_85),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_79),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_98),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_92),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_122),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_120),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_120),
.A2(n_154),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_205),
.B(n_210),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_155),
.B(n_204),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_144),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_128),
.B(n_144),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_136),
.C(n_141),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_129),
.B(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_136),
.A2(n_141),
.B1(n_142),
.B2(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_145),
.B(n_151),
.C(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_198),
.B(n_203),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_174),
.B(n_197),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_168),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_168),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_164),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_163),
.C(n_164),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_184),
.B(n_196),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_182),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_178),
.A2(n_180),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_189),
.B(n_195),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_187),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_202),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_209),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);


endmodule