module fake_jpeg_5144_n_250 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_28),
.B(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_16),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_20),
.B1(n_15),
.B2(n_32),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_32),
.B1(n_26),
.B2(n_20),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_26),
.B1(n_36),
.B2(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_34),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_41),
.B1(n_36),
.B2(n_25),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_33),
.C(n_25),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_23),
.B(n_40),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_72),
.C(n_77),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_41),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_52),
.B1(n_54),
.B2(n_51),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_40),
.C(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_38),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_14),
.B(n_19),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_62),
.C(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_57),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_72),
.B(n_12),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_95),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_37),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_96),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_67),
.A2(n_53),
.B1(n_35),
.B2(n_29),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_79),
.B1(n_78),
.B2(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_59),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

BUFx24_ASAP7_75t_SL g95 ( 
.A(n_61),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_48),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_69),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_107),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_66),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_112),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_79),
.B1(n_93),
.B2(n_83),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_104),
.B(n_61),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_130),
.C(n_131),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_110),
.Y(n_119)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_122),
.B1(n_124),
.B2(n_127),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_96),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_93),
.B1(n_81),
.B2(n_91),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_81),
.B1(n_92),
.B2(n_93),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_99),
.B(n_98),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_128),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_93),
.B1(n_91),
.B2(n_87),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_96),
.B(n_89),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_134),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_87),
.B(n_77),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_48),
.B(n_19),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_35),
.C(n_37),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_21),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_137),
.Y(n_172)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_109),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_133),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_110),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_106),
.B1(n_102),
.B2(n_108),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_130),
.B1(n_118),
.B2(n_128),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_102),
.B1(n_59),
.B2(n_45),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_64),
.B1(n_68),
.B2(n_36),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_149),
.B(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_131),
.B(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_64),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_152),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_125),
.C(n_115),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_161),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_164),
.B1(n_168),
.B2(n_13),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_153),
.C(n_142),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_37),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_174),
.B1(n_137),
.B2(n_155),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_37),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_170),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_41),
.B1(n_36),
.B2(n_35),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_169),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_36),
.B1(n_41),
.B2(n_13),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_151),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_39),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_45),
.B1(n_22),
.B2(n_21),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_191),
.C(n_39),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_149),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_177),
.A2(n_186),
.B(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_185),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_142),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_152),
.B1(n_155),
.B2(n_138),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_143),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_39),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_189),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_173),
.B(n_22),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_39),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_39),
.C(n_38),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_14),
.B1(n_35),
.B2(n_18),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_167),
.C(n_163),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_194),
.B(n_195),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_179),
.A2(n_157),
.B(n_164),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.C(n_205),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_187),
.A2(n_46),
.B(n_39),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_38),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_46),
.C(n_38),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_38),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_181),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_46),
.C(n_38),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_191),
.A2(n_46),
.B1(n_38),
.B2(n_17),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_38),
.B1(n_30),
.B2(n_29),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_208),
.A2(n_209),
.B(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_180),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_199),
.B(n_182),
.Y(n_213)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_216),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_30),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_0),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_1),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_211),
.A3(n_216),
.B1(n_202),
.B2(n_206),
.C1(n_30),
.C2(n_29),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_222),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_30),
.A3(n_29),
.B1(n_8),
.B2(n_9),
.C1(n_12),
.C2(n_6),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_224),
.B(n_225),
.C(n_228),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_0),
.C(n_1),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_3),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_3),
.C(n_4),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_9),
.B(n_12),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_231),
.A2(n_11),
.B(n_4),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_9),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_236),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_8),
.B(n_11),
.C(n_10),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_10),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_3),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_7),
.Y(n_236)
);

NAND2xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_227),
.Y(n_237)
);

NOR3xp33_ASAP7_75t_SL g243 ( 
.A(n_237),
.B(n_235),
.C(n_29),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_11),
.B(n_5),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_230),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_241),
.B(n_242),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_5),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_246),
.C(n_239),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_4),
.B(n_5),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_245),
.Y(n_250)
);


endmodule