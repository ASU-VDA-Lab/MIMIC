module fake_jpeg_29442_n_41 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_41);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_37;
wire n_32;

INVx11_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_9),
.B(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_3),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_20),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_23),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_23),
.B(n_18),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_32),
.B(n_33),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_21),
.B(n_17),
.Y(n_38)
);

OAI31xp33_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_1),
.A3(n_4),
.B(n_25),
.Y(n_39)
);

OAI311xp33_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_6),
.A3(n_13),
.B1(n_14),
.C1(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);


endmodule