module real_jpeg_7149_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g199 ( 
.A(n_0),
.Y(n_199)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_0),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_0),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_0),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B1(n_23),
.B2(n_26),
.Y(n_19)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_2),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_2),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_2),
.Y(n_330)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_2),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_2),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_3),
.A2(n_282),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_3),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_3),
.A2(n_284),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_3),
.A2(n_284),
.B1(n_289),
.B2(n_392),
.Y(n_391)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_3),
.A2(n_52),
.B1(n_284),
.B2(n_457),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_4),
.A2(n_213),
.B1(n_217),
.B2(n_218),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_4),
.A2(n_205),
.B1(n_217),
.B2(n_239),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_4),
.A2(n_91),
.B1(n_217),
.B2(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_4),
.A2(n_217),
.B1(n_329),
.B2(n_429),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_97),
.B1(n_98),
.B2(n_101),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_5),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_101),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_60),
.B1(n_101),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_5),
.A2(n_101),
.B1(n_382),
.B2(n_383),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_8),
.A2(n_133),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_8),
.A2(n_173),
.B1(n_205),
.B2(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_8),
.A2(n_173),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_8),
.A2(n_152),
.B1(n_173),
.B2(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_11),
.A2(n_164),
.B1(n_166),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_11),
.B(n_180),
.C(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_11),
.B(n_78),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_11),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_11),
.B(n_131),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_11),
.B(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_12),
.Y(n_186)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_88),
.B1(n_91),
.B2(n_94),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_14),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_94),
.B1(n_141),
.B2(n_146),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_14),
.A2(n_94),
.B1(n_182),
.B2(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_14),
.A2(n_94),
.B1(n_407),
.B2(n_411),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_15),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_15),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_15),
.A2(n_133),
.B1(n_192),
.B2(n_214),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_15),
.A2(n_192),
.B1(n_289),
.B2(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_15),
.A2(n_55),
.B1(n_62),
.B2(n_192),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_16),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_16),
.A2(n_56),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_16),
.A2(n_56),
.B1(n_213),
.B2(n_368),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_16),
.A2(n_56),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_18),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_18),
.A2(n_63),
.B1(n_342),
.B2(n_344),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_18),
.A2(n_63),
.B1(n_135),
.B2(n_388),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_18),
.A2(n_63),
.B1(n_392),
.B2(n_442),
.Y(n_441)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_534),
.B(n_537),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_153),
.B(n_533),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_150),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_29),
.B(n_150),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_139),
.C(n_147),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_30),
.A2(n_31),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_64),
.C(n_102),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_32),
.B(n_521),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_51),
.B1(n_57),
.B2(n_59),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_33),
.A2(n_57),
.B1(n_59),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_33),
.A2(n_57),
.B1(n_140),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_33),
.A2(n_354),
.B(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_33),
.A2(n_57),
.B1(n_402),
.B2(n_428),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_33),
.A2(n_51),
.B1(n_57),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_34),
.A2(n_351),
.B(n_353),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_34),
.B(n_355),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_34),
.A2(n_58),
.B(n_536),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_40),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_35)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_36),
.Y(n_332)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx8_ASAP7_75t_L g352 ( 
.A(n_37),
.Y(n_352)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_43),
.Y(n_334)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_46),
.Y(n_273)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_57),
.B(n_169),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_57),
.A2(n_428),
.B(n_460),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_58),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_58),
.B(n_456),
.Y(n_455)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_60),
.Y(n_146)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_64),
.A2(n_102),
.B1(n_103),
.B2(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_64),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_87),
.B1(n_95),
.B2(n_96),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_65),
.A2(n_95),
.B1(n_307),
.B2(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_65),
.A2(n_95),
.B1(n_391),
.B2(n_395),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_65),
.A2(n_87),
.B1(n_95),
.B2(n_510),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_78),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_69),
.B1(n_73),
.B2(n_76),
.Y(n_66)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_67),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_69),
.Y(n_276)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_72),
.Y(n_268)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_72),
.Y(n_328)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_72),
.Y(n_444)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_78)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_75),
.Y(n_294)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_77),
.Y(n_400)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_78),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

AOI22x1_ASAP7_75t_L g431 ( 
.A1(n_78),
.A2(n_148),
.B1(n_310),
.B2(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_78),
.A2(n_148),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_82),
.Y(n_410)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_88),
.B(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_90),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_90),
.Y(n_397)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_92),
.Y(n_277)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_95),
.B(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_95),
.A2(n_307),
.B(n_309),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_97),
.Y(n_289)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_102),
.A2(n_103),
.B1(n_508),
.B2(n_509),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_102),
.B(n_505),
.C(n_508),
.Y(n_516)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_130),
.B(n_132),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_163),
.B(n_170),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_104),
.A2(n_130),
.B1(n_212),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_104),
.A2(n_170),
.B(n_264),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_104),
.A2(n_130),
.B1(n_365),
.B2(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_105),
.B(n_171),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_105),
.A2(n_131),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_105),
.A2(n_131),
.B1(n_387),
.B2(n_406),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_105),
.A2(n_131),
.B1(n_406),
.B2(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_117),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_112),
.B2(n_115),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g368 ( 
.A(n_107),
.Y(n_368)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_108),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_116),
.Y(n_292)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_117),
.A2(n_212),
.B(n_221),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_123),
.Y(n_286)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_123),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_125),
.Y(n_241)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_130),
.A2(n_221),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_131),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_132),
.Y(n_447)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp33_ASAP7_75t_SL g295 ( 
.A(n_136),
.B(n_296),
.Y(n_295)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_138),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_138),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_138),
.Y(n_367)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_138),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_139),
.B(n_147),
.Y(n_530)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_142),
.B(n_169),
.Y(n_335)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_145),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_148),
.A2(n_267),
.B(n_274),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_148),
.B(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_148),
.A2(n_274),
.B(n_473),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_150),
.B(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_150),
.B(n_535),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_151),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_527),
.B(n_532),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_499),
.B(n_524),
.Y(n_154)
);

OAI311xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_371),
.A3(n_475),
.B1(n_493),
.C1(n_494),
.Y(n_155)
);

AOI21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_321),
.B(n_370),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_298),
.B(n_320),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_258),
.B(n_297),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_224),
.B(n_257),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_187),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_161),
.B(n_187),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_174),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_162),
.A2(n_174),
.B1(n_175),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_162),
.Y(n_255)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_169),
.A2(n_196),
.B(n_202),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_SL g267 ( 
.A1(n_169),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_SL g351 ( 
.A1(n_169),
.A2(n_335),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_184),
.Y(n_343)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_209),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_188),
.B(n_210),
.C(n_223),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_196),
.B(n_202),
.Y(n_188)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_195),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_196),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_196),
.A2(n_252),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_196),
.A2(n_381),
.B(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_204),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_197),
.A2(n_281),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_197),
.A2(n_317),
.B1(n_341),
.B2(n_425),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_199),
.Y(n_318)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_207),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_222),
.B2(n_223),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_247),
.B(n_256),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_236),
.B(n_246),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_235),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_233),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_232),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_245),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_245),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_242),
.B(n_244),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_244),
.A2(n_280),
.B(n_287),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_254),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_254),
.Y(n_256)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_260),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_278),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_265),
.B2(n_266),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_265),
.C(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_289),
.A3(n_290),
.B1(n_293),
.B2(n_295),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_288),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx5_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_299),
.B(n_300),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_305),
.B2(n_319),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_304),
.C(n_319),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_306),
.B(n_312),
.C(n_313),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_322),
.B(n_323),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_348),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_345),
.B1(n_346),
.B2(n_347),
.Y(n_324)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_336),
.B2(n_337),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_327),
.B(n_336),
.Y(n_471)
);

OAI32xp33_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.A3(n_331),
.B1(n_333),
.B2(n_335),
.Y(n_327)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_342),
.Y(n_382)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_345),
.B(n_346),
.C(n_348),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_359),
.B2(n_369),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_349),
.B(n_360),
.C(n_364),
.Y(n_484)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_359),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_364),
.Y(n_359)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_361),
.Y(n_473)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_363),
.Y(n_394)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_461),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_SL g494 ( 
.A1(n_372),
.A2(n_461),
.B(n_495),
.C(n_498),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_433),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_373),
.B(n_433),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_403),
.C(n_420),
.Y(n_373)
);

FAx1_ASAP7_75t_L g474 ( 
.A(n_374),
.B(n_403),
.CI(n_420),
.CON(n_474),
.SN(n_474)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_389),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_375),
.B(n_390),
.C(n_401),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_385),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_376),
.B(n_385),
.Y(n_467)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_386),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_401),
.Y(n_389)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_SL g393 ( 
.A(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_395),
.Y(n_440)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_415),
.B2(n_419),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_415),
.Y(n_451)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx8_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_415),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_415),
.A2(n_419),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_415),
.A2(n_451),
.B(n_454),
.Y(n_502)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_426),
.C(n_431),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_424),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_422),
.B(n_424),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_426),
.A2(n_427),
.B1(n_431),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_431),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_434),
.B(n_437),
.C(n_449),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_449),
.B2(n_450),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_445),
.B(n_448),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_439),
.B(n_446),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_441),
.Y(n_510)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g501 ( 
.A(n_448),
.B(n_502),
.CI(n_503),
.CON(n_501),
.SN(n_501)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_448),
.B(n_502),
.C(n_503),
.Y(n_523)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_460),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_456),
.Y(n_506)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_474),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_462),
.B(n_474),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_467),
.C(n_468),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_463),
.A2(n_464),
.B1(n_467),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_467),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.C(n_472),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_471),
.B(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_472),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_474),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_488),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_477),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_485),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_478),
.B(n_485),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.C(n_484),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_491),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_484),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_490),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_513),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_512),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_512),
.Y(n_525)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_501),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B1(n_507),
.B2(n_511),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_504),
.A2(n_505),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_515),
.C(n_519),
.Y(n_531)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_507),
.Y(n_511)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_513),
.A2(n_525),
.B(n_526),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_523),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_523),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_531),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_531),
.Y(n_532)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_538),
.Y(n_537)
);


endmodule