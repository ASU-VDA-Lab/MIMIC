module fake_jpeg_4362_n_186 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_186);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx12_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx5_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_27),
.B(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_13),
.B1(n_22),
.B2(n_15),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_17),
.B(n_18),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_23),
.A2(n_22),
.B1(n_13),
.B2(n_12),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_27),
.B1(n_12),
.B2(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_40),
.B(n_29),
.C(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_48),
.A2(n_51),
.B1(n_38),
.B2(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_50),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_41),
.B1(n_35),
.B2(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_30),
.C(n_25),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_36),
.C(n_35),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_69),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_45),
.Y(n_79)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_49),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_32),
.B(n_36),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_61),
.C(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_54),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_47),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_53),
.C(n_51),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_64),
.B(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_51),
.B1(n_47),
.B2(n_52),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_51),
.B1(n_66),
.B2(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_87),
.A2(n_92),
.B1(n_77),
.B2(n_80),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_76),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_65),
.B1(n_64),
.B2(n_62),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_86),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_74),
.B(n_79),
.Y(n_96)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_84),
.CI(n_75),
.CON(n_103),
.SN(n_103)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_68),
.B(n_46),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_106),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_110),
.B(n_115),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_80),
.B(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_97),
.C(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_71),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_114),
.B(n_60),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

OAI322xp33_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_88),
.A3(n_97),
.B1(n_96),
.B2(n_94),
.C1(n_93),
.C2(n_85),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_125),
.C(n_130),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_109),
.A2(n_98),
.B(n_71),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_101),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_110),
.A2(n_18),
.B(n_91),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_112),
.B(n_16),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_44),
.B1(n_38),
.B2(n_60),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_127),
.B1(n_102),
.B2(n_108),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_50),
.C(n_100),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_106),
.A2(n_38),
.B1(n_60),
.B2(n_33),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_0),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_36),
.C(n_30),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_117),
.A2(n_103),
.B1(n_115),
.B2(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_14),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_135),
.B(n_141),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_143),
.B(n_120),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_30),
.C(n_33),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_128),
.C(n_127),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_58),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_142),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_139),
.A2(n_140),
.B1(n_122),
.B2(n_7),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_33),
.B1(n_58),
.B2(n_24),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_125),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_153),
.B(n_131),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_147),
.C(n_149),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_119),
.C(n_121),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_6),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_134),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_152),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_132),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_157),
.A2(n_162),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_160),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_14),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_163),
.Y(n_165)
);

FAx1_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_0),
.CI(n_1),
.CON(n_161),
.SN(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_8),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_7),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_148),
.C(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_157),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_169),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_168),
.B(n_171),
.CI(n_8),
.CON(n_177),
.SN(n_177)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_2),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_175),
.B(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_9),
.C(n_10),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_8),
.C(n_9),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_165),
.C(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_177),
.B(n_11),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_180),
.B(n_181),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_2),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_172),
.C(n_184),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_182),
.Y(n_186)
);


endmodule