module fake_jpeg_14088_n_580 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_580);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_580;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_54),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_57),
.Y(n_146)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_58),
.Y(n_156)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_40),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_78),
.Y(n_114)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_28),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_97),
.Y(n_116)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_83),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_32),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_84),
.B(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

BUFx24_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_34),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_25),
.B1(n_37),
.B2(n_43),
.Y(n_131)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_16),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_100),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_15),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_107),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_52),
.Y(n_120)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_38),
.Y(n_104)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_0),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_44),
.B(n_1),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_31),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_111),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_52),
.Y(n_145)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_50),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_119),
.B(n_123),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_120),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_19),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_19),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_127),
.B(n_164),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_50),
.B1(n_23),
.B2(n_31),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_130),
.B(n_153),
.C(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_131),
.A2(n_147),
.B1(n_165),
.B2(n_176),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_145),
.B(n_85),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_112),
.A2(n_23),
.B1(n_43),
.B2(n_37),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_71),
.A2(n_23),
.B1(n_49),
.B2(n_47),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_148),
.A2(n_159),
.B1(n_93),
.B2(n_75),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_55),
.B(n_25),
.Y(n_151)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_81),
.B(n_1),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_67),
.A2(n_52),
.B1(n_49),
.B2(n_47),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_22),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_60),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_61),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_54),
.A2(n_46),
.B1(n_42),
.B2(n_45),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_102),
.B(n_45),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_92),
.B(n_27),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_80),
.B(n_27),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_46),
.Y(n_204)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_186),
.Y(n_296)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_188),
.Y(n_267)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_125),
.A2(n_90),
.B1(n_110),
.B2(n_70),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_190),
.A2(n_158),
.B1(n_5),
.B2(n_6),
.Y(n_294)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_191),
.Y(n_285)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_192),
.Y(n_252)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

BUFx2_ASAP7_75t_SL g256 ( 
.A(n_194),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_149),
.A2(n_82),
.B1(n_65),
.B2(n_98),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_195),
.A2(n_198),
.B1(n_160),
.B2(n_162),
.Y(n_260)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_153),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_197),
.A2(n_204),
.B(n_232),
.Y(n_276)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_200),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_124),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_221),
.Y(n_253)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_207),
.Y(n_263)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_208),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_116),
.B(n_26),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_209),
.B(n_213),
.Y(n_266)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_150),
.Y(n_210)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_211),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_212),
.B(n_140),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_114),
.B(n_24),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_135),
.Y(n_214)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_214),
.Y(n_279)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_215),
.Y(n_280)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_133),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_217),
.Y(n_271)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_117),
.B(n_91),
.C(n_74),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g273 ( 
.A(n_222),
.B(n_126),
.C(n_162),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_118),
.Y(n_223)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_135),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_227),
.A2(n_229),
.B1(n_243),
.B2(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_111),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_228),
.B(n_235),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_231),
.B(n_233),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_144),
.A2(n_2),
.B(n_3),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_128),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_161),
.B(n_2),
.Y(n_235)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_239),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g265 ( 
.A(n_238),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_173),
.Y(n_239)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_242),
.Y(n_298)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_169),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_134),
.Y(n_244)
);

CKINVDCx9p33_ASAP7_75t_R g289 ( 
.A(n_244),
.Y(n_289)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_106),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_246),
.B(n_136),
.Y(n_288)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_247),
.A2(n_248),
.B1(n_175),
.B2(n_157),
.Y(n_278)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_152),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_198),
.A2(n_159),
.B1(n_148),
.B2(n_72),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_251),
.A2(n_260),
.B1(n_196),
.B2(n_244),
.Y(n_308)
);

AO22x1_ASAP7_75t_SL g254 ( 
.A1(n_201),
.A2(n_160),
.B1(n_140),
.B2(n_126),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_254),
.B(n_274),
.Y(n_320)
);

AND2x6_ASAP7_75t_L g259 ( 
.A(n_193),
.B(n_132),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_259),
.B(n_185),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_232),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_212),
.C(n_216),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_201),
.B(n_141),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_187),
.B(n_170),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_223),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_199),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_211),
.A2(n_136),
.B1(n_170),
.B2(n_168),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_221),
.A2(n_168),
.B1(n_163),
.B2(n_94),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_187),
.A2(n_163),
.B1(n_175),
.B2(n_158),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_184),
.B(n_3),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_5),
.Y(n_317)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_305),
.B(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_266),
.B(n_202),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_307),
.B(n_315),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_308),
.A2(n_309),
.B1(n_325),
.B2(n_341),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_251),
.A2(n_195),
.B1(n_241),
.B2(n_247),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g362 ( 
.A1(n_310),
.A2(n_317),
.B(n_11),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_258),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_253),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_240),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_316),
.B(n_318),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_267),
.B(n_239),
.Y(n_318)
);

OAI22x1_ASAP7_75t_SL g319 ( 
.A1(n_259),
.A2(n_261),
.B1(n_299),
.B2(n_254),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_319),
.A2(n_332),
.B1(n_333),
.B2(n_255),
.Y(n_357)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_263),
.Y(n_321)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_321),
.Y(n_368)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_271),
.Y(n_323)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_287),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_324),
.B(n_340),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_272),
.A2(n_189),
.B1(n_237),
.B2(n_229),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_270),
.Y(n_326)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_326),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_289),
.A2(n_203),
.B1(n_186),
.B2(n_238),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_281),
.Y(n_329)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_289),
.A2(n_223),
.B1(n_227),
.B2(n_8),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_268),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_294),
.A2(n_274),
.B1(n_273),
.B2(n_276),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_334),
.Y(n_351)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_335),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_254),
.A2(n_5),
.B(n_7),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_336),
.A2(n_269),
.B(n_283),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_249),
.B(n_9),
.C(n_10),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_249),
.B(n_9),
.C(n_10),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_267),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_345),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_285),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_305),
.A2(n_262),
.B1(n_285),
.B2(n_255),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_347),
.A2(n_361),
.B1(n_365),
.B2(n_369),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_275),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_375),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_318),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_350),
.B(n_355),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_331),
.Y(n_355)
);

OAI21xp33_ASAP7_75t_SL g356 ( 
.A1(n_320),
.A2(n_296),
.B(n_297),
.Y(n_356)
);

AO21x1_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_357),
.B(n_325),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_332),
.A2(n_250),
.B1(n_271),
.B2(n_286),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_304),
.B1(n_311),
.B2(n_323),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_308),
.A2(n_250),
.B1(n_286),
.B2(n_256),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_310),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_309),
.A2(n_301),
.B1(n_319),
.B2(n_336),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_306),
.A2(n_329),
.B1(n_322),
.B2(n_303),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_315),
.Y(n_375)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_379),
.Y(n_419)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_381),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_345),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_383),
.B(n_399),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_310),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_397),
.C(n_400),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g423 ( 
.A(n_386),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_312),
.Y(n_387)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_387),
.Y(n_434)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_316),
.C(n_317),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_388),
.B(n_342),
.C(n_372),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_348),
.B(n_353),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_377),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_390),
.A2(n_398),
.B1(n_412),
.B2(n_374),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_391),
.A2(n_394),
.B1(n_402),
.B2(n_351),
.Y(n_417)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_349),
.Y(n_392)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_392),
.Y(n_442)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_357),
.A2(n_300),
.B1(n_302),
.B2(n_326),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_396),
.B(n_403),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_328),
.Y(n_397)
);

AOI32xp33_ASAP7_75t_L g398 ( 
.A1(n_375),
.A2(n_334),
.A3(n_335),
.B1(n_339),
.B2(n_338),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_367),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_321),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_367),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_405),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_358),
.A2(n_314),
.B1(n_333),
.B2(n_307),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_376),
.B(n_297),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_404),
.B(n_410),
.C(n_377),
.Y(n_429)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_341),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_406),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_364),
.B(n_283),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_408),
.Y(n_444)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_340),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_409),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_252),
.C(n_296),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_343),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_350),
.B(n_337),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_413),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_403),
.A2(n_411),
.B1(n_390),
.B2(n_382),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_414),
.A2(n_415),
.B1(n_402),
.B2(n_413),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_411),
.A2(n_346),
.B1(n_365),
.B2(n_373),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_395),
.A2(n_346),
.B1(n_363),
.B2(n_361),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_416),
.A2(n_420),
.B(n_437),
.Y(n_447)
);

OAI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_417),
.A2(n_438),
.B1(n_257),
.B2(n_252),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_395),
.A2(n_359),
.B(n_363),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_387),
.A2(n_344),
.B(n_371),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_426),
.B(n_427),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_385),
.A2(n_371),
.B(n_351),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_428),
.B(n_429),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_380),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_433),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_380),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_440),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_385),
.B(n_372),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_436),
.B(n_406),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_394),
.A2(n_342),
.B(n_374),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_386),
.A2(n_342),
.B1(n_374),
.B2(n_366),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_384),
.B(n_397),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_441),
.B(n_446),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_410),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_409),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_386),
.A2(n_268),
.B(n_277),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_418),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_455),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_425),
.Y(n_451)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_400),
.Y(n_452)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_453),
.Y(n_499)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_444),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_464),
.B1(n_465),
.B2(n_469),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_425),
.B(n_404),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_458),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_439),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_460),
.Y(n_488)
);

AO22x1_ASAP7_75t_SL g460 ( 
.A1(n_434),
.A2(n_389),
.B1(n_396),
.B2(n_379),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_461),
.B(n_463),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_439),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_434),
.Y(n_464)
);

INVx13_ASAP7_75t_L g465 ( 
.A(n_426),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_415),
.A2(n_388),
.B1(n_257),
.B2(n_284),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_466),
.A2(n_416),
.B1(n_417),
.B2(n_457),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_431),
.B(n_284),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_467),
.B(n_419),
.Y(n_495)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_471),
.A2(n_414),
.B1(n_421),
.B2(n_420),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_290),
.C(n_265),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_429),
.C(n_440),
.Y(n_481)
);

NOR4xp25_ASAP7_75t_L g473 ( 
.A(n_433),
.B(n_268),
.C(n_264),
.D(n_265),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_473),
.A2(n_474),
.B1(n_475),
.B2(n_438),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_430),
.B(n_268),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_442),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_437),
.Y(n_477)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_489),
.C(n_461),
.Y(n_502)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_482),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_483),
.A2(n_500),
.B1(n_475),
.B2(n_469),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_470),
.B(n_422),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g507 ( 
.A(n_484),
.B(n_487),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_486),
.A2(n_463),
.B1(n_456),
.B2(n_453),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_468),
.B(n_435),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_472),
.B(n_443),
.C(n_428),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_449),
.A2(n_421),
.B1(n_445),
.B2(n_442),
.Y(n_490)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_490),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_448),
.A2(n_445),
.B1(n_423),
.B2(n_419),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_470),
.B(n_427),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_455),
.A2(n_446),
.B1(n_290),
.B2(n_264),
.Y(n_496)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_496),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_277),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_464),
.A2(n_277),
.B1(n_265),
.B2(n_14),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_476),
.B(n_454),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_501),
.B(n_502),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_483),
.A2(n_462),
.B(n_465),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_503),
.A2(n_514),
.B(n_450),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_476),
.B(n_456),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_504),
.B(n_505),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_481),
.B(n_466),
.C(n_447),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_498),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_508),
.B(n_510),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_512),
.A2(n_477),
.B1(n_486),
.B2(n_518),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_477),
.A2(n_447),
.B(n_450),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_515),
.A2(n_460),
.B1(n_467),
.B2(n_485),
.Y(n_533)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_478),
.Y(n_519)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_519),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_489),
.C(n_484),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_521),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_506),
.A2(n_491),
.B1(n_499),
.B2(n_488),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_515),
.Y(n_522)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_522),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_488),
.B1(n_485),
.B2(n_498),
.Y(n_523)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_524),
.A2(n_509),
.B(n_512),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_480),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_525),
.B(n_535),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_493),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_533),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_497),
.C(n_494),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g544 ( 
.A1(n_528),
.A2(n_514),
.B(n_518),
.Y(n_544)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_519),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_474),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_532),
.B(n_503),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_460),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_487),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_536),
.B(n_507),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g561 ( 
.A(n_539),
.B(n_543),
.Y(n_561)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_529),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_541),
.B(n_495),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_511),
.C(n_507),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_548),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_533),
.Y(n_559)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_545),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_546),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_531),
.A2(n_509),
.B(n_511),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_547),
.A2(n_528),
.B(n_536),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_526),
.B(n_500),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_534),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_551),
.A2(n_537),
.B(n_550),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_538),
.A2(n_534),
.B(n_524),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_552),
.B(n_558),
.Y(n_564)
);

OA21x2_ASAP7_75t_SL g554 ( 
.A1(n_542),
.A2(n_522),
.B(n_527),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_554),
.B(n_540),
.Y(n_563)
);

A2O1A1Ixp33_ASAP7_75t_SL g567 ( 
.A1(n_555),
.A2(n_545),
.B(n_473),
.C(n_14),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_540),
.B(n_532),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_559),
.B(n_539),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_560),
.B(n_543),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_562),
.B(n_563),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_566),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_567),
.B(n_551),
.C(n_556),
.Y(n_570)
);

INVx6_ASAP7_75t_L g568 ( 
.A(n_557),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_568),
.A2(n_553),
.B(n_559),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_570),
.B(n_561),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_571),
.A2(n_564),
.B(n_562),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_573),
.B(n_574),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_575),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_569),
.B(n_572),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_577),
.A2(n_561),
.B1(n_567),
.B2(n_14),
.Y(n_578)
);

MAJx2_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_12),
.C(n_13),
.Y(n_579)
);

AO21x1_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_12),
.B(n_448),
.Y(n_580)
);


endmodule