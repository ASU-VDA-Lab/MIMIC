module fake_jpeg_10198_n_56 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_56);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_56;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_32;

INVx2_ASAP7_75t_SL g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_34),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_3),
.B(n_28),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_1),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_2),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_39),
.B(n_42),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_43),
.B(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_5),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_26),
.B1(n_25),
.B2(n_27),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_48),
.C(n_9),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_38),
.B1(n_41),
.B2(n_40),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_7),
.B(n_8),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_49),
.B2(n_45),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.C(n_18),
.Y(n_54)
);

OAI321xp33_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_16),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_37),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_55),
.Y(n_56)
);


endmodule