module real_aes_15731_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g108 ( .A(n_0), .B(n_109), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_1), .A2(n_4), .B1(n_282), .B2(n_283), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_2), .A2(n_43), .B1(n_183), .B2(n_231), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_3), .A2(n_24), .B1(n_231), .B2(n_265), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_16), .B1(n_532), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_6), .A2(n_62), .B1(n_168), .B2(n_169), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_7), .A2(n_17), .B1(n_183), .B2(n_184), .Y(n_182) );
INVx1_ASAP7_75t_L g109 ( .A(n_8), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_9), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_10), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_11), .A2(n_18), .B1(n_533), .B2(n_577), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_12), .A2(n_66), .B1(n_141), .B2(n_142), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_12), .Y(n_141) );
BUFx2_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
OR2x2_ASAP7_75t_L g130 ( .A(n_13), .B(n_38), .Y(n_130) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_14), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g561 ( .A(n_15), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_19), .A2(n_99), .B1(n_283), .B2(n_532), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_20), .A2(n_39), .B1(n_161), .B2(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_21), .B(n_159), .Y(n_593) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_22), .A2(n_60), .B(n_174), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_23), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_25), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_26), .B(n_156), .Y(n_223) );
INVx4_ASAP7_75t_R g207 ( .A(n_27), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_28), .A2(n_47), .B1(n_187), .B2(n_280), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_29), .A2(n_55), .B1(n_187), .B2(n_532), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_30), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_31), .B(n_557), .Y(n_595) );
CKINVDCx5p33_ASAP7_75t_R g538 ( .A(n_32), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_33), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g287 ( .A(n_34), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_SL g262 ( .A1(n_35), .A2(n_155), .B(n_183), .C(n_263), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_36), .A2(n_56), .B1(n_183), .B2(n_187), .Y(n_271) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_37), .Y(n_810) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_40), .A2(n_87), .B1(n_183), .B2(n_524), .Y(n_523) );
OAI22xp5_ASAP7_75t_SL g828 ( .A1(n_41), .A2(n_54), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_41), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_42), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_44), .A2(n_46), .B1(n_183), .B2(n_184), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_45), .A2(n_61), .B1(n_532), .B2(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g227 ( .A(n_48), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_49), .B(n_183), .Y(n_229) );
INVx1_ASAP7_75t_L g832 ( .A(n_50), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_51), .Y(n_241) );
INVx2_ASAP7_75t_L g135 ( .A(n_52), .Y(n_135) );
INVx1_ASAP7_75t_L g111 ( .A(n_53), .Y(n_111) );
BUFx3_ASAP7_75t_L g138 ( .A(n_53), .Y(n_138) );
INVx1_ASAP7_75t_L g829 ( .A(n_54), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_57), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_58), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g186 ( .A1(n_59), .A2(n_88), .B1(n_183), .B2(n_187), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_63), .A2(n_76), .B1(n_280), .B2(n_549), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_64), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_65), .A2(n_79), .B1(n_183), .B2(n_184), .Y(n_534) );
INVx1_ASAP7_75t_L g142 ( .A(n_66), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_67), .A2(n_98), .B1(n_532), .B2(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g174 ( .A(n_68), .Y(n_174) );
AND2x4_ASAP7_75t_L g177 ( .A(n_69), .B(n_178), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_70), .A2(n_90), .B1(n_187), .B2(n_280), .Y(n_279) );
AO22x1_ASAP7_75t_L g157 ( .A1(n_71), .A2(n_77), .B1(n_158), .B2(n_161), .Y(n_157) );
INVx1_ASAP7_75t_L g178 ( .A(n_72), .Y(n_178) );
AND2x2_ASAP7_75t_L g266 ( .A(n_73), .B(n_219), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_74), .B(n_168), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_75), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_78), .B(n_231), .Y(n_242) );
INVx2_ASAP7_75t_L g156 ( .A(n_80), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_81), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_82), .B(n_219), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_83), .A2(n_97), .B1(n_168), .B2(n_187), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_84), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_85), .B(n_172), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_86), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_89), .B(n_219), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_91), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_92), .B(n_219), .Y(n_238) );
INVx1_ASAP7_75t_L g113 ( .A(n_93), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_93), .B(n_128), .Y(n_127) );
NAND2xp33_ASAP7_75t_L g596 ( .A(n_94), .B(n_159), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_95), .A2(n_168), .B(n_189), .C(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g212 ( .A(n_96), .B(n_213), .Y(n_212) );
NAND2xp33_ASAP7_75t_L g246 ( .A(n_100), .B(n_208), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_118), .B(n_831), .Y(n_101) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx4_ASAP7_75t_L g833 ( .A(n_104), .Y(n_833) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_114), .Y(n_105) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .C(n_112), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g504 ( .A(n_113), .Y(n_504) );
NOR2x1p5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2x1p5_ASAP7_75t_L g118 ( .A(n_119), .B(n_817), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_131), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_121), .A2(n_823), .B(n_825), .Y(n_822) );
NOR2x1_ASAP7_75t_R g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx3_ASAP7_75t_L g824 ( .A(n_124), .Y(n_824) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
CKINVDCx8_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
AND2x6_ASAP7_75t_SL g126 ( .A(n_127), .B(n_129), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_129), .B(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_130), .B(n_138), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_809), .Y(n_131) );
BUFx12f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x6_ASAP7_75t_SL g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_135), .B(n_814), .Y(n_813) );
INVx3_ASAP7_75t_L g821 ( .A(n_135), .Y(n_821) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OAI22xp33_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_143), .B1(n_144), .B2(n_808), .Y(n_139) );
INVx1_ASAP7_75t_L g808 ( .A(n_140), .Y(n_808) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_502), .B1(n_505), .B2(n_807), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_412), .Y(n_146) );
NOR3xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_341), .C(n_383), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_149), .B(n_315), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_214), .B1(n_290), .B2(n_301), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OR2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_195), .Y(n_151) );
AOI21xp33_ASAP7_75t_L g334 ( .A1(n_152), .A2(n_335), .B(n_337), .Y(n_334) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_152), .A2(n_408), .B(n_409), .Y(n_407) );
OR2x2_ASAP7_75t_L g152 ( .A(n_153), .B(n_179), .Y(n_152) );
INVx2_ASAP7_75t_L g327 ( .A(n_153), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_153), .B(n_180), .Y(n_357) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_163), .C(n_175), .Y(n_154) );
INVx6_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_155), .A2(n_246), .B(n_247), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_155), .B(n_157), .Y(n_299) );
O2A1O1Ixp5_ASAP7_75t_L g591 ( .A1(n_155), .A2(n_184), .B(n_592), .C(n_593), .Y(n_591) );
BUFx8_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g166 ( .A(n_156), .Y(n_166) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
INVx1_ASAP7_75t_L g226 ( .A(n_156), .Y(n_226) );
INVxp67_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g532 ( .A(n_159), .Y(n_532) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g162 ( .A(n_160), .Y(n_162) );
INVx1_ASAP7_75t_L g168 ( .A(n_160), .Y(n_168) );
INVx1_ASAP7_75t_L g170 ( .A(n_160), .Y(n_170) );
INVx3_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_160), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_160), .Y(n_209) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_160), .Y(n_231) );
INVx1_ASAP7_75t_L g259 ( .A(n_160), .Y(n_259) );
INVx2_ASAP7_75t_L g265 ( .A(n_160), .Y(n_265) );
OAI21xp33_ASAP7_75t_SL g222 ( .A1(n_161), .A2(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g298 ( .A(n_163), .Y(n_298) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_171), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_164), .A2(n_229), .B(n_230), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_164), .A2(n_185), .B1(n_270), .B2(n_271), .Y(n_269) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g515 ( .A(n_165), .Y(n_515) );
BUFx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g244 ( .A(n_166), .Y(n_244) );
INVx1_ASAP7_75t_L g577 ( .A(n_169), .Y(n_577) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_170), .B(n_204), .Y(n_203) );
OAI21xp33_ASAP7_75t_L g175 ( .A1(n_171), .A2(n_172), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g190 ( .A(n_172), .Y(n_190) );
INVx2_ASAP7_75t_L g194 ( .A(n_172), .Y(n_194) );
INVx2_ASAP7_75t_L g200 ( .A(n_172), .Y(n_200) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_173), .Y(n_220) );
INVx1_ASAP7_75t_L g300 ( .A(n_175), .Y(n_300) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_176), .A2(n_255), .B(n_262), .Y(n_254) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx10_ASAP7_75t_L g191 ( .A(n_177), .Y(n_191) );
BUFx10_ASAP7_75t_L g233 ( .A(n_177), .Y(n_233) );
INVx1_ASAP7_75t_L g285 ( .A(n_177), .Y(n_285) );
AND2x2_ASAP7_75t_L g397 ( .A(n_179), .B(n_236), .Y(n_397) );
INVx1_ASAP7_75t_L g430 ( .A(n_179), .Y(n_430) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g292 ( .A(n_180), .B(n_237), .Y(n_292) );
AND2x2_ASAP7_75t_L g323 ( .A(n_180), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g332 ( .A(n_180), .Y(n_332) );
OR2x2_ASAP7_75t_L g351 ( .A(n_180), .B(n_197), .Y(n_351) );
AND2x2_ASAP7_75t_L g366 ( .A(n_180), .B(n_197), .Y(n_366) );
AO31x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_190), .A3(n_191), .B(n_192), .Y(n_180) );
OAI22x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_185), .B1(n_186), .B2(n_188), .Y(n_181) );
INVx4_ASAP7_75t_L g184 ( .A(n_183), .Y(n_184) );
INVx1_ASAP7_75t_L g533 ( .A(n_183), .Y(n_533) );
INVx1_ASAP7_75t_L g549 ( .A(n_183), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_184), .A2(n_241), .B(n_242), .C(n_243), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_185), .A2(n_188), .B1(n_279), .B2(n_281), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_185), .A2(n_514), .B1(n_515), .B2(n_516), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_185), .A2(n_188), .B1(n_523), .B2(n_525), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_185), .A2(n_531), .B1(n_534), .B2(n_535), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_185), .A2(n_515), .B1(n_547), .B2(n_548), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_185), .A2(n_515), .B1(n_556), .B2(n_558), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_185), .A2(n_515), .B1(n_566), .B2(n_567), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_185), .A2(n_535), .B1(n_576), .B2(n_578), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_185), .A2(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_187), .B(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g282 ( .A(n_187), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_188), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_SL g535 ( .A(n_189), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_190), .B(n_551), .Y(n_550) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_190), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g211 ( .A(n_191), .Y(n_211) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_191), .A2(n_272), .A3(n_513), .B(n_517), .Y(n_512) );
AO31x2_ASAP7_75t_L g554 ( .A1(n_191), .A2(n_521), .A3(n_555), .B(n_560), .Y(n_554) );
AO31x2_ASAP7_75t_L g574 ( .A1(n_191), .A2(n_253), .A3(n_575), .B(n_579), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
INVx2_ASAP7_75t_L g213 ( .A(n_194), .Y(n_213) );
BUFx2_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_194), .B(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_194), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_196), .B(n_365), .Y(n_408) );
OR2x2_ASAP7_75t_L g496 ( .A(n_196), .B(n_357), .Y(n_496) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g324 ( .A(n_197), .Y(n_324) );
AND2x2_ASAP7_75t_L g333 ( .A(n_197), .B(n_296), .Y(n_333) );
AND2x2_ASAP7_75t_L g336 ( .A(n_197), .B(n_237), .Y(n_336) );
AND2x2_ASAP7_75t_L g355 ( .A(n_197), .B(n_236), .Y(n_355) );
AND2x4_ASAP7_75t_L g374 ( .A(n_197), .B(n_297), .Y(n_374) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_201), .B(n_212), .Y(n_197) );
AO31x2_ASAP7_75t_L g545 ( .A1(n_198), .A2(n_536), .A3(n_546), .B(n_550), .Y(n_545) );
AO31x2_ASAP7_75t_L g564 ( .A1(n_198), .A2(n_284), .A3(n_565), .B(n_568), .Y(n_564) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_200), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_SL g579 ( .A(n_200), .B(n_580), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_205), .B(n_211), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_206) );
INVx2_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
INVx1_ASAP7_75t_L g557 ( .A(n_208), .Y(n_557) );
INVx1_ASAP7_75t_L g559 ( .A(n_209), .Y(n_559) );
INVx1_ASAP7_75t_L g536 ( .A(n_211), .Y(n_536) );
OAI21xp33_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_234), .B(n_275), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_215), .B(n_369), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_217), .B(n_289), .Y(n_288) );
INVx3_ASAP7_75t_L g305 ( .A(n_217), .Y(n_305) );
OR2x2_ASAP7_75t_L g313 ( .A(n_217), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_217), .B(n_306), .Y(n_338) );
AND2x2_ASAP7_75t_L g363 ( .A(n_217), .B(n_277), .Y(n_363) );
AND2x2_ASAP7_75t_L g381 ( .A(n_217), .B(n_311), .Y(n_381) );
INVx1_ASAP7_75t_L g420 ( .A(n_217), .Y(n_420) );
AND2x2_ASAP7_75t_L g422 ( .A(n_217), .B(n_423), .Y(n_422) );
NAND2x1p5_ASAP7_75t_SL g441 ( .A(n_217), .B(n_362), .Y(n_441) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_221), .Y(n_217) );
NOR2x1_ASAP7_75t_L g248 ( .A(n_219), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g272 ( .A(n_219), .Y(n_272) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g232 ( .A(n_220), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_220), .B(n_518), .Y(n_517) );
BUFx3_ASAP7_75t_L g521 ( .A(n_220), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_220), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_220), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_SL g589 ( .A(n_220), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .B(n_232), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
BUFx4f_ASAP7_75t_L g261 ( .A(n_226), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_231), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g249 ( .A(n_233), .Y(n_249) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_233), .A2(n_269), .A3(n_272), .B(n_273), .Y(n_268) );
OAI32xp33_ASAP7_75t_L g325 ( .A1(n_234), .A2(n_317), .A3(n_326), .B1(n_328), .B2(n_330), .Y(n_325) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_250), .Y(n_234) );
INVx1_ASAP7_75t_L g365 ( .A(n_235), .Y(n_365) );
AND2x2_ASAP7_75t_L g373 ( .A(n_235), .B(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g372 ( .A(n_236), .B(n_296), .Y(n_372) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
BUFx3_ASAP7_75t_L g322 ( .A(n_237), .Y(n_322) );
AND2x2_ASAP7_75t_L g331 ( .A(n_237), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g437 ( .A(n_237), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_245), .B(n_248), .Y(n_239) );
INVx2_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g307 ( .A(n_250), .Y(n_307) );
OR2x2_ASAP7_75t_L g317 ( .A(n_250), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g439 ( .A(n_250), .Y(n_439) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_267), .Y(n_250) );
AND2x2_ASAP7_75t_L g340 ( .A(n_251), .B(n_268), .Y(n_340) );
INVx2_ASAP7_75t_L g362 ( .A(n_251), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_251), .B(n_277), .Y(n_382) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g289 ( .A(n_252), .Y(n_289) );
AOI21x1_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_266), .Y(n_252) );
AO31x2_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_278), .A3(n_284), .B(n_286), .Y(n_277) );
AO31x2_ASAP7_75t_L g529 ( .A1(n_253), .A2(n_530), .A3(n_536), .B(n_537), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_258), .B(n_261), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g283 ( .A(n_259), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_SL g524 ( .A(n_265), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_267), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g371 ( .A(n_267), .Y(n_371) );
INVx2_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g311 ( .A(n_268), .Y(n_311) );
OR2x2_ASAP7_75t_L g377 ( .A(n_268), .B(n_277), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_268), .B(n_277), .Y(n_410) );
INVx2_ASAP7_75t_L g358 ( .A(n_275), .Y(n_358) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_288), .Y(n_275) );
OR2x2_ASAP7_75t_L g345 ( .A(n_276), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g423 ( .A(n_276), .Y(n_423) );
INVx1_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
INVx1_ASAP7_75t_L g314 ( .A(n_277), .Y(n_314) );
INVx1_ASAP7_75t_L g329 ( .A(n_277), .Y(n_329) );
AO31x2_ASAP7_75t_L g520 ( .A1(n_284), .A2(n_521), .A3(n_522), .B(n_526), .Y(n_520) );
INVx2_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_SL g597 ( .A(n_285), .Y(n_597) );
OR2x2_ASAP7_75t_L g433 ( .A(n_288), .B(n_410), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_289), .B(n_305), .Y(n_346) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_289), .Y(n_348) );
OR2x2_ASAP7_75t_L g447 ( .A(n_289), .B(n_371), .Y(n_447) );
INVxp67_ASAP7_75t_L g471 ( .A(n_289), .Y(n_471) );
INVx2_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
NAND2x1_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_292), .B(n_333), .Y(n_400) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g349 ( .A(n_294), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g462 ( .A(n_295), .Y(n_462) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g491 ( .A(n_296), .B(n_324), .Y(n_491) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g417 ( .A(n_297), .B(n_324), .Y(n_417) );
AOI21x1_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_300), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_304), .B(n_340), .Y(n_454) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g318 ( .A(n_305), .Y(n_318) );
AND2x2_ASAP7_75t_L g368 ( .A(n_305), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_305), .B(n_362), .Y(n_411) );
OR2x2_ASAP7_75t_L g483 ( .A(n_305), .B(n_370), .Y(n_483) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g394 ( .A(n_310), .Y(n_394) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g384 ( .A(n_313), .B(n_385), .Y(n_384) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_313), .Y(n_395) );
OR2x2_ASAP7_75t_L g446 ( .A(n_313), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g501 ( .A(n_313), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B(n_325), .C(n_334), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g390 ( .A(n_318), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_318), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g463 ( .A(n_318), .B(n_340), .Y(n_463) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_321), .B(n_366), .Y(n_388) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_321), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g473 ( .A(n_321), .B(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g416 ( .A(n_322), .Y(n_416) );
AND2x2_ASAP7_75t_L g444 ( .A(n_323), .B(n_372), .Y(n_444) );
INVx2_ASAP7_75t_L g467 ( .A(n_323), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_323), .B(n_365), .Y(n_499) );
AND2x4_ASAP7_75t_SL g453 ( .A(n_326), .B(n_331), .Y(n_453) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g406 ( .A(n_327), .B(n_332), .Y(n_406) );
OR2x2_ASAP7_75t_L g458 ( .A(n_327), .B(n_351), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_328), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_328), .B(n_340), .Y(n_494) );
BUFx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g442 ( .A(n_329), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
INVx1_ASAP7_75t_L g425 ( .A(n_331), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_331), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g475 ( .A(n_332), .Y(n_475) );
BUFx2_ASAP7_75t_L g343 ( .A(n_333), .Y(n_343) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g461 ( .A(n_336), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_340), .Y(n_402) );
NAND3xp33_ASAP7_75t_SL g341 ( .A(n_342), .B(n_352), .C(n_367), .Y(n_341) );
AOI22xp33_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_344), .B1(n_347), .B2(n_349), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g455 ( .A1(n_349), .A2(n_375), .B1(n_456), .B2(n_459), .C1(n_461), .C2(n_463), .Y(n_455) );
AND2x2_ASAP7_75t_L g487 ( .A(n_350), .B(n_436), .Y(n_487) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g435 ( .A(n_351), .B(n_436), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_358), .B1(n_359), .B2(n_364), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx2_ASAP7_75t_SL g431 ( .A(n_355), .Y(n_431) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
AND2x2_ASAP7_75t_L g418 ( .A(n_360), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g376 ( .A(n_361), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g370 ( .A(n_362), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g485 ( .A(n_363), .Y(n_485) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_366), .B(n_462), .Y(n_481) );
INVx1_ASAP7_75t_L g498 ( .A(n_366), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_372), .B1(n_373), .B2(n_375), .C1(n_378), .C2(n_379), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_374), .Y(n_378) );
AND2x2_ASAP7_75t_L g396 ( .A(n_374), .B(n_397), .Y(n_396) );
INVx3_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g391 ( .A(n_377), .Y(n_391) );
OR2x2_ASAP7_75t_L g460 ( .A(n_377), .B(n_441), .Y(n_460) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_389), .C(n_398), .Y(n_383) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_396), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_390), .A2(n_428), .B1(n_477), .B2(n_480), .C(n_482), .Y(n_476) );
AND2x4_ASAP7_75t_L g419 ( .A(n_391), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g450 ( .A(n_397), .Y(n_450) );
AOI211x1_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_403), .C(n_407), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g468 ( .A(n_406), .Y(n_468) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_409), .B(n_457), .C(n_458), .Y(n_456) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g492 ( .A(n_410), .Y(n_492) );
NOR2x1_ASAP7_75t_L g412 ( .A(n_413), .B(n_464), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_421), .C(n_443), .D(n_455), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND2x2_ASAP7_75t_L g474 ( .A(n_417), .B(n_475), .Y(n_474) );
AOI221x1_ASAP7_75t_L g443 ( .A1(n_419), .A2(n_444), .B1(n_445), .B2(n_448), .C(n_451), .Y(n_443) );
AND2x2_ASAP7_75t_L g469 ( .A(n_419), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g479 ( .A(n_420), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B1(n_428), .B2(n_432), .C(n_434), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_426), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_431), .A2(n_435), .B1(n_438), .B2(n_440), .Y(n_434) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_435), .A2(n_452), .B(n_454), .Y(n_451) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVxp67_ASAP7_75t_L g478 ( .A(n_447), .Y(n_478) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g497 ( .A1(n_460), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .C(n_488), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_469), .B1(n_472), .B2(n_473), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g484 ( .A(n_471), .B(n_485), .Y(n_484) );
NAND2x1_ASAP7_75t_L g500 ( .A(n_471), .B(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B1(n_493), .B2(n_495), .C(n_497), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g807 ( .A(n_502), .Y(n_807) );
BUFx12f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g815 ( .A(n_504), .B(n_816), .Y(n_815) );
XNOR2xp5_ASAP7_75t_L g827 ( .A(n_505), .B(n_828), .Y(n_827) );
NOR2x1p5_ASAP7_75t_L g505 ( .A(n_506), .B(n_717), .Y(n_505) );
NAND4xp75_ASAP7_75t_L g506 ( .A(n_507), .B(n_662), .C(n_682), .D(n_698), .Y(n_506) );
NOR2x1p5_ASAP7_75t_SL g507 ( .A(n_508), .B(n_632), .Y(n_507) );
NAND4xp75_ASAP7_75t_L g508 ( .A(n_509), .B(n_570), .C(n_609), .D(n_618), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_539), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_519), .Y(n_510) );
AND2x4_ASAP7_75t_L g742 ( .A(n_511), .B(n_669), .Y(n_742) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_512), .Y(n_585) );
INVx2_ASAP7_75t_L g603 ( .A(n_512), .Y(n_603) );
AND2x2_ASAP7_75t_L g626 ( .A(n_512), .B(n_588), .Y(n_626) );
OR2x2_ASAP7_75t_L g681 ( .A(n_512), .B(n_520), .Y(n_681) );
AND2x2_ASAP7_75t_L g599 ( .A(n_519), .B(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g749 ( .A(n_519), .B(n_626), .Y(n_749) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .Y(n_519) );
OR2x2_ASAP7_75t_L g586 ( .A(n_520), .B(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g617 ( .A(n_520), .Y(n_617) );
AND2x2_ASAP7_75t_L g623 ( .A(n_520), .B(n_529), .Y(n_623) );
INVx1_ASAP7_75t_L g641 ( .A(n_520), .Y(n_641) );
INVx2_ASAP7_75t_L g670 ( .A(n_520), .Y(n_670) );
INVx3_ASAP7_75t_L g646 ( .A(n_528), .Y(n_646) );
INVx2_ASAP7_75t_L g651 ( .A(n_528), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_528), .B(n_602), .Y(n_656) );
AND2x2_ASAP7_75t_L g679 ( .A(n_528), .B(n_658), .Y(n_679) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_528), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_528), .B(n_734), .Y(n_733) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g668 ( .A(n_529), .Y(n_668) );
AND2x2_ASAP7_75t_L g716 ( .A(n_529), .B(n_670), .Y(n_716) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_552), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_541), .B(n_660), .Y(n_707) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g704 ( .A(n_542), .B(n_660), .Y(n_704) );
INVx1_ASAP7_75t_L g805 ( .A(n_542), .Y(n_805) );
INVx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g755 ( .A(n_543), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g608 ( .A(n_544), .Y(n_608) );
OR2x2_ASAP7_75t_L g689 ( .A(n_544), .B(n_563), .Y(n_689) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g631 ( .A(n_545), .Y(n_631) );
AND2x4_ASAP7_75t_L g637 ( .A(n_545), .B(n_638), .Y(n_637) );
AOI32xp33_ASAP7_75t_L g775 ( .A1(n_552), .A2(n_678), .A3(n_776), .B1(n_778), .B2(n_779), .Y(n_775) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g724 ( .A(n_553), .B(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_562), .Y(n_553) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_554), .Y(n_572) );
OR2x2_ASAP7_75t_L g606 ( .A(n_554), .B(n_564), .Y(n_606) );
INVx1_ASAP7_75t_L g621 ( .A(n_554), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_554), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g636 ( .A(n_554), .Y(n_636) );
INVx2_ASAP7_75t_L g661 ( .A(n_554), .Y(n_661) );
AND2x2_ASAP7_75t_L g780 ( .A(n_554), .B(n_574), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_562), .B(n_613), .Y(n_700) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g573 ( .A(n_564), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g629 ( .A(n_564), .Y(n_629) );
INVx2_ASAP7_75t_L g638 ( .A(n_564), .Y(n_638) );
AND2x4_ASAP7_75t_L g660 ( .A(n_564), .B(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_564), .Y(n_752) );
AOI22x1_ASAP7_75t_SL g570 ( .A1(n_571), .A2(n_581), .B1(n_599), .B2(n_604), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_573), .B(n_730), .C(n_731), .D(n_732), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_573), .B(n_630), .Y(n_760) );
INVx4_ASAP7_75t_SL g613 ( .A(n_574), .Y(n_613) );
BUFx2_ASAP7_75t_L g676 ( .A(n_574), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_574), .B(n_621), .Y(n_739) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g701 ( .A(n_583), .B(n_650), .Y(n_701) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_L g624 ( .A(n_587), .B(n_602), .Y(n_624) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_588), .B(n_603), .Y(n_648) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_598), .Y(n_588) );
OAI21x1_ASAP7_75t_L g643 ( .A1(n_589), .A2(n_590), .B(n_598), .Y(n_643) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_594), .B(n_597), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_600), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g666 ( .A(n_600), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g705 ( .A(n_601), .B(n_623), .Y(n_705) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g748 ( .A(n_603), .B(n_658), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_604), .A2(n_721), .B1(n_723), .B2(n_726), .C(n_728), .Y(n_720) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g614 ( .A(n_606), .Y(n_614) );
OR2x2_ASAP7_75t_L g714 ( .A(n_606), .B(n_653), .Y(n_714) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_610), .A2(n_736), .B1(n_740), .B2(n_743), .Y(n_735) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
AND2x4_ASAP7_75t_L g659 ( .A(n_611), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g771 ( .A(n_611), .B(n_689), .Y(n_771) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g619 ( .A(n_613), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g635 ( .A(n_613), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g694 ( .A(n_613), .B(n_631), .Y(n_694) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_613), .Y(n_711) );
INVx1_ASAP7_75t_L g725 ( .A(n_613), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_613), .B(n_638), .Y(n_768) );
AND2x4_ASAP7_75t_L g675 ( .A(n_614), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g673 ( .A(n_616), .Y(n_673) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_617), .B(n_658), .Y(n_657) );
NAND2x1_ASAP7_75t_L g777 ( .A(n_617), .B(n_679), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_622), .B1(n_625), .B2(n_627), .Y(n_618) );
AND2x2_ASAP7_75t_L g644 ( .A(n_619), .B(n_637), .Y(n_644) );
INVx1_ASAP7_75t_L g685 ( .A(n_619), .Y(n_685) );
AND2x2_ASAP7_75t_L g792 ( .A(n_619), .B(n_653), .Y(n_792) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x4_ASAP7_75t_SL g622 ( .A(n_623), .B(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g625 ( .A(n_623), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g765 ( .A(n_623), .Y(n_765) );
AND2x2_ASAP7_75t_L g782 ( .A(n_623), .B(n_642), .Y(n_782) );
AND2x2_ASAP7_75t_L g798 ( .A(n_623), .B(n_748), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_624), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g721 ( .A(n_624), .B(n_722), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_624), .A2(n_714), .B1(n_729), .B2(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g684 ( .A(n_626), .Y(n_684) );
AND2x2_ASAP7_75t_L g715 ( .A(n_626), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_626), .B(n_722), .Y(n_744) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g750 ( .A(n_630), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_630), .A2(n_654), .B1(n_759), .B2(n_761), .Y(n_758) );
INVx3_ASAP7_75t_L g653 ( .A(n_631), .Y(n_653) );
AND2x2_ASAP7_75t_L g785 ( .A(n_631), .B(n_638), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_649), .Y(n_632) );
AOI32xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_639), .A3(n_642), .B1(n_644), .B2(n_645), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_636), .Y(n_731) );
INVx1_ASAP7_75t_L g756 ( .A(n_636), .Y(n_756) );
INVx3_ASAP7_75t_L g712 ( .A(n_637), .Y(n_712) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_640), .A2(n_788), .B1(n_789), .B2(n_790), .C(n_791), .Y(n_787) );
BUFx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g764 ( .A(n_642), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g800 ( .A(n_642), .B(n_761), .Y(n_800) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g658 ( .A(n_643), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_645), .B(n_673), .Y(n_672) );
AO22x1_ASAP7_75t_L g702 ( .A1(n_645), .A2(n_703), .B1(n_705), .B2(n_706), .Y(n_702) );
NAND2x1p5_ASAP7_75t_L g806 ( .A(n_645), .B(n_673), .Y(n_806) );
AND2x4_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_L g722 ( .A(n_646), .Y(n_722) );
INVx1_ASAP7_75t_L g732 ( .A(n_646), .Y(n_732) );
AND2x2_ASAP7_75t_L g652 ( .A(n_647), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_648), .Y(n_734) );
INVx1_ASAP7_75t_L g774 ( .A(n_648), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B(n_654), .C(n_659), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NOR2x1p5_ASAP7_75t_L g761 ( .A(n_651), .B(n_681), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_652), .B(n_711), .Y(n_788) );
AOI31xp33_ASAP7_75t_L g671 ( .A1(n_653), .A2(n_672), .A3(n_674), .B(n_677), .Y(n_671) );
INVx4_ASAP7_75t_L g730 ( .A(n_653), .Y(n_730) );
OR2x2_ASAP7_75t_L g767 ( .A(n_653), .B(n_768), .Y(n_767) );
INVx2_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
AND2x4_ASAP7_75t_L g669 ( .A(n_658), .B(n_670), .Y(n_669) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_660), .Y(n_665) );
AND2x2_ASAP7_75t_L g696 ( .A(n_660), .B(n_694), .Y(n_696) );
NOR2xp67_ASAP7_75t_L g662 ( .A(n_663), .B(n_671), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
INVx1_ASAP7_75t_L g789 ( .A(n_666), .Y(n_789) );
INVx1_ASAP7_75t_L g697 ( .A(n_667), .Y(n_697) );
AND2x4_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g727 ( .A(n_668), .Y(n_727) );
AND2x2_ASAP7_75t_L g726 ( .A(n_669), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI322xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_685), .A3(n_686), .B1(n_690), .B2(n_693), .C1(n_695), .C2(n_697), .Y(n_683) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI211x1_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_702), .C(n_708), .Y(n_698) );
INVx1_ASAP7_75t_L g803 ( .A(n_699), .Y(n_803) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g757 ( .A(n_701), .Y(n_757) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OA21x2_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_713), .B(n_715), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx2_ASAP7_75t_L g778 ( .A(n_712), .Y(n_778) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND2xp33_ASAP7_75t_L g773 ( .A(n_716), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_786), .Y(n_717) );
NOR3xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_753), .C(n_769), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_735), .C(n_745), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_722), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI21xp33_ASAP7_75t_L g781 ( .A1(n_726), .A2(n_782), .B(n_783), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g736 ( .A(n_730), .B(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_730), .B(n_780), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_731), .B(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_732), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_742), .A2(n_792), .B(n_793), .Y(n_791) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B(n_750), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI211xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_757), .B(n_758), .C(n_762), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_SL g772 ( .A(n_764), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_768), .Y(n_790) );
OAI211xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_772), .B(n_775), .C(n_781), .Y(n_769) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_780), .B(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g801 ( .A(n_780), .Y(n_801) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g797 ( .A(n_785), .Y(n_797) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_795), .C(n_802), .Y(n_786) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
AOI21xp33_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_799), .B(n_801), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
AOI21xp33_ASAP7_75t_R g802 ( .A1(n_803), .A2(n_804), .B(n_806), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx6_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx10_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_822), .Y(n_817) );
INVxp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
BUFx2_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
BUFx6f_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
endmodule