module real_jpeg_22264_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_0),
.A2(n_6),
.B1(n_24),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_0),
.A2(n_5),
.B1(n_39),
.B2(n_51),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_0),
.A2(n_4),
.B1(n_35),
.B2(n_51),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_5),
.B1(n_39),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_1),
.A2(n_4),
.B1(n_35),
.B2(n_41),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_21),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_2),
.A2(n_10),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_2),
.A2(n_21),
.B(n_26),
.C(n_113),
.Y(n_112)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_9),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_65),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_4),
.A2(n_10),
.B1(n_26),
.B2(n_35),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_4),
.A2(n_9),
.B(n_10),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_5),
.A2(n_9),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_5),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_7),
.B1(n_39),
.B2(n_48),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_10),
.B1(n_26),
.B2(n_39),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_5),
.A2(n_26),
.B(n_36),
.C(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_6),
.A2(n_8),
.B1(n_21),
.B2(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_6),
.A2(n_10),
.B1(n_24),
.B2(n_26),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_6),
.A2(n_7),
.B1(n_24),
.B2(n_48),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_10),
.B(n_114),
.Y(n_113)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_10),
.B(n_24),
.C(n_159),
.Y(n_158)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_10),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_10),
.B(n_49),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_91),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_89),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_73),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_14),
.B(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_60),
.B1(n_61),
.B2(n_72),
.Y(n_14)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_53),
.B2(n_54),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_18),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_18),
.A2(n_62),
.B(n_68),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_57),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_18),
.A2(n_52),
.B1(n_62),
.B2(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_18),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_18),
.A2(n_52),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_18),
.A2(n_57),
.B(n_82),
.C(n_110),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_23),
.Y(n_19)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_23),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_26),
.B(n_34),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_26),
.B(n_79),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_26),
.A2(n_39),
.B(n_48),
.Y(n_159)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_33),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_37),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

OA22x2_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_37),
.B1(n_40),
.B2(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_34),
.A2(n_37),
.B1(n_56),
.B2(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_35),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_58),
.Y(n_81)
);

AOI211xp5_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_80),
.B(n_83),
.C(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_55),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_57),
.A2(n_58),
.B1(n_80),
.B2(n_100),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_57),
.A2(n_100),
.B(n_161),
.C(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_57),
.A2(n_58),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_115),
.C(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_62),
.A2(n_69),
.B1(n_88),
.B2(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_67),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_78),
.B1(n_79),
.B2(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_69),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.C(n_86),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_74),
.A2(n_75),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_81),
.B(n_82),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_76),
.A2(n_108),
.B1(n_109),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_76),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_77),
.A2(n_80),
.B1(n_100),
.B2(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_77),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_100),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_100),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_80),
.A2(n_100),
.B1(n_136),
.B2(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_115),
.C(n_140),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_80),
.A2(n_100),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_80),
.B(n_167),
.C(n_173),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_80),
.B(n_103),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_81),
.A2(n_82),
.B(n_192),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_86),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_209),
.B(n_214),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_199),
.B(n_208),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_129),
.B(n_184),
.C(n_198),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_117),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_95),
.B(n_117),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_101),
.B2(n_102),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_97),
.B(n_102),
.C(n_107),
.Y(n_185)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_99),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_103),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_116),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_108),
.A2(n_109),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_124),
.B1(n_139),
.B2(n_142),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_124),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_115),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_170)
);

NAND2x1_ASAP7_75t_SL g174 ( 
.A(n_115),
.B(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_125),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_118),
.A2(n_119),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_121),
.B1(n_157),
.B2(n_161),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_124),
.B(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_125),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_183),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_176),
.B(n_182),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_163),
.B(n_175),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_154),
.B(n_162),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_143),
.B(n_153),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_139),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_150),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_158),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_164),
.B(n_166),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_171),
.B2(n_172),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_196),
.B2(n_197),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_195),
.C(n_197),
.Y(n_200)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_191),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_192),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_201),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_202),
.B(n_210),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.CI(n_207),
.CON(n_202),
.SN(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);


endmodule