module real_jpeg_24665_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_213;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_49),
.B1(n_52),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_1),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_3),
.A2(n_27),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_3),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_3),
.A2(n_27),
.B1(n_49),
.B2(n_52),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_5),
.A2(n_49),
.B1(n_52),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_5),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_86),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_49),
.B1(n_52),
.B2(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_9),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_9),
.A2(n_43),
.B1(n_49),
.B2(n_52),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_10),
.A2(n_57),
.B1(n_64),
.B2(n_75),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_10),
.A2(n_49),
.B1(n_52),
.B2(n_57),
.Y(n_142)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_12),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_12),
.B(n_66),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_12),
.B(n_36),
.C(n_38),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_12),
.A2(n_28),
.B1(n_31),
.B2(n_69),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_12),
.B(n_41),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_69),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_12),
.B(n_49),
.C(n_51),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_12),
.A2(n_80),
.B(n_173),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_14),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_100)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_132),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_20),
.B(n_103),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_92),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_21),
.A2(n_22),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_58),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_25),
.B(n_44),
.C(n_58),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_26),
.Y(n_94)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_28),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_28),
.A2(n_31),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_28),
.B(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_28),
.B(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_31),
.A2(n_63),
.A3(n_68),
.B1(n_71),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_33),
.A2(n_108),
.B(n_109),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_33),
.A2(n_109),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_34),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_55)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_36),
.B(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_41),
.B(n_96),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_42),
.Y(n_108)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_53),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_46),
.A2(n_48),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_48),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_48),
.A2(n_53),
.B(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_48),
.B(n_69),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_52),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_54),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_56),
.B(n_147),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_73),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_65),
.A2(n_111),
.B(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_69),
.B(n_125),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_77),
.B(n_92),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_90),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_90),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_79),
.A2(n_184),
.B1(n_186),
.B2(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_85),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_80),
.A2(n_172),
.B(n_173),
.Y(n_171)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_99),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_93),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_117),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_129),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_127),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_127),
.A2(n_161),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_210),
.B(n_215),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_162),
.B(n_209),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_151),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_135),
.B(n_151),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.C(n_148),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_136),
.B(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_143),
.A2(n_148),
.B1(n_149),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_146),
.Y(n_160)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_152),
.B(n_158),
.C(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_203),
.B(n_208),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_181),
.B(n_202),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_175),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_175),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_207)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_179),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_191),
.B(n_201),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_189),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_187),
.B(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_196),
.B(n_200),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_194),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_207),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_214),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);


endmodule