module fake_jpeg_7428_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_1),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_0),
.C(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_38),
.Y(n_51)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_54),
.B1(n_61),
.B2(n_29),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_18),
.B1(n_31),
.B2(n_17),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_55),
.B1(n_29),
.B2(n_23),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_56),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_18),
.B1(n_15),
.B2(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_31),
.B1(n_15),
.B2(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_19),
.B1(n_20),
.B2(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

OR2x4_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_30),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_40),
.B1(n_37),
.B2(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_77),
.Y(n_87)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_66),
.Y(n_85)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_42),
.B1(n_39),
.B2(n_40),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_73),
.B1(n_54),
.B2(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_72),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_29),
.B(n_73),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_37),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_41),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_56),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_58),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_84),
.A2(n_77),
.B1(n_64),
.B2(n_33),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_47),
.C(n_56),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_101),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_95),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_71),
.B(n_80),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_72),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_16),
.Y(n_97)
);

NOR3xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_26),
.C(n_19),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_104),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_65),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_47),
.C(n_41),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_14),
.C(n_3),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_26),
.C(n_25),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_68),
.Y(n_108)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_120),
.B(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_117),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_89),
.B1(n_98),
.B2(n_104),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_53),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_100),
.C(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_62),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_20),
.Y(n_126)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_116),
.B1(n_112),
.B2(n_106),
.C(n_114),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_105),
.B1(n_95),
.B2(n_81),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_123),
.B1(n_76),
.B2(n_48),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_86),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_138),
.B(n_130),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_144),
.C(n_123),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_136),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_93),
.C(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_135),
.B(n_2),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_93),
.B(n_87),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_87),
.B1(n_84),
.B2(n_90),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_143),
.B1(n_124),
.B2(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_145),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_94),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_76),
.B1(n_48),
.B2(n_81),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_62),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_129),
.A3(n_134),
.B1(n_132),
.B2(n_139),
.C1(n_137),
.C2(n_33),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_118),
.B1(n_115),
.B2(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_155),
.B1(n_165),
.B2(n_136),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_115),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_129),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_164),
.C(n_131),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_60),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_60),
.Y(n_161)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_60),
.C(n_94),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_172),
.C(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_132),
.C(n_134),
.Y(n_172)
);

NOR4xp25_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_160),
.C(n_157),
.D(n_151),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_60),
.C(n_36),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_149),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_46),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_153),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_177),
.A3(n_179),
.B1(n_176),
.B2(n_180),
.C1(n_167),
.C2(n_21),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_166),
.B(n_159),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_185),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_162),
.B1(n_154),
.B2(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_170),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_175),
.A2(n_165),
.B(n_4),
.Y(n_189)
);

NAND4xp25_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_5),
.C(n_6),
.D(n_9),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_4),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_27),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_27),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_177),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_195),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_198),
.A2(n_197),
.B(n_22),
.Y(n_206)
);

OA21x2_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_181),
.B(n_182),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_183),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_205),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_181),
.B1(n_182),
.B2(n_46),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_199),
.B1(n_24),
.B2(n_46),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_202),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_5),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_22),
.B(n_21),
.C(n_10),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_212),
.A2(n_207),
.B(n_6),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_24),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_204),
.A2(n_199),
.B1(n_205),
.B2(n_208),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_211),
.A2(n_207),
.B(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_5),
.C(n_11),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_11),
.B(n_12),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_213),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_12),
.B(n_13),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_11),
.C(n_12),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_225),
.B(n_220),
.Y(n_226)
);


endmodule