module fake_jpeg_29035_n_412 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_412);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_46),
.Y(n_118)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_17),
.B(n_7),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_48),
.B(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_0),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_35),
.C(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g127 ( 
.A(n_60),
.Y(n_127)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_33),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_71),
.Y(n_114)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_40),
.B(n_8),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_77),
.B(n_83),
.Y(n_138)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_8),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_87),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_65),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_98),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_42),
.B1(n_20),
.B2(n_36),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_106),
.B1(n_126),
.B2(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_41),
.B1(n_44),
.B2(n_39),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_100),
.A2(n_129),
.B1(n_131),
.B2(n_73),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_41),
.B1(n_44),
.B2(n_39),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_105),
.B(n_9),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_57),
.A2(n_42),
.B1(n_36),
.B2(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_16),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_120),
.Y(n_154)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_45),
.B(n_0),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_34),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_46),
.B(n_2),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_50),
.C(n_47),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_58),
.A2(n_42),
.B1(n_34),
.B2(n_31),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_64),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_27),
.B1(n_18),
.B2(n_10),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_78),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_49),
.A2(n_10),
.B1(n_13),
.B2(n_11),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_81),
.B1(n_80),
.B2(n_88),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_60),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_79),
.B1(n_54),
.B2(n_56),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_141),
.A2(n_157),
.B1(n_132),
.B2(n_113),
.Y(n_212)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_144),
.B(n_147),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_67),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_150),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_72),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_60),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_151),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_152),
.B(n_155),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_72),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_153),
.B(n_159),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_101),
.B(n_59),
.Y(n_159)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_62),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_177),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_106),
.B1(n_99),
.B2(n_140),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_70),
.B1(n_76),
.B2(n_75),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_163),
.A2(n_186),
.B1(n_188),
.B2(n_187),
.Y(n_225)
);

INVx5_ASAP7_75t_SL g164 ( 
.A(n_127),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_164),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_118),
.A2(n_66),
.B(n_86),
.Y(n_165)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_185),
.B(n_5),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_113),
.C(n_135),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_94),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_167),
.B(n_175),
.Y(n_224)
);

BUFx8_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

BUFx8_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_109),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_178),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_174),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_116),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_104),
.B(n_13),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_4),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_126),
.Y(n_178)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_107),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_51),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_96),
.B(n_61),
.Y(n_183)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_102),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_184),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_122),
.A2(n_63),
.B1(n_14),
.B2(n_6),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_104),
.B(n_14),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_136),
.A2(n_5),
.B1(n_6),
.B2(n_139),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_96),
.B(n_5),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_93),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_190),
.A2(n_93),
.B1(n_95),
.B2(n_123),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_195),
.B1(n_225),
.B2(n_171),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_193),
.B(n_200),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_140),
.B1(n_135),
.B2(n_132),
.Y(n_195)
);

CKINVDCx12_ASAP7_75t_R g197 ( 
.A(n_168),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_202),
.B(n_212),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_146),
.B(n_107),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_226),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_213),
.A2(n_219),
.B1(n_173),
.B2(n_220),
.Y(n_252)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_143),
.B(n_95),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g266 ( 
.A1(n_214),
.A2(n_198),
.B(n_202),
.C(n_193),
.D(n_210),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_149),
.A2(n_6),
.B1(n_164),
.B2(n_155),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_157),
.A2(n_163),
.B1(n_148),
.B2(n_154),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_223),
.A2(n_186),
.B1(n_188),
.B2(n_167),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_177),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_185),
.B(n_143),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_232),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_150),
.B(n_143),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_166),
.B(n_175),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_158),
.B(n_156),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_152),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_239),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_232),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_235),
.B(n_238),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_237),
.A2(n_240),
.B1(n_263),
.B2(n_218),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_176),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_181),
.B1(n_160),
.B2(n_169),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_245),
.B1(n_252),
.B2(n_233),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_180),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_244),
.B(n_247),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_225),
.A2(n_179),
.B1(n_184),
.B2(n_151),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_172),
.B(n_190),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_246),
.A2(n_256),
.B(n_207),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_142),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_201),
.B(n_173),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_168),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_251),
.B(n_254),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_217),
.B(n_173),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_226),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_201),
.B(n_229),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_261),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_199),
.A2(n_200),
.B(n_214),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_209),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_215),
.B(n_204),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_227),
.A2(n_211),
.B1(n_198),
.B2(n_215),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_210),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_270),
.Y(n_303)
);

OAI21x1_ASAP7_75t_SL g289 ( 
.A1(n_266),
.A2(n_192),
.B(n_207),
.Y(n_289)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_218),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_203),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_282),
.C(n_287),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_237),
.A2(n_220),
.B1(n_222),
.B2(n_233),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_276),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_277),
.A2(n_278),
.B(n_286),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_248),
.A2(n_243),
.B(n_251),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_296),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_242),
.B(n_243),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_238),
.A2(n_222),
.B(n_196),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_290),
.B(n_265),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_280),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_196),
.B(n_207),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_192),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_289),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_294),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_297),
.B1(n_245),
.B2(n_249),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_236),
.B(n_208),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_265),
.A2(n_208),
.B1(n_231),
.B2(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_301),
.Y(n_323)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_302),
.Y(n_325)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_304),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_241),
.B1(n_290),
.B2(n_235),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_305),
.A2(n_311),
.B1(n_318),
.B2(n_328),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_271),
.B(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_309),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_244),
.Y(n_312)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_316),
.A2(n_276),
.B(n_281),
.Y(n_348)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_303),
.B(n_246),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_317),
.A2(n_283),
.B(n_273),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_302),
.A2(n_265),
.B1(n_266),
.B2(n_254),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_247),
.Y(n_319)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_319),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_303),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_321),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_293),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_255),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_326),
.Y(n_339)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_261),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_272),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_256),
.C(n_287),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_336),
.C(n_337),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_320),
.B(n_308),
.C(n_296),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_275),
.C(n_282),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_278),
.C(n_236),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_340),
.C(n_343),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_315),
.B(n_286),
.C(n_298),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_281),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_304),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_330),
.C(n_321),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_307),
.B(n_284),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_SL g355 ( 
.A(n_344),
.B(n_319),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_351),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_329),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_311),
.A2(n_240),
.B1(n_266),
.B2(n_300),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_350),
.A2(n_325),
.B1(n_312),
.B2(n_317),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_327),
.B(n_259),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_313),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_354),
.A2(n_357),
.B(n_332),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_355),
.B(n_368),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_309),
.Y(n_356)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

NAND5xp2_ASAP7_75t_SL g357 ( 
.A(n_344),
.B(n_324),
.C(n_343),
.D(n_335),
.E(n_339),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_334),
.Y(n_358)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_349),
.A2(n_346),
.B1(n_342),
.B2(n_324),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_360),
.A2(n_350),
.B1(n_332),
.B2(n_328),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_333),
.Y(n_362)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_362),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_322),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_363),
.B(n_367),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_331),
.B(n_325),
.C(n_314),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_365),
.C(n_369),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_340),
.C(n_337),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_366),
.A2(n_326),
.B1(n_323),
.B2(n_313),
.Y(n_374)
);

BUFx12_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_306),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_345),
.C(n_348),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_370),
.B(n_352),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_371),
.A2(n_357),
.B1(n_353),
.B2(n_359),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_374),
.A2(n_383),
.B1(n_382),
.B2(n_372),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_323),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_378),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_376),
.B(n_352),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_361),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_310),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_381),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_369),
.B(n_310),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_389),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_386),
.B(n_388),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_291),
.C(n_301),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_367),
.B(n_299),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_374),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_367),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_380),
.C(n_381),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_292),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_393),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_394),
.B(n_257),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_379),
.C(n_375),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_392),
.C(n_385),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_376),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_400),
.B(n_288),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_392),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_401),
.B(n_402),
.Y(n_406)
);

OAI21x1_ASAP7_75t_SL g407 ( 
.A1(n_404),
.A2(n_398),
.B(n_357),
.Y(n_407)
);

AOI322xp5_ASAP7_75t_L g405 ( 
.A1(n_403),
.A2(n_399),
.A3(n_398),
.B1(n_397),
.B2(n_262),
.C1(n_258),
.C2(n_231),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_405),
.B(n_407),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_406),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_408),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_410),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_411),
.Y(n_412)
);


endmodule