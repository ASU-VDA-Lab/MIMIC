module fake_jpeg_27120_n_87 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_87);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_0),
.B(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_20),
.B1(n_18),
.B2(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_2),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_13),
.Y(n_37)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_19),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_15),
.B(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_21),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_3),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_20),
.B(n_17),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_35),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_36),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_22),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_27),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_45),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_28),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_64),
.B1(n_30),
.B2(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_52),
.B(n_47),
.Y(n_59)
);

AO21x1_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_60),
.B(n_25),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_43),
.B1(n_46),
.B2(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_65),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OAI221xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_68),
.B1(n_73),
.B2(n_59),
.C(n_61),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_48),
.B(n_49),
.C(n_30),
.D(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_73),
.A3(n_69),
.B1(n_26),
.B2(n_18),
.C(n_9),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_77),
.B(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_18),
.B1(n_11),
.B2(n_17),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_14),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

OAI322xp33_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_79),
.A3(n_9),
.B1(n_10),
.B2(n_16),
.C1(n_5),
.C2(n_6),
.Y(n_86)
);

AOI221xp5_ASAP7_75t_L g87 ( 
.A1(n_86),
.A2(n_7),
.B1(n_84),
.B2(n_83),
.C(n_81),
.Y(n_87)
);


endmodule