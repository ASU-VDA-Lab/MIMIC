module fake_jpeg_10625_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_33),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_19),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_22),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_32),
.B1(n_21),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_55),
.B1(n_56),
.B2(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_32),
.B1(n_19),
.B2(n_30),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_32),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_16),
.B1(n_22),
.B2(n_28),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_27),
.B1(n_34),
.B2(n_28),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_17),
.B1(n_24),
.B2(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_16),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_68),
.Y(n_71)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_35),
.A2(n_34),
.B1(n_30),
.B2(n_27),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_20),
.B1(n_38),
.B2(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_66),
.B(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_21),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_70),
.B(n_88),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_83),
.B(n_87),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_82),
.B(n_93),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_43),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_18),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_29),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_38),
.B1(n_49),
.B2(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_94),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_48),
.B(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_46),
.B(n_51),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_29),
.Y(n_97)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_75),
.B(n_23),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_40),
.B(n_23),
.Y(n_143)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_79),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_49),
.B1(n_38),
.B2(n_58),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_72),
.B1(n_41),
.B2(n_24),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_52),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_122),
.C(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_121),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_63),
.B1(n_59),
.B2(n_38),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_81),
.B1(n_96),
.B2(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_52),
.C(n_59),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_96),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_135),
.B1(n_138),
.B2(n_151),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_112),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_133),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_93),
.B(n_74),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_144),
.B(n_145),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_90),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_102),
.A2(n_73),
.B1(n_76),
.B2(n_84),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_0),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_150),
.Y(n_177)
);

INVxp33_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_140),
.B1(n_104),
.B2(n_124),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_102),
.A2(n_73),
.B1(n_84),
.B2(n_41),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_78),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_149),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_23),
.A3(n_26),
.B1(n_33),
.B2(n_24),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_113),
.B1(n_155),
.B2(n_106),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_147),
.B(n_100),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_119),
.B(n_108),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_0),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_23),
.B(n_26),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_152),
.C(n_124),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_108),
.B(n_72),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_41),
.B1(n_51),
.B2(n_67),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_85),
.C(n_40),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_85),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_29),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_120),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_0),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_169),
.B(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_164),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_172),
.B1(n_173),
.B2(n_179),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_103),
.B(n_98),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_152),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_171),
.B(n_175),
.C(n_178),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_109),
.B1(n_107),
.B2(n_99),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_131),
.B(n_125),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_51),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_189),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_105),
.B1(n_12),
.B2(n_13),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_40),
.C(n_67),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_143),
.C(n_132),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_126),
.A2(n_40),
.B1(n_26),
.B2(n_23),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_181),
.A2(n_154),
.B1(n_128),
.B2(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_127),
.B(n_29),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_183),
.Y(n_193)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_29),
.Y(n_185)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_135),
.A2(n_40),
.B1(n_26),
.B2(n_23),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_186),
.B1(n_142),
.B2(n_190),
.Y(n_206)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_130),
.B(n_18),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_144),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_190),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_188),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_195),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_199),
.B(n_157),
.Y(n_225)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_177),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_203),
.A2(n_219),
.B1(n_173),
.B2(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_129),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_205),
.B(n_210),
.C(n_214),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_206),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_215),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_145),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_146),
.B1(n_141),
.B2(n_132),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_213),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_167),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_146),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_163),
.B(n_177),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_160),
.A2(n_168),
.B1(n_169),
.B2(n_176),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_178),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_227),
.C(n_241),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_221),
.B(n_222),
.Y(n_260)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_217),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_234),
.Y(n_259)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_161),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_163),
.B1(n_169),
.B2(n_161),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_229),
.A2(n_194),
.B1(n_208),
.B2(n_212),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_237),
.B1(n_238),
.B2(n_240),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_193),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_233),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_170),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx8_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_192),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_180),
.C(n_170),
.Y(n_241)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_242),
.A2(n_199),
.B1(n_195),
.B2(n_216),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_189),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_214),
.C(n_198),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_250),
.C(n_254),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_245),
.B1(n_236),
.B2(n_229),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_238),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_198),
.C(n_218),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_197),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_218),
.C(n_202),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_262),
.C(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_261),
.A2(n_228),
.B1(n_235),
.B2(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_145),
.C(n_204),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_145),
.C(n_140),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_225),
.B(n_136),
.C(n_18),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_1),
.C(n_2),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_265),
.A2(n_242),
.B(n_224),
.Y(n_270)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_276),
.B1(n_278),
.B2(n_281),
.Y(n_286)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_240),
.B(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_258),
.A2(n_226),
.B1(n_136),
.B2(n_3),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_258),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_4),
.B1(n_26),
.B2(n_6),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_264),
.C(n_262),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_248),
.A2(n_1),
.B(n_2),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_263),
.Y(n_291)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_290),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_269),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_246),
.C(n_256),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_297),
.C(n_276),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_289),
.A2(n_4),
.B1(n_26),
.B2(n_7),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_274),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_291),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_259),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_294),
.B(n_295),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_250),
.C(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_247),
.C(n_259),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_275),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_305),
.Y(n_313)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_301),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_277),
.B1(n_282),
.B2(n_267),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_307),
.B1(n_291),
.B2(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_278),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_306),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_296),
.A2(n_280),
.B(n_5),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_9),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_8),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_9),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_303),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_11),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_317),
.A2(n_288),
.B(n_299),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_287),
.B(n_285),
.Y(n_318)
);

AOI211xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_310),
.B(n_300),
.C(n_33),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_9),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_317),
.B(n_313),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_18),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_330),
.A2(n_321),
.B(n_322),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_328),
.A3(n_326),
.B1(n_13),
.B2(n_14),
.C1(n_12),
.C2(n_11),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_332),
.B(n_13),
.CI(n_324),
.CON(n_333),
.SN(n_333)
);


endmodule