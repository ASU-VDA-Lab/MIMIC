module real_jpeg_14357_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_3),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_3),
.A2(n_33),
.B1(n_36),
.B2(n_57),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_3),
.A2(n_57),
.B1(n_77),
.B2(n_78),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_82),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_82),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_82),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_5),
.A2(n_77),
.B1(n_78),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_5),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_5),
.A2(n_74),
.B(n_77),
.C(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_5),
.B(n_84),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_5),
.B(n_63),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_SL g214 ( 
.A1(n_5),
.A2(n_63),
.B(n_200),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_33),
.C(n_51),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_144),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_5),
.B(n_90),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_48),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_48),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_9),
.A2(n_48),
.B1(n_77),
.B2(n_78),
.Y(n_290)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_77),
.B1(n_78),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_147),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_147),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_11),
.A2(n_33),
.B1(n_36),
.B2(n_147),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_13),
.A2(n_77),
.B1(n_78),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_13),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_135),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_13),
.A2(n_33),
.B1(n_36),
.B2(n_135),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_14),
.A2(n_35),
.B1(n_77),
.B2(n_78),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_14),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_14),
.A2(n_35),
.B1(n_63),
.B2(n_64),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_15),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_15),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_15),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_15),
.A2(n_41),
.B1(n_77),
.B2(n_78),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_321),
.C(n_325),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_319),
.B(n_323),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_312),
.B(n_318),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_278),
.B(n_309),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_136),
.B(n_277),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_114),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_22),
.B(n_114),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_86),
.B2(n_113),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_23),
.B(n_87),
.C(n_98),
.Y(n_307)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_58),
.C(n_71),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_25),
.A2(n_26),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_27),
.A2(n_28),
.B1(n_42),
.B2(n_43),
.Y(n_266)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_30),
.A2(n_38),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_31),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_31),
.A2(n_124),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_31),
.A2(n_37),
.B(n_162),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_31),
.A2(n_161),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_32),
.A2(n_126),
.B(n_161),
.Y(n_203)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_54)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_36),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_38),
.A2(n_39),
.B(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_38),
.A2(n_123),
.B(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_38),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_38),
.A2(n_39),
.B1(n_229),
.B2(n_237),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_39),
.B(n_40),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_39),
.B(n_144),
.Y(n_235)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_45),
.A2(n_54),
.B(n_95),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_SL g201 ( 
.A(n_46),
.B(n_60),
.C(n_64),
.Y(n_201)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_47),
.A2(n_61),
.B(n_199),
.C(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_47),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_56),
.B(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_49),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_49),
.A2(n_55),
.B1(n_195),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_49),
.A2(n_55),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_49),
.A2(n_55),
.B1(n_216),
.B2(n_226),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_54),
.B(n_144),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_54),
.A2(n_154),
.B(n_155),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_96),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_58),
.B(n_71),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_66),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_59),
.B(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_59),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_59),
.A2(n_68),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_59),
.A2(n_68),
.B1(n_150),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_59),
.A2(n_68),
.B1(n_172),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_69)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_64),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_63),
.A2(n_75),
.B(n_144),
.Y(n_165)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_66),
.B(n_178),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_67),
.A2(n_90),
.B(n_179),
.Y(n_315)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_68),
.A2(n_151),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_68),
.A2(n_131),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_70),
.B(n_90),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_81),
.B(n_83),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_72),
.A2(n_110),
.B(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_73),
.B1(n_81),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_72),
.A2(n_73),
.B1(n_134),
.B2(n_146),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_72),
.A2(n_73),
.B1(n_290),
.B2(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_72),
.A2(n_111),
.B(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_73),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_83),
.B(n_291),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_84),
.A2(n_85),
.B(n_142),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_98),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B(n_97),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_90),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_91),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_93),
.A2(n_154),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_97),
.B(n_281),
.C(n_293),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_97),
.B(n_281),
.CI(n_293),
.CON(n_308),
.SN(n_308)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g293 ( 
.A1(n_99),
.A2(n_100),
.B(n_108),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_100),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_102),
.B1(n_103),
.B2(n_107),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_105),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_112),
.B(n_142),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_119),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_120),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.C(n_132),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_121),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_127),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_128),
.A2(n_129),
.B1(n_132),
.B2(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_271),
.B(n_276),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_184),
.B(n_262),
.C(n_270),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_173),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_139),
.B(n_173),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_157),
.C(n_166),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_152),
.C(n_156),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_152),
.B1(n_153),
.B2(n_156),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_158),
.B1(n_166),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_163),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_174),
.B(n_182),
.C(n_183),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_176),
.B(n_177),
.C(n_180),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_260),
.B(n_261),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_204),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_190),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_187),
.B(n_190),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_196),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_193),
.A2(n_196),
.B1(n_197),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_202),
.B1(n_203),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_217),
.B(n_259),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_206),
.B(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_215),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_253),
.B(n_258),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_243),
.B(n_252),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_232),
.B(n_242),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_227),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_224),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_241),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_245),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_248),
.C(n_251),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_266),
.C(n_267),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_306),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_279),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_294),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_294),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_289),
.B2(n_292),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_288),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_288),
.C(n_289),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_288),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_301),
.C(n_303),
.Y(n_317)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_292),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_295),
.C(n_298),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_308),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_314),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_321),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.CI(n_317),
.CON(n_314),
.SN(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_322),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);


endmodule