module fake_netlist_6_2731_n_662 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_662);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_662;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_229;
wire n_542;
wire n_644;
wire n_621;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_659;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_624;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_550;
wire n_487;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_612;
wire n_633;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_655;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_26),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_71),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_49),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_11),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_4),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_19),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_51),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_53),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_138),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_41),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_8),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_46),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_81),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_2),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_70),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_43),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_0),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_91),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_60),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_39),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_23),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_17),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_140),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_95),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_136),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_74),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_54),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_68),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_48),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_69),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_143),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_44),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_13),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_64),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_85),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_103),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_80),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_57),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_21),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_67),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_79),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_31),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_1),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_110),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_105),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_20),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_0),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

XNOR2x2_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_1),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_2),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_175),
.Y(n_221)
);

AND2x4_ASAP7_75t_SL g222 ( 
.A(n_213),
.B(n_15),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_3),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_154),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_16),
.Y(n_225)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_149),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_150),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_3),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_175),
.B(n_4),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_5),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_5),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_173),
.B(n_6),
.Y(n_237)
);

AND2x6_ASAP7_75t_L g238 ( 
.A(n_148),
.B(n_18),
.Y(n_238)
);

BUFx8_ASAP7_75t_SL g239 ( 
.A(n_188),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_188),
.B(n_6),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_175),
.B(n_7),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_175),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_156),
.B(n_9),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_9),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_155),
.B(n_162),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_171),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_145),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_196),
.B(n_10),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_10),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_12),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_12),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_146),
.B(n_14),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_186),
.B(n_14),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_22),
.Y(n_258)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_147),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_153),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_24),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_157),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_202),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_266)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_151),
.B1(n_168),
.B2(n_206),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

AO22x2_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_214),
.B1(n_212),
.B2(n_210),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_226),
.B(n_158),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_159),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

AO22x2_ASAP7_75t_L g276 ( 
.A1(n_256),
.A2(n_209),
.B1(n_200),
.B2(n_199),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_197),
.B1(n_194),
.B2(n_193),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_224),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_229),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_160),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_230),
.B(n_163),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_243),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_166),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_226),
.B(n_167),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_235),
.A2(n_181),
.B1(n_190),
.B2(n_185),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_223),
.A2(n_191),
.B1(n_183),
.B2(n_178),
.Y(n_286)
);

OR2x6_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_169),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_172),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_236),
.A2(n_177),
.B1(n_27),
.B2(n_28),
.Y(n_289)
);

CKINVDCx6p67_ASAP7_75t_R g290 ( 
.A(n_226),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_236),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_252),
.A2(n_234),
.B1(n_253),
.B2(n_227),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_32),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_33),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g296 ( 
.A1(n_215),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

AND2x6_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_225),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

BUFx6f_ASAP7_75t_SL g300 ( 
.A(n_245),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_252),
.A2(n_246),
.B1(n_245),
.B2(n_222),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_231),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_254),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

OAI22xp33_ASAP7_75t_L g306 ( 
.A1(n_255),
.A2(n_50),
.B1(n_52),
.B2(n_55),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_257),
.A2(n_242),
.B1(n_232),
.B2(n_233),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g308 ( 
.A1(n_218),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_261),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_65),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_251),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_218),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

OAI22xp33_ASAP7_75t_L g314 ( 
.A1(n_233),
.A2(n_75),
.B1(n_77),
.B2(n_82),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_274),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_279),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_222),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_262),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_267),
.B(n_217),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_307),
.A2(n_238),
.B(n_241),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_259),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_298),
.B(n_219),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_260),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_239),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_269),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_285),
.B(n_260),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_R g334 ( 
.A(n_287),
.B(n_239),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_260),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_273),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_259),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_278),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_270),
.B(n_86),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_301),
.B(n_260),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_266),
.B(n_259),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_251),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_272),
.B(n_221),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_241),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_287),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_292),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_311),
.Y(n_352)
);

NAND2x1p5_ASAP7_75t_L g353 ( 
.A(n_291),
.B(n_244),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_270),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_280),
.B(n_244),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_276),
.B(n_87),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_281),
.B(n_238),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_276),
.B(n_244),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_291),
.B(n_244),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_310),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_300),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_294),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_277),
.B(n_89),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_302),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_298),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_298),
.A2(n_238),
.B(n_92),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_271),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_284),
.B(n_238),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_289),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

NAND2x1p5_ASAP7_75t_L g380 ( 
.A(n_303),
.B(n_238),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_312),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_330),
.B(n_90),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_320),
.B(n_94),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_320),
.B(n_96),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_349),
.B(n_97),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_98),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_321),
.B(n_100),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_335),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_350),
.B(n_101),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_345),
.B(n_314),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_363),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_309),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_322),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_102),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_316),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_317),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_104),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_357),
.Y(n_404)
);

OR2x2_ASAP7_75t_L g405 ( 
.A(n_372),
.B(n_296),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_378),
.B(n_306),
.Y(n_406)
);

AND2x4_ASAP7_75t_SL g407 ( 
.A(n_367),
.B(n_108),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_362),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_324),
.B(n_109),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_324),
.B(n_111),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_364),
.B(n_112),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_347),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_144),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_382),
.B(n_115),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_347),
.A2(n_377),
.B(n_327),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_339),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_116),
.Y(n_419)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_374),
.A2(n_327),
.B(n_342),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_319),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

AND2x4_ASAP7_75t_SL g424 ( 
.A(n_348),
.B(n_375),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_315),
.B(n_120),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_344),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_353),
.B(n_121),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_353),
.B(n_122),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_123),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_124),
.Y(n_430)
);

AND2x6_ASAP7_75t_L g431 ( 
.A(n_333),
.B(n_125),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_323),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_361),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_340),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_319),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_365),
.B(n_126),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_325),
.B(n_127),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_380),
.B(n_132),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_326),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_380),
.B(n_133),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_331),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_337),
.B(n_135),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_336),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_374),
.A2(n_137),
.B(n_141),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_338),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_343),
.B(n_318),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_332),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_370),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_341),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_359),
.Y(n_450)
);

NAND2x1p5_ASAP7_75t_L g451 ( 
.A(n_392),
.B(n_346),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_409),
.B(n_351),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_394),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_434),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_444),
.B(n_328),
.Y(n_456)
);

AO21x2_ASAP7_75t_L g457 ( 
.A1(n_417),
.A2(n_352),
.B(n_329),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_434),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_392),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_394),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_392),
.Y(n_461)
);

BUFx4f_ASAP7_75t_L g462 ( 
.A(n_429),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_142),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_426),
.B(n_334),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g467 ( 
.A(n_383),
.Y(n_467)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_406),
.B(n_396),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_420),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_410),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_446),
.B(n_439),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_392),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_397),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

OR2x6_ASAP7_75t_L g482 ( 
.A(n_429),
.B(n_413),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_416),
.B(n_403),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_448),
.B(n_405),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_424),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_403),
.B(n_390),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_416),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_413),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_416),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_409),
.B(n_410),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_406),
.B(n_420),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_489),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_466),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_455),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_472),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_388),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_492),
.Y(n_501)
);

OR2x6_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_413),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_476),
.Y(n_503)
);

BUFx12f_ASAP7_75t_L g504 ( 
.A(n_485),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_432),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_458),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_474),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_476),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_476),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_468),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_489),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_431),
.B1(n_442),
.B2(n_414),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_488),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g514 ( 
.A(n_488),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_477),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_476),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_388),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

BUFx12f_ASAP7_75t_L g519 ( 
.A(n_465),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_470),
.B(n_414),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_481),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_459),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_482),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_494),
.Y(n_524)
);

BUFx8_ASAP7_75t_L g525 ( 
.A(n_506),
.Y(n_525)
);

INVx11_ASAP7_75t_L g526 ( 
.A(n_519),
.Y(n_526)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_504),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_508),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_500),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_520),
.A2(n_491),
.B1(n_469),
.B2(n_456),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_520),
.A2(n_491),
.B1(n_456),
.B2(n_490),
.Y(n_533)
);

BUFx2_ASAP7_75t_R g534 ( 
.A(n_496),
.Y(n_534)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_519),
.Y(n_535)
);

CKINVDCx6p67_ASAP7_75t_R g536 ( 
.A(n_506),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_512),
.A2(n_490),
.B1(n_431),
.B2(n_486),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_505),
.A2(n_431),
.B1(n_442),
.B2(n_405),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_496),
.Y(n_539)
);

CKINVDCx11_ASAP7_75t_R g540 ( 
.A(n_504),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_494),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_495),
.B(n_480),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

BUFx12f_ASAP7_75t_L g544 ( 
.A(n_499),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_497),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_510),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_501),
.Y(n_548)
);

CKINVDCx11_ASAP7_75t_R g549 ( 
.A(n_510),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_500),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_525),
.A2(n_462),
.B1(n_418),
.B2(n_431),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_538),
.A2(n_457),
.B1(n_431),
.B2(n_462),
.Y(n_552)
);

BUFx4f_ASAP7_75t_SL g553 ( 
.A(n_544),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_542),
.A2(n_464),
.B1(n_457),
.B2(n_471),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_538),
.A2(n_431),
.B1(n_467),
.B2(n_479),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_524),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_539),
.A2(n_471),
.B1(n_408),
.B2(n_482),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_532),
.A2(n_431),
.B1(n_523),
.B2(n_498),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_532),
.A2(n_523),
.B1(n_498),
.B2(n_390),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_537),
.A2(n_502),
.B1(n_484),
.B2(n_473),
.Y(n_560)
);

OAI21xp33_ASAP7_75t_L g561 ( 
.A1(n_533),
.A2(n_391),
.B(n_395),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_541),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_537),
.A2(n_502),
.B1(n_483),
.B2(n_473),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_528),
.B(n_475),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_475),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_549),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_545),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_533),
.A2(n_498),
.B1(n_517),
.B2(n_502),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_536),
.A2(n_498),
.B1(n_517),
.B2(n_424),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_535),
.A2(n_517),
.B1(n_502),
.B2(n_463),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_530),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_550),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_547),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_574)
);

AND2x4_ASAP7_75t_SL g575 ( 
.A(n_529),
.B(n_508),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_525),
.A2(n_430),
.B1(n_440),
.B2(n_438),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_528),
.Y(n_577)
);

AOI222xp33_ASAP7_75t_L g578 ( 
.A1(n_540),
.A2(n_413),
.B1(n_430),
.B2(n_440),
.C1(n_438),
.C2(n_384),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_547),
.B(n_463),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_535),
.A2(n_407),
.B1(n_453),
.B2(n_411),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_535),
.A2(n_411),
.B1(n_478),
.B2(n_387),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_578),
.A2(n_453),
.B1(n_527),
.B2(n_540),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_578),
.A2(n_453),
.B1(n_402),
.B2(n_436),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_577),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_561),
.A2(n_453),
.B1(n_428),
.B2(n_427),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_574),
.A2(n_407),
.B1(n_386),
.B2(n_387),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_554),
.B(n_501),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_560),
.A2(n_443),
.B1(n_445),
.B2(n_421),
.Y(n_588)
);

OAI221xp5_ASAP7_75t_L g589 ( 
.A1(n_576),
.A2(n_437),
.B1(n_514),
.B2(n_513),
.C(n_433),
.Y(n_589)
);

OAI21xp33_ASAP7_75t_L g590 ( 
.A1(n_552),
.A2(n_565),
.B(n_581),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_560),
.A2(n_443),
.B1(n_445),
.B2(n_421),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_557),
.A2(n_534),
.B1(n_547),
.B2(n_526),
.Y(n_592)
);

OAI221xp5_ASAP7_75t_L g593 ( 
.A1(n_570),
.A2(n_433),
.B1(n_423),
.B2(n_441),
.C(n_518),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_568),
.A2(n_423),
.B1(n_441),
.B2(n_385),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_SL g595 ( 
.A1(n_563),
.A2(n_516),
.B1(n_518),
.B2(n_531),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_566),
.A2(n_516),
.B1(n_531),
.B2(n_546),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_559),
.A2(n_551),
.B1(n_558),
.B2(n_555),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_580),
.A2(n_450),
.B1(n_419),
.B2(n_449),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_556),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_572),
.B(n_507),
.Y(n_600)
);

OAI222xp33_ASAP7_75t_L g601 ( 
.A1(n_569),
.A2(n_515),
.B1(n_507),
.B2(n_522),
.C1(n_521),
.C2(n_450),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_562),
.B(n_515),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_567),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_571),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_564),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_599),
.B(n_573),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_599),
.B(n_579),
.Y(n_607)
);

AOI21x1_ASAP7_75t_L g608 ( 
.A1(n_587),
.A2(n_449),
.B(n_425),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_604),
.B(n_566),
.Y(n_609)
);

OAI221xp5_ASAP7_75t_L g610 ( 
.A1(n_582),
.A2(n_566),
.B1(n_521),
.B2(n_511),
.C(n_522),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_589),
.B(n_549),
.C(n_493),
.Y(n_611)
);

AO22x1_ASAP7_75t_L g612 ( 
.A1(n_592),
.A2(n_553),
.B1(n_546),
.B2(n_529),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_584),
.B(n_575),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_604),
.B(n_546),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_602),
.B(n_546),
.Y(n_615)
);

OA21x2_ASAP7_75t_L g616 ( 
.A1(n_601),
.A2(n_400),
.B(n_404),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_586),
.B(n_531),
.C(n_529),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_531),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_595),
.B(n_529),
.Y(n_619)
);

NAND4xp75_ASAP7_75t_L g620 ( 
.A(n_619),
.B(n_600),
.C(n_596),
.D(n_511),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_617),
.A2(n_597),
.B1(n_583),
.B2(n_593),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_607),
.B(n_590),
.Y(n_622)
);

NAND4xp75_ASAP7_75t_L g623 ( 
.A(n_609),
.B(n_400),
.C(n_404),
.D(n_598),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_611),
.B(n_591),
.C(n_588),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_594),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_585),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_618),
.B(n_493),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_627),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_622),
.B(n_610),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_627),
.Y(n_630)
);

NAND4xp75_ASAP7_75t_L g631 ( 
.A(n_626),
.B(n_614),
.C(n_606),
.D(n_616),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_625),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_620),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_623),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_628),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_633),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_632),
.B(n_612),
.Y(n_637)
);

NOR2x1_ASAP7_75t_R g638 ( 
.A(n_634),
.B(n_503),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_630),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_635),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_636),
.B(n_629),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_636),
.A2(n_621),
.B1(n_631),
.B2(n_624),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_639),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_637),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_643),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_640),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_644),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_647),
.Y(n_648)
);

OA22x2_ASAP7_75t_L g649 ( 
.A1(n_645),
.A2(n_642),
.B1(n_641),
.B2(n_638),
.Y(n_649)
);

OAI211xp5_ASAP7_75t_L g650 ( 
.A1(n_648),
.A2(n_646),
.B(n_617),
.C(n_615),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_650),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_651),
.Y(n_652)
);

AO22x1_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_649),
.B1(n_493),
.B2(n_508),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_608),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_654),
.A2(n_616),
.B1(n_509),
.B2(n_503),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_655),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_656),
.A2(n_509),
.B1(n_503),
.B2(n_489),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_657),
.Y(n_658)
);

AO22x2_ASAP7_75t_L g659 ( 
.A1(n_658),
.A2(n_509),
.B1(n_487),
.B2(n_461),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_659),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g661 ( 
.A1(n_660),
.A2(n_422),
.B1(n_393),
.B2(n_435),
.C(n_451),
.Y(n_661)
);

AOI211xp5_ASAP7_75t_L g662 ( 
.A1(n_661),
.A2(n_447),
.B(n_451),
.C(n_393),
.Y(n_662)
);


endmodule