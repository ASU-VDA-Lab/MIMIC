module real_jpeg_20595_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_346, n_347, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_346;
input n_347;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_0),
.A2(n_24),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_0),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_0),
.A2(n_35),
.B1(n_71),
.B2(n_72),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_1),
.A2(n_24),
.B1(n_26),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_1),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_1),
.A2(n_71),
.B1(n_72),
.B2(n_95),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_95),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_71),
.B1(n_72),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_2),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_131),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_131),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_2),
.A2(n_24),
.B1(n_26),
.B2(n_131),
.Y(n_268)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_4),
.A2(n_24),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_62),
.B1(n_71),
.B2(n_72),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_4),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_62),
.Y(n_284)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_55),
.B(n_67),
.C(n_111),
.D(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_5),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_5),
.B(n_53),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_5),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_132),
.B(n_134),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_5),
.A2(n_32),
.B(n_48),
.C(n_171),
.D(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_5),
.B(n_32),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_5),
.B(n_36),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_5),
.A2(n_24),
.B1(n_26),
.B2(n_155),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_5),
.A2(n_33),
.B(n_224),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_24),
.B1(n_26),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_6),
.A2(n_64),
.B1(n_71),
.B2(n_72),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_6),
.A2(n_54),
.B1(n_55),
.B2(n_64),
.Y(n_259)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_7),
.Y(n_133)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_7),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_7),
.A2(n_153),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_144),
.B1(n_181),
.B2(n_196),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_9),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_9),
.A2(n_71),
.B1(n_72),
.B2(n_114),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_114),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_9),
.A2(n_24),
.B1(n_26),
.B2(n_114),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_11),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_71),
.B1(n_72),
.B2(n_126),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_126),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_11),
.A2(n_24),
.B1(n_26),
.B2(n_126),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_12),
.A2(n_23),
.B1(n_32),
.B2(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_12),
.A2(n_23),
.B1(n_71),
.B2(n_72),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_12),
.A2(n_23),
.B1(n_54),
.B2(n_55),
.Y(n_291)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_38),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_21),
.B(n_42),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_34),
.B2(n_36),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_22),
.A2(n_27),
.B1(n_36),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_24),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_29),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_24),
.A2(n_29),
.B(n_155),
.C(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_34),
.B(n_36),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_27),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_28),
.A2(n_31),
.B1(n_239),
.B2(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_28),
.A2(n_217),
.B(n_268),
.Y(n_286)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_29),
.Y(n_224)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_31),
.A2(n_239),
.B(n_240),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_31),
.A2(n_94),
.B(n_240),
.Y(n_310)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_52),
.C(n_53),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_36),
.B(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

OAI21x1_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_81),
.B(n_344),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_76),
.C(n_78),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_44),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_59),
.C(n_65),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_46),
.B1(n_65),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_56),
.B1(n_57),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_47),
.A2(n_57),
.B1(n_190),
.B2(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_47),
.A2(n_212),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_53),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_48),
.B(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_48),
.A2(n_53),
.B1(n_265),
.B2(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_48),
.A2(n_53),
.B1(n_100),
.B2(n_284),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_49),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_50),
.B(n_54),
.Y(n_178)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_52),
.Y(n_179)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_68),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_55),
.A2(n_171),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_57),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_57),
.A2(n_190),
.B(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_57),
.A2(n_191),
.B(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_60),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_65),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B(n_75),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_66),
.A2(n_74),
.B1(n_125),
.B2(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_66),
.A2(n_169),
.B(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_66),
.A2(n_74),
.B1(n_209),
.B2(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_66),
.A2(n_74),
.B1(n_250),
.B2(n_259),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_66),
.A2(n_74),
.B1(n_259),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_67),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_67),
.A2(n_70),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_68),
.B(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_71),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_71),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_72),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_74),
.B(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_74),
.A2(n_127),
.B(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_75),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21x1_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_101),
.B(n_343),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_83),
.B(n_87),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.C(n_96),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_329),
.Y(n_335)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_93),
.C(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_93),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_93),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_96),
.B(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

OAI321xp33_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_326),
.A3(n_336),
.B1(n_341),
.B2(n_342),
.C(n_346),
.Y(n_101)
);

AOI321xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_276),
.A3(n_314),
.B1(n_320),
.B2(n_325),
.C(n_347),
.Y(n_102)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_233),
.C(n_272),
.Y(n_103)
);

AOI21x1_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_203),
.B(n_232),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_184),
.B(n_202),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_163),
.B(n_183),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_139),
.B(n_162),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_109),
.B(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_115),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_115),
.B1(n_116),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_129),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_124),
.C(n_129),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_132),
.B(n_134),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_136),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_132),
.A2(n_151),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_132),
.A2(n_151),
.B1(n_228),
.B2(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_132),
.A2(n_133),
.B1(n_248),
.B2(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_132),
.A2(n_133),
.B(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_148),
.B(n_161),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_146),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_151),
.B(n_152),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_156),
.B(n_160),
.Y(n_148)
);

NOR2xp67_ASAP7_75t_R g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_155),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_164),
.B(n_165),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_176),
.B2(n_182),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_175),
.C(n_182),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_172),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_173),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_185),
.B(n_186),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_198),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_199),
.C(n_200),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_197),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_194),
.C(n_195),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_205),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_220),
.C(n_231),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_213),
.C(n_214),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_225),
.B2(n_226),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_226),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_234),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_252),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_235),
.B(n_252),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_246),
.C(n_251),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_236),
.B(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_245),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_270)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_251),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_249),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_270),
.B2(n_271),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_255),
.B(n_260),
.C(n_271),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_258),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_266),
.C(n_269),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_263),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_274),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_294),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_277),
.B(n_294),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.C(n_293),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_278),
.A2(n_279),
.B1(n_287),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_283),
.C(n_285),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_292),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_288),
.A2(n_289),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_288),
.A2(n_306),
.B(n_310),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_290),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_290),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_291),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_312),
.B2(n_313),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_304),
.B2(n_305),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_305),
.C(n_313),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_302),
.B(n_303),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_302),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_303),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_303),
.A2(n_328),
.B1(n_332),
.B2(n_340),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_308),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_312),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_315),
.A2(n_321),
.B(n_324),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_316),
.B(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_334),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_334),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.C(n_333),
.Y(n_327)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_328),
.Y(n_340)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);


endmodule