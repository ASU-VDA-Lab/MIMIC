module fake_jpeg_8973_n_175 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_53),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_32),
.A2(n_19),
.B1(n_18),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_24),
.C(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_16),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_25),
.C(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_41),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_27),
.B1(n_19),
.B2(n_31),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_41),
.B1(n_15),
.B2(n_26),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_74),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_68),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_42),
.B1(n_40),
.B2(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_48),
.B(n_60),
.C(n_46),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_38),
.B1(n_31),
.B2(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_24),
.B1(n_15),
.B2(n_23),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_29),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_79),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_28),
.B1(n_20),
.B2(n_41),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_21),
.B1(n_36),
.B2(n_28),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_43),
.B(n_47),
.C(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_48),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_70),
.C(n_72),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_50),
.B(n_60),
.C(n_36),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_78),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_112),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_74),
.C(n_67),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_113),
.Y(n_129)
);

INVxp33_ASAP7_75t_SL g107 ( 
.A(n_95),
.Y(n_107)
);

OAI22x1_ASAP7_75t_L g122 ( 
.A1(n_107),
.A2(n_110),
.B1(n_83),
.B2(n_80),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_68),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_86),
.B1(n_87),
.B2(n_97),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_118),
.B1(n_99),
.B2(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_86),
.B1(n_87),
.B2(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_125),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_123),
.B1(n_102),
.B2(n_108),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_112),
.A2(n_93),
.B1(n_88),
.B2(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_104),
.B(n_89),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_135),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_122),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_136),
.B(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_141),
.B1(n_115),
.B2(n_77),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_92),
.C(n_90),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_116),
.C(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_22),
.B(n_1),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_128),
.B(n_115),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_141),
.B1(n_133),
.B2(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_100),
.B1(n_91),
.B2(n_55),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_147),
.A2(n_150),
.B1(n_96),
.B2(n_22),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_100),
.B1(n_91),
.B2(n_79),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_153),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_149),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_155),
.C(n_150),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_147),
.C(n_146),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_152),
.B1(n_155),
.B2(n_154),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_2),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_144),
.B(n_145),
.C(n_148),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_163),
.B1(n_8),
.B2(n_9),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_162),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_158),
.A2(n_142),
.B1(n_1),
.B2(n_2),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_161),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_168),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_165),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_166),
.A2(n_159),
.B(n_160),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_161),
.B(n_10),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.C(n_14),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.C(n_5),
.Y(n_175)
);


endmodule