module fake_netlist_6_681_n_892 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_892);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_892;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_465;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_248;
wire n_222;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_544;
wire n_468;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_608;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_474;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_598;
wire n_496;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_663;
wire n_508;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_8),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_51),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_44),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_74),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_111),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_154),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_189),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_115),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_179),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_85),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_16),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_66),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_75),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_40),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_170),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_175),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_52),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_100),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_73),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_168),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_6),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_5),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_19),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_120),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_156),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_104),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_160),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_148),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_64),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_7),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_108),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_173),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_101),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_48),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_15),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_33),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_177),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_176),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_71),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_63),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_87),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_78),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_178),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

INVx4_ASAP7_75t_R g249 ( 
.A(n_172),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_103),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_35),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_20),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_180),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_159),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_76),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_188),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_18),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_136),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_144),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_162),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_118),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_130),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_164),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_132),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_0),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_200),
.B(n_0),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_200),
.B(n_29),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_30),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_202),
.B(n_1),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_228),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_193),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_1),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_195),
.B(n_2),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_197),
.B(n_2),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_199),
.Y(n_288)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_242),
.B(n_3),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_204),
.B(n_3),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_206),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_208),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_194),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_198),
.B(n_4),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_212),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_237),
.B(n_4),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_220),
.B(n_5),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_6),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_215),
.Y(n_303)
);

BUFx8_ASAP7_75t_SL g304 ( 
.A(n_209),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_223),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_214),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_216),
.B(n_7),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_232),
.B(n_8),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_31),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_231),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_194),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_9),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

BUFx12f_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_10),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_234),
.B(n_10),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_251),
.B(n_32),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_261),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_263),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_278),
.A2(n_209),
.B1(n_244),
.B2(n_257),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

NAND3x1_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_265),
.C(n_11),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_283),
.A2(n_244),
.B1(n_257),
.B2(n_230),
.Y(n_327)
);

AO22x2_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_L g331 ( 
.A1(n_289),
.A2(n_269),
.B1(n_196),
.B2(n_230),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_269),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_271),
.A2(n_268),
.B1(n_267),
.B2(n_264),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_319),
.B1(n_301),
.B2(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_276),
.A2(n_262),
.B1(n_260),
.B2(n_258),
.Y(n_336)
);

AO22x2_ASAP7_75t_L g337 ( 
.A1(n_275),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_279),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g339 ( 
.A1(n_276),
.A2(n_256),
.B1(n_252),
.B2(n_250),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_297),
.A2(n_247),
.B1(n_246),
.B2(n_245),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_241),
.B1(n_240),
.B2(n_238),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_217),
.B1(n_235),
.B2(n_227),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

AO22x2_ASAP7_75t_L g346 ( 
.A1(n_275),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_300),
.B(n_192),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_R g348 ( 
.A1(n_303),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_348)
);

OR2x6_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_17),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_201),
.Y(n_350)
);

BUFx6f_ASAP7_75t_SL g351 ( 
.A(n_275),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_203),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_317),
.A2(n_218),
.B1(n_226),
.B2(n_222),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_299),
.A2(n_236),
.B1(n_219),
.B2(n_213),
.Y(n_355)
);

AND2x4_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_205),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_284),
.A2(n_210),
.B1(n_207),
.B2(n_22),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_280),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_273),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_276),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_270),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_362)
);

AO22x2_ASAP7_75t_L g363 ( 
.A1(n_310),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_307),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_273),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_286),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_310),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_305),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_304),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_286),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_277),
.Y(n_373)
);

OA22x2_ASAP7_75t_L g374 ( 
.A1(n_307),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_300),
.B(n_47),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_276),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_54),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_324),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_325),
.A2(n_272),
.B(n_322),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_353),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_373),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_353),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_327),
.B(n_316),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_335),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

BUFx6f_ASAP7_75t_SL g397 ( 
.A(n_349),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_334),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_354),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_296),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_372),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_333),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_312),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_347),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_342),
.B(n_291),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_351),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_310),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_320),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_351),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_369),
.B(n_320),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_375),
.B(n_320),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_343),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_357),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_346),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_349),
.B(n_291),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_376),
.A2(n_323),
.B(n_282),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_346),
.B(n_291),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_363),
.B(n_291),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_371),
.B(n_55),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_368),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_336),
.A2(n_293),
.B(n_318),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_328),
.Y(n_437)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_328),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_326),
.B(n_302),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_348),
.B(n_309),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_362),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_348),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_330),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_324),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_329),
.B(n_288),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_330),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_334),
.B(n_285),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_330),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_381),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_384),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_290),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_403),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_439),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_389),
.B(n_274),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_385),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_287),
.B(n_315),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_447),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_447),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_405),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_419),
.B(n_409),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_386),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_391),
.B(n_290),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_312),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_415),
.B(n_312),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_420),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_308),
.B(n_274),
.Y(n_471)
);

AND2x2_ASAP7_75t_SL g472 ( 
.A(n_418),
.B(n_410),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_298),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_415),
.B(n_313),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_406),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_274),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_442),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_270),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_418),
.B(n_288),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_421),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_421),
.B(n_313),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_434),
.B(n_431),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_429),
.B(n_281),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_421),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_421),
.B(n_274),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_395),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g491 ( 
.A(n_411),
.B(n_288),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_399),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_413),
.B(n_281),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_428),
.B(n_390),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_428),
.A2(n_274),
.B(n_313),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_401),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_392),
.B(n_313),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_423),
.B(n_294),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_427),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_379),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_422),
.B(n_56),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_436),
.B(n_294),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_383),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_441),
.B(n_294),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_393),
.B(n_394),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_388),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_380),
.B(n_294),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_380),
.B(n_295),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_451),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_425),
.B(n_321),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_411),
.B(n_295),
.Y(n_515)
);

BUFx4f_ASAP7_75t_SL g516 ( 
.A(n_400),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_441),
.B(n_295),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_430),
.B(n_57),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_435),
.B(n_295),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_416),
.A2(n_321),
.B(n_311),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_396),
.B(n_306),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_398),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_398),
.B(n_306),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_417),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_400),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_473),
.B(n_440),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_483),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_396),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_444),
.Y(n_532)
);

BUFx12f_ASAP7_75t_L g533 ( 
.A(n_522),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_483),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_466),
.B(n_402),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_522),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_463),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_503),
.B(n_397),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_477),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_469),
.B(n_424),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_489),
.Y(n_542)
);

NAND2x1_ASAP7_75t_L g543 ( 
.A(n_488),
.B(n_306),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_503),
.B(n_424),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_479),
.B(n_306),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_463),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_464),
.B(n_432),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_473),
.B(n_311),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_522),
.Y(n_549)
);

INVx5_ASAP7_75t_L g550 ( 
.A(n_522),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_489),
.Y(n_551)
);

BUFx8_ASAP7_75t_SL g552 ( 
.A(n_524),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_504),
.B(n_311),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_475),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_475),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_518),
.B(n_397),
.Y(n_556)
);

AND2x2_ASAP7_75t_SL g557 ( 
.A(n_472),
.B(n_378),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_460),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_522),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_504),
.B(n_311),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_487),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_378),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_482),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_518),
.B(n_446),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_491),
.B(n_461),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_524),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_518),
.B(n_446),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_453),
.B(n_58),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_466),
.B(n_321),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_481),
.B(n_59),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_492),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_492),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_519),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_485),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_454),
.B(n_60),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_454),
.B(n_61),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_479),
.B(n_321),
.Y(n_578)
);

NAND2x1_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_62),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_491),
.B(n_65),
.Y(n_580)
);

CKINVDCx8_ASAP7_75t_R g581 ( 
.A(n_494),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_462),
.B(n_67),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_459),
.B(n_68),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_443),
.Y(n_584)
);

CKINVDCx8_ASAP7_75t_R g585 ( 
.A(n_494),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_485),
.B(n_443),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_517),
.B(n_69),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_552),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_537),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_542),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_537),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_542),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_532),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_533),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_575),
.B(n_586),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_538),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_559),
.Y(n_597)
);

BUFx12f_ASAP7_75t_L g598 ( 
.A(n_541),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_541),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_528),
.B(n_514),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_527),
.Y(n_601)
);

BUFx2_ASAP7_75t_R g602 ( 
.A(n_547),
.Y(n_602)
);

INVx5_ASAP7_75t_SL g603 ( 
.A(n_529),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_530),
.B(n_498),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_584),
.A2(n_456),
.B1(n_472),
.B2(n_471),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_550),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_566),
.B(n_507),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_572),
.B(n_507),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_540),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_514),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_576),
.B(n_478),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_551),
.B(n_520),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_527),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_550),
.B(n_489),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_564),
.B(n_520),
.Y(n_616)
);

BUFx2_ASAP7_75t_R g617 ( 
.A(n_535),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_529),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_559),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_538),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_558),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_551),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_554),
.Y(n_623)
);

BUFx12f_ASAP7_75t_L g624 ( 
.A(n_544),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_576),
.B(n_478),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_529),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_534),
.Y(n_627)
);

BUFx24_ASAP7_75t_L g628 ( 
.A(n_544),
.Y(n_628)
);

BUFx6f_ASAP7_75t_SL g629 ( 
.A(n_568),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_554),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_577),
.B(n_498),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_563),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_559),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_550),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_581),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_555),
.Y(n_636)
);

INVx6_ASAP7_75t_L g637 ( 
.A(n_534),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_589),
.Y(n_638)
);

BUFx2_ASAP7_75t_SL g639 ( 
.A(n_610),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_SL g640 ( 
.A1(n_604),
.A2(n_557),
.B1(n_584),
.B2(n_516),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_568),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_589),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_605),
.A2(n_585),
.B1(n_612),
.B2(n_631),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_620),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_610),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_632),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_620),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_630),
.Y(n_648)
);

AOI22xp5_ASAP7_75t_L g649 ( 
.A1(n_600),
.A2(n_565),
.B1(n_493),
.B2(n_452),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_635),
.A2(n_565),
.B1(n_458),
.B2(n_570),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_634),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_630),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_606),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_600),
.A2(n_625),
.B1(n_631),
.B2(n_595),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_608),
.B(n_577),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_625),
.A2(n_532),
.B1(n_583),
.B2(n_555),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_636),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_591),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_606),
.B(n_493),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_637),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_SL g661 ( 
.A1(n_629),
.A2(n_532),
.B1(n_580),
.B2(n_569),
.Y(n_661)
);

BUFx8_ASAP7_75t_SL g662 ( 
.A(n_588),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_SL g663 ( 
.A1(n_629),
.A2(n_532),
.B1(n_569),
.B2(n_486),
.Y(n_663)
);

BUFx4_ASAP7_75t_R g664 ( 
.A(n_588),
.Y(n_664)
);

CKINVDCx6p67_ASAP7_75t_R g665 ( 
.A(n_628),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_618),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_591),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_634),
.Y(n_668)
);

INVx6_ASAP7_75t_L g669 ( 
.A(n_637),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_613),
.A2(n_536),
.B1(n_549),
.B2(n_556),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_634),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_613),
.A2(n_536),
.B1(n_549),
.B2(n_556),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_596),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_618),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_609),
.A2(n_546),
.B1(n_531),
.B2(n_611),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_636),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_598),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_629),
.A2(n_486),
.B1(n_571),
.B2(n_539),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_616),
.A2(n_515),
.B1(n_548),
.B2(n_561),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_598),
.Y(n_681)
);

INVx3_ASAP7_75t_SL g682 ( 
.A(n_665),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_649),
.A2(n_601),
.B1(n_599),
.B2(n_614),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_645),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_643),
.A2(n_635),
.B1(n_624),
.B2(n_614),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_651),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_641),
.B(n_654),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_645),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_640),
.A2(n_602),
.B1(n_635),
.B2(n_617),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_659),
.B(n_635),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_639),
.A2(n_635),
.B1(n_624),
.B2(n_599),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_638),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_655),
.A2(n_601),
.B1(n_593),
.B2(n_594),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_644),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_680),
.A2(n_582),
.B(n_587),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_663),
.A2(n_539),
.B1(n_545),
.B2(n_526),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_644),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_665),
.A2(n_593),
.B1(n_623),
.B2(n_574),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_647),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_650),
.A2(n_623),
.B1(n_613),
.B2(n_496),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_647),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_L g702 ( 
.A1(n_679),
.A2(n_500),
.B(n_508),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_648),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_642),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_646),
.A2(n_571),
.B1(n_494),
.B2(n_465),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_SL g706 ( 
.A1(n_661),
.A2(n_495),
.B(n_621),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_656),
.A2(n_526),
.B1(n_593),
.B2(n_594),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_SL g708 ( 
.A1(n_681),
.A2(n_593),
.B1(n_603),
.B2(n_627),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_656),
.A2(n_496),
.B1(n_553),
.B2(n_560),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_680),
.A2(n_562),
.B1(n_561),
.B2(n_578),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_651),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_653),
.A2(n_593),
.B1(n_603),
.B2(n_534),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_675),
.A2(n_603),
.B1(n_626),
.B2(n_637),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_675),
.A2(n_603),
.B1(n_626),
.B2(n_637),
.Y(n_714)
);

OAI22xp5_ASAP7_75t_L g715 ( 
.A1(n_678),
.A2(n_590),
.B1(n_592),
.B2(n_622),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_658),
.A2(n_562),
.B1(n_480),
.B2(n_490),
.Y(n_716)
);

BUFx4f_ASAP7_75t_SL g717 ( 
.A(n_666),
.Y(n_717)
);

AOI22xp33_ASAP7_75t_L g718 ( 
.A1(n_667),
.A2(n_509),
.B1(n_506),
.B2(n_505),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_660),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_673),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_666),
.B(n_501),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_670),
.A2(n_622),
.B1(n_590),
.B2(n_592),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_648),
.B(n_590),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_676),
.A2(n_592),
.B1(n_622),
.B2(n_457),
.Y(n_724)
);

INVx5_ASAP7_75t_SL g725 ( 
.A(n_651),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_652),
.Y(n_726)
);

BUFx4f_ASAP7_75t_SL g727 ( 
.A(n_674),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_672),
.A2(n_615),
.B1(n_607),
.B2(n_467),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_674),
.A2(n_615),
.B1(n_607),
.B2(n_634),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_657),
.A2(n_457),
.B1(n_579),
.B2(n_619),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_702),
.A2(n_457),
.B1(n_513),
.B2(n_484),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_705),
.A2(n_671),
.B1(n_669),
.B2(n_660),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_689),
.A2(n_677),
.B1(n_657),
.B2(n_669),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_688),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_687),
.A2(n_671),
.B1(n_668),
.B2(n_651),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_683),
.A2(n_669),
.B1(n_660),
.B2(n_468),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_685),
.A2(n_700),
.B1(n_690),
.B2(n_695),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_706),
.A2(n_677),
.B1(n_671),
.B2(n_668),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_696),
.A2(n_474),
.B1(n_497),
.B2(n_668),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_700),
.A2(n_671),
.B1(n_615),
.B2(n_668),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_693),
.A2(n_513),
.B1(n_476),
.B2(n_510),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_684),
.B(n_686),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_709),
.A2(n_662),
.B1(n_671),
.B2(n_513),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_686),
.B(n_597),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_707),
.A2(n_513),
.B1(n_476),
.B2(n_510),
.Y(n_747)
);

OAI222xp33_ASAP7_75t_L g748 ( 
.A1(n_691),
.A2(n_543),
.B1(n_476),
.B2(n_664),
.C1(n_512),
.C2(n_511),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_721),
.A2(n_513),
.B1(n_597),
.B2(n_619),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_711),
.B(n_597),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_694),
.B(n_597),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_711),
.B(n_597),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_SL g753 ( 
.A1(n_698),
.A2(n_634),
.B(n_633),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_698),
.A2(n_633),
.B1(n_619),
.B2(n_502),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_L g755 ( 
.A1(n_682),
.A2(n_633),
.B1(n_619),
.B2(n_502),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_715),
.A2(n_633),
.B1(n_619),
.B2(n_502),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_697),
.B(n_633),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_L g758 ( 
.A1(n_682),
.A2(n_499),
.B1(n_470),
.B2(n_664),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_709),
.A2(n_662),
.B1(n_499),
.B2(n_470),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_717),
.A2(n_499),
.B1(n_72),
.B2(n_77),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_SL g761 ( 
.A1(n_717),
.A2(n_70),
.B1(n_79),
.B2(n_80),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_L g762 ( 
.A1(n_727),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_727),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_699),
.B(n_86),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_712),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_692),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_701),
.B(n_91),
.Y(n_767)
);

AOI211xp5_ASAP7_75t_L g768 ( 
.A1(n_713),
.A2(n_714),
.B(n_729),
.C(n_722),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_L g769 ( 
.A1(n_718),
.A2(n_716),
.B1(n_704),
.B2(n_720),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_735),
.B(n_728),
.Y(n_770)
);

AOI221xp5_ASAP7_75t_L g771 ( 
.A1(n_739),
.A2(n_718),
.B1(n_716),
.B2(n_719),
.C(n_730),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_766),
.B(n_703),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_740),
.B(n_708),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_736),
.B(n_726),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_744),
.B(n_769),
.Y(n_775)
);

OAI21xp33_ASAP7_75t_L g776 ( 
.A1(n_734),
.A2(n_769),
.B(n_759),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_736),
.B(n_725),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_734),
.B(n_723),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_736),
.B(n_746),
.Y(n_779)
);

OAI21xp33_ASAP7_75t_L g780 ( 
.A1(n_759),
.A2(n_724),
.B(n_710),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_736),
.B(n_725),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_SL g782 ( 
.A(n_748),
.B(n_725),
.C(n_724),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_738),
.A2(n_733),
.B1(n_758),
.B2(n_760),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_768),
.B(n_710),
.Y(n_784)
);

INVx1_ASAP7_75t_SL g785 ( 
.A(n_763),
.Y(n_785)
);

OAI221xp5_ASAP7_75t_SL g786 ( 
.A1(n_745),
.A2(n_731),
.B1(n_93),
.B2(n_94),
.C(n_96),
.Y(n_786)
);

NAND3xp33_ASAP7_75t_L g787 ( 
.A(n_761),
.B(n_731),
.C(n_97),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_765),
.B(n_92),
.C(n_98),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_745),
.A2(n_99),
.B1(n_102),
.B2(n_105),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_750),
.B(n_185),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_740),
.B(n_106),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_752),
.B(n_184),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_SL g793 ( 
.A1(n_762),
.A2(n_107),
.B(n_109),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_741),
.B(n_110),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_751),
.B(n_113),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_757),
.B(n_737),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_764),
.B(n_116),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_767),
.B(n_117),
.Y(n_798)
);

OA21x2_ASAP7_75t_L g799 ( 
.A1(n_754),
.A2(n_119),
.B(n_121),
.Y(n_799)
);

NAND4xp25_ASAP7_75t_L g800 ( 
.A(n_732),
.B(n_124),
.C(n_125),
.D(n_128),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_779),
.B(n_753),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_775),
.B(n_747),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_770),
.B(n_742),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_SL g804 ( 
.A1(n_784),
.A2(n_755),
.B1(n_743),
.B2(n_749),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_796),
.B(n_756),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_785),
.B(n_182),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_777),
.B(n_129),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_L g808 ( 
.A(n_794),
.B(n_131),
.C(n_134),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_772),
.B(n_135),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_774),
.Y(n_810)
);

OA21x2_ASAP7_75t_L g811 ( 
.A1(n_773),
.A2(n_137),
.B(n_138),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_778),
.B(n_139),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_781),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_776),
.B(n_140),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_783),
.B(n_141),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_773),
.B(n_142),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_803),
.B(n_795),
.Y(n_817)
);

NOR2x1_ASAP7_75t_L g818 ( 
.A(n_811),
.B(n_799),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_813),
.B(n_790),
.Y(n_819)
);

XNOR2xp5_ASAP7_75t_L g820 ( 
.A(n_807),
.B(n_792),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_810),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_803),
.B(n_794),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_801),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_801),
.Y(n_824)
);

INVx3_ASAP7_75t_SL g825 ( 
.A(n_807),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_821),
.Y(n_826)
);

XOR2x2_ASAP7_75t_L g827 ( 
.A(n_820),
.B(n_816),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_824),
.Y(n_828)
);

XNOR2x2_ASAP7_75t_L g829 ( 
.A(n_818),
.B(n_816),
.Y(n_829)
);

XOR2x2_ASAP7_75t_L g830 ( 
.A(n_825),
.B(n_815),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_826),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_829),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_826),
.Y(n_833)
);

AOI22x1_ASAP7_75t_L g834 ( 
.A1(n_828),
.A2(n_822),
.B1(n_825),
.B2(n_823),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_833),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_833),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_831),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_835),
.A2(n_832),
.B1(n_830),
.B2(n_827),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_836),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_839),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_838),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_SL g842 ( 
.A1(n_839),
.A2(n_832),
.B(n_837),
.C(n_806),
.Y(n_842)
);

NAND4xp25_ASAP7_75t_SL g843 ( 
.A(n_841),
.B(n_823),
.C(n_814),
.D(n_834),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_840),
.B(n_817),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_842),
.Y(n_845)
);

AO22x1_ASAP7_75t_L g846 ( 
.A1(n_841),
.A2(n_807),
.B1(n_791),
.B2(n_809),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_840),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_840),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_847),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_845),
.A2(n_811),
.B1(n_805),
.B2(n_808),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_819),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_848),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_846),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_843),
.Y(n_854)
);

OAI21xp5_ASAP7_75t_L g855 ( 
.A1(n_853),
.A2(n_811),
.B(n_793),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_849),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_852),
.Y(n_857)
);

OAI22x1_ASAP7_75t_L g858 ( 
.A1(n_854),
.A2(n_791),
.B1(n_788),
.B2(n_787),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_851),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_850),
.B(n_812),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_857),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_856),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_859),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_858),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_855),
.B(n_800),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_860),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_L g867 ( 
.A(n_859),
.B(n_797),
.C(n_798),
.Y(n_867)
);

INVxp67_ASAP7_75t_SL g868 ( 
.A(n_857),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_857),
.Y(n_869)
);

OAI22x1_ASAP7_75t_L g870 ( 
.A1(n_859),
.A2(n_809),
.B1(n_799),
.B2(n_805),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_861),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_869),
.A2(n_789),
.B1(n_799),
.B2(n_771),
.Y(n_872)
);

OAI22x1_ASAP7_75t_L g873 ( 
.A1(n_868),
.A2(n_802),
.B1(n_786),
.B2(n_782),
.Y(n_873)
);

AO22x2_ASAP7_75t_L g874 ( 
.A1(n_864),
.A2(n_802),
.B1(n_782),
.B2(n_804),
.Y(n_874)
);

AO22x2_ASAP7_75t_L g875 ( 
.A1(n_862),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_SL g876 ( 
.A1(n_866),
.A2(n_780),
.B1(n_149),
.B2(n_150),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_863),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_865),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_870),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_871),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_879),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_878),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_875),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_876),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_874),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_881),
.A2(n_872),
.B1(n_867),
.B2(n_877),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_880),
.A2(n_873),
.B1(n_157),
.B2(n_158),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_887),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_SL g889 ( 
.A1(n_888),
.A2(n_885),
.B1(n_882),
.B2(n_884),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_889),
.Y(n_890)
);

AOI221xp5_ASAP7_75t_L g891 ( 
.A1(n_890),
.A2(n_886),
.B1(n_883),
.B2(n_163),
.C(n_165),
.Y(n_891)
);

AOI211xp5_ASAP7_75t_L g892 ( 
.A1(n_891),
.A2(n_155),
.B(n_161),
.C(n_167),
.Y(n_892)
);


endmodule