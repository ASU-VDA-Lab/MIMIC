module fake_jpeg_289_n_161 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_161);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_42),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_63),
.B1(n_54),
.B2(n_51),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_40),
.C(n_50),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_56),
.C(n_71),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_46),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_43),
.B1(n_54),
.B2(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_47),
.B1(n_45),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_68),
.B1(n_5),
.B2(n_6),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_43),
.B1(n_48),
.B2(n_55),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_66),
.B1(n_65),
.B2(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_87),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_40),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_84),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_83),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_81),
.B1(n_91),
.B2(n_3),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_82),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_66),
.A2(n_52),
.B1(n_41),
.B2(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_0),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_R g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_89),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_39),
.C(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_95),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_68),
.B(n_5),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_12),
.B(n_13),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_68),
.B1(n_6),
.B2(n_7),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_96),
.A2(n_102),
.B(n_103),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_15),
.B1(n_17),
.B2(n_21),
.Y(n_121)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

OA21x2_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_19),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_37),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_11),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_9),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_9),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_108),
.A2(n_80),
.B1(n_12),
.B2(n_13),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_118),
.B1(n_125),
.B2(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_11),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_121),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_14),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_111),
.B(n_115),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_25),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_24),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_29),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_33),
.B1(n_34),
.B2(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_102),
.B1(n_104),
.B2(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_138),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_120),
.B1(n_112),
.B2(n_125),
.Y(n_137)
);

INVxp33_ASAP7_75t_SL g142 ( 
.A(n_137),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_120),
.B(n_127),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_127),
.Y(n_139)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_119),
.C(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.C(n_135),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_137),
.C(n_136),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_148),
.B(n_149),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_130),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_151),
.B1(n_142),
.B2(n_141),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_141),
.B1(n_129),
.B2(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_153),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_154),
.B(n_152),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_142),
.B(n_133),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_131),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_128),
.Y(n_161)
);


endmodule