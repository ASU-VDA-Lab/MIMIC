module fake_aes_11901_n_38 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx8_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_4), .A2(n_12), .B1(n_1), .B2(n_8), .Y(n_16) );
INVxp67_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_0), .B(n_2), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_7), .Y(n_19) );
BUFx2_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_8), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
A2O1A1Ixp33_ASAP7_75t_L g23 ( .A1(n_18), .A2(n_0), .B(n_1), .C(n_2), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_15), .Y(n_24) );
O2A1O1Ixp33_ASAP7_75t_SL g25 ( .A1(n_23), .A2(n_17), .B(n_21), .C(n_16), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_22), .B(n_20), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
OAI32xp33_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_22), .A3(n_24), .B1(n_25), .B2(n_16), .Y(n_30) );
OAI221xp5_ASAP7_75t_SL g31 ( .A1(n_29), .A2(n_26), .B1(n_15), .B2(n_5), .C(n_6), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g32 ( .A(n_30), .B(n_3), .Y(n_32) );
NAND2x1_ASAP7_75t_L g33 ( .A(n_31), .B(n_14), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_3), .Y(n_34) );
AOI22xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
OAI22xp33_ASAP7_75t_SL g37 ( .A1(n_36), .A2(n_7), .B1(n_9), .B2(n_35), .Y(n_37) );
INVxp67_ASAP7_75t_L g38 ( .A(n_37), .Y(n_38) );
endmodule