module real_jpeg_25522_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_4),
.A2(n_53),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_59),
.B1(n_64),
.B2(n_107),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_36),
.B1(n_38),
.B2(n_107),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_4),
.A2(n_26),
.B1(n_30),
.B2(n_107),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_35),
.B1(n_59),
.B2(n_64),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_6),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_6),
.B(n_58),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_6),
.B(n_36),
.C(n_78),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_6),
.A2(n_59),
.B1(n_64),
.B2(n_173),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_6),
.B(n_123),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_6),
.A2(n_36),
.B1(n_38),
.B2(n_173),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_6),
.B(n_26),
.C(n_41),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_6),
.A2(n_25),
.B(n_263),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_59),
.B1(n_64),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_7),
.A2(n_36),
.B1(n_38),
.B2(n_82),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_53),
.B1(n_82),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_7),
.A2(n_26),
.B1(n_30),
.B2(n_82),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_9),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_9),
.A2(n_56),
.B1(n_59),
.B2(n_64),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_9),
.A2(n_36),
.B1(n_38),
.B2(n_56),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_56),
.Y(n_213)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_11),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_59),
.B1(n_64),
.B2(n_147),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_11),
.A2(n_36),
.B1(n_38),
.B2(n_147),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_11),
.A2(n_26),
.B1(n_30),
.B2(n_147),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_13),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_14),
.A2(n_59),
.B1(n_64),
.B2(n_69),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_14),
.A2(n_36),
.B1(n_38),
.B2(n_69),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_14),
.A2(n_26),
.B1(n_30),
.B2(n_69),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_15),
.A2(n_36),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_26),
.B1(n_30),
.B2(n_45),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_15),
.A2(n_45),
.B1(n_59),
.B2(n_64),
.Y(n_125)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_16),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_137),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_135),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_21),
.B(n_112),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_73),
.C(n_89),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_22),
.A2(n_73),
.B1(n_74),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_22),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_24),
.A2(n_32),
.B1(n_33),
.B2(n_48),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_29),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_25),
.A2(n_29),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_25),
.A2(n_94),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_25),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_25),
.A2(n_179),
.B1(n_181),
.B2(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_25),
.B(n_233),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_25),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_27),
.Y(n_277)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_28),
.Y(n_157)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_28),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_30),
.B(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_44),
.B2(n_46),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_34),
.A2(n_39),
.B1(n_46),
.B2(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_36),
.A2(n_38),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_36),
.B(n_271),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_39),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_39),
.A2(n_46),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_39),
.B(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_39),
.A2(n_46),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_43),
.A2(n_85),
.B1(n_101),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_43),
.A2(n_159),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_43),
.A2(n_200),
.B(n_236),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_43),
.B(n_173),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_46),
.B(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_65),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_51),
.A2(n_57),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_62),
.B1(n_63),
.B2(n_68),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_55),
.B(n_173),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_67),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_57),
.A2(n_65),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_58),
.A2(n_71),
.B1(n_106),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_59),
.A2(n_63),
.B(n_172),
.C(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_59),
.B(n_228),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_SL g174 ( 
.A(n_62),
.B(n_64),
.C(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_71),
.A2(n_111),
.B(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_84),
.B(n_88),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_84),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_83),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_76),
.A2(n_166),
.B(n_168),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_76),
.A2(n_168),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_77),
.A2(n_103),
.B(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_77),
.A2(n_150),
.B(n_209),
.Y(n_208)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_85),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_85),
.A2(n_251),
.B(n_269),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_89),
.A2(n_90),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.C(n_104),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_91),
.A2(n_92),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_93),
.A2(n_98),
.B1(n_99),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_93),
.Y(n_161)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_97),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_102),
.B(n_104),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_110),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_134),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_122),
.A2(n_123),
.B1(n_167),
.B2(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_123),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_130),
.Y(n_134)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_314),
.B(n_320),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_189),
.B(n_313),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_182),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_140),
.B(n_182),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_160),
.C(n_162),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_141),
.A2(n_142),
.B1(n_160),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_148),
.C(n_152),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_158),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_177),
.B1(n_178),
.B2(n_180),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_156),
.B(n_173),
.Y(n_288)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_160),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_162),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_169),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_163),
.B(n_165),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_169),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_170),
.A2(n_171),
.B1(n_176),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_173),
.B(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_177),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_181),
.A2(n_276),
.B(n_285),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_188),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_184),
.B(n_185),
.C(n_188),
.Y(n_319)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_220),
.B(n_307),
.C(n_312),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_214),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_214),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_204),
.C(n_207),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_192),
.A2(n_193),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_202),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_198),
.C(n_202),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_207),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_212),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_212),
.Y(n_245)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_300),
.B(n_306),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_252),
.B(n_299),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_241),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_225),
.B(n_241),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.C(n_238),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_226),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_229),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B(n_232),
.Y(n_229)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_234),
.A2(n_238),
.B1(n_239),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_242),
.B(n_248),
.C(n_249),
.Y(n_305)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_293),
.B(n_298),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_272),
.B(n_292),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_266),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_255),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_260),
.C(n_261),
.Y(n_297)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_262),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_270),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_281),
.B(n_291),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_279),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_286),
.B(n_290),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_297),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_305),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_305),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_319),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_319),
.Y(n_320)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);


endmodule