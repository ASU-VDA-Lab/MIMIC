module real_aes_9162_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_639;
wire n_546;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_686;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_0), .Y(n_588) );
XOR2x2_ASAP7_75t_L g368 ( .A(n_1), .B(n_369), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_2), .A2(n_175), .B1(n_317), .B2(n_514), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_3), .A2(n_133), .B1(n_265), .B2(n_269), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_4), .A2(n_49), .B1(n_372), .B2(n_527), .Y(n_558) );
INVx1_ASAP7_75t_L g496 ( .A(n_5), .Y(n_496) );
AOI222xp33_ASAP7_75t_L g391 ( .A1(n_6), .A2(n_18), .B1(n_182), .B2(n_364), .C1(n_392), .C2(n_393), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_7), .A2(n_131), .B1(n_318), .B2(n_378), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_8), .B(n_373), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_9), .A2(n_79), .B1(n_269), .B2(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_10), .A2(n_237), .B1(n_330), .B2(n_331), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g330 ( .A(n_10), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_11), .A2(n_60), .B1(n_380), .B2(n_382), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_12), .A2(n_436), .B1(n_484), .B2(n_485), .Y(n_435) );
INVx1_ASAP7_75t_L g484 ( .A(n_12), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_13), .A2(n_137), .B1(n_342), .B2(n_714), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_14), .A2(n_71), .B1(n_263), .B2(n_393), .Y(n_530) );
INVx1_ASAP7_75t_L g564 ( .A(n_15), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_16), .B(n_412), .Y(n_708) );
AO22x2_ASAP7_75t_L g245 ( .A1(n_17), .A2(n_65), .B1(n_246), .B2(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g669 ( .A(n_17), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g361 ( .A1(n_19), .A2(n_77), .B1(n_96), .B2(n_282), .C1(n_362), .C2(n_364), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_20), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_21), .A2(n_188), .B1(n_356), .B2(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g424 ( .A(n_22), .Y(n_424) );
CKINVDCx20_ASAP7_75t_R g306 ( .A(n_23), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_24), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_25), .A2(n_146), .B1(n_290), .B2(n_566), .Y(n_565) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_26), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_27), .A2(n_28), .B1(n_372), .B2(n_373), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_29), .A2(n_43), .B1(n_552), .B2(n_553), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_30), .A2(n_169), .B1(n_322), .B2(n_378), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_31), .A2(n_118), .B1(n_339), .B2(n_340), .Y(n_338) );
AO22x2_ASAP7_75t_L g249 ( .A1(n_32), .A2(n_67), .B1(n_246), .B2(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g670 ( .A(n_32), .Y(n_670) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_33), .A2(n_138), .B1(n_265), .B2(n_414), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_34), .A2(n_101), .B1(n_512), .B2(n_514), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_35), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_36), .A2(n_59), .B1(n_340), .B2(n_426), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g536 ( .A1(n_37), .A2(n_40), .B1(n_537), .B2(n_538), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_38), .A2(n_90), .B1(n_356), .B2(n_380), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_39), .A2(n_162), .B1(n_553), .B2(n_635), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_41), .Y(n_703) );
AOI22xp33_ASAP7_75t_SL g524 ( .A1(n_42), .A2(n_210), .B1(n_362), .B2(n_364), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_44), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_45), .B(n_372), .Y(n_614) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_46), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_47), .A2(n_70), .B1(n_454), .B2(n_455), .Y(n_453) );
AOI22xp5_ASAP7_75t_SL g546 ( .A1(n_48), .A2(n_206), .B1(n_547), .B2(n_549), .Y(n_546) );
AOI22xp33_ASAP7_75t_SL g533 ( .A1(n_50), .A2(n_160), .B1(n_446), .B2(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_51), .Y(n_650) );
XOR2x2_ASAP7_75t_L g518 ( .A(n_52), .B(n_519), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_53), .A2(n_209), .B1(n_290), .B2(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_54), .A2(n_168), .B1(n_318), .B2(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_55), .B(n_412), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_56), .A2(n_205), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_57), .A2(n_163), .B1(n_357), .B2(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_58), .A2(n_120), .B1(n_359), .B2(n_360), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_61), .A2(n_149), .B1(n_402), .B2(n_555), .Y(n_677) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_62), .A2(n_114), .B1(n_470), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_63), .A2(n_75), .B1(n_324), .B2(n_327), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_64), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_66), .A2(n_132), .B1(n_263), .B2(n_269), .Y(n_262) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_68), .A2(n_174), .B1(n_386), .B2(n_445), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_69), .A2(n_167), .B1(n_555), .B2(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g230 ( .A(n_72), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_73), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_74), .A2(n_148), .B1(n_327), .B2(n_388), .Y(n_623) );
INVx1_ASAP7_75t_L g226 ( .A(n_76), .Y(n_226) );
INVx1_ASAP7_75t_L g567 ( .A(n_78), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_80), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_81), .A2(n_116), .B1(n_291), .B2(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_82), .A2(n_110), .B1(n_386), .B2(n_429), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_83), .A2(n_190), .B1(n_343), .B2(n_378), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_84), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_85), .Y(n_633) );
INVx1_ASAP7_75t_L g427 ( .A(n_86), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g256 ( .A(n_87), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_88), .A2(n_161), .B1(n_317), .B2(n_320), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_89), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_91), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_92), .A2(n_98), .B1(n_353), .B2(n_363), .Y(n_375) );
INVx1_ASAP7_75t_L g417 ( .A(n_93), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_94), .A2(n_176), .B1(n_455), .B2(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_SL g573 ( .A1(n_95), .A2(n_574), .B1(n_575), .B2(n_601), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_95), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_97), .B(n_431), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_99), .A2(n_216), .B1(n_386), .B2(n_388), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_100), .Y(n_452) );
INVx1_ASAP7_75t_L g422 ( .A(n_102), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_103), .A2(n_104), .B1(n_402), .B2(n_403), .Y(n_401) );
AOI222xp33_ASAP7_75t_L g430 ( .A1(n_105), .A2(n_144), .B1(n_151), .B2(n_284), .C1(n_363), .C2(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_106), .A2(n_135), .B1(n_407), .B2(n_534), .Y(n_678) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_107), .A2(n_136), .B1(n_177), .B2(n_284), .C1(n_289), .C2(n_498), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_108), .A2(n_192), .B1(n_444), .B2(n_549), .Y(n_595) );
AOI22x1_ASAP7_75t_L g627 ( .A1(n_109), .A2(n_628), .B1(n_654), .B2(n_655), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_109), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_111), .Y(n_465) );
AND2x2_ASAP7_75t_L g229 ( .A(n_112), .B(n_230), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_113), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_115), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_117), .A2(n_204), .B1(n_308), .B2(n_342), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_119), .A2(n_193), .B1(n_263), .B2(n_612), .Y(n_682) );
AND2x6_ASAP7_75t_L g225 ( .A(n_121), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_121), .Y(n_663) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_122), .A2(n_185), .B1(n_246), .B2(n_250), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_123), .A2(n_208), .B1(n_405), .B2(n_407), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_124), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_125), .A2(n_673), .B1(n_674), .B2(n_689), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_125), .Y(n_689) );
CKINVDCx20_ASAP7_75t_R g280 ( .A(n_126), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_127), .A2(n_186), .B1(n_308), .B2(n_312), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_128), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_129), .B(n_349), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_130), .Y(n_478) );
INVx1_ASAP7_75t_L g624 ( .A(n_134), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_139), .A2(n_215), .B1(n_325), .B2(n_340), .Y(n_684) );
INVx1_ASAP7_75t_L g409 ( .A(n_140), .Y(n_409) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_141), .A2(n_223), .B(n_231), .C(n_671), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_142), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_143), .A2(n_180), .B1(n_444), .B2(n_446), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_145), .Y(n_366) );
INVx1_ASAP7_75t_L g432 ( .A(n_147), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_150), .A2(n_200), .B1(n_339), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g620 ( .A1(n_152), .A2(n_183), .B1(n_380), .B2(n_508), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_153), .B(n_373), .Y(n_615) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_154), .Y(n_698) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_155), .A2(n_194), .B1(n_246), .B2(n_247), .Y(n_253) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_156), .A2(n_198), .B1(n_325), .B2(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_157), .B(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_158), .Y(n_639) );
AOI22xp33_ASAP7_75t_SL g507 ( .A1(n_159), .A2(n_164), .B1(n_390), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_165), .A2(n_202), .B1(n_263), .B2(n_414), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_166), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_170), .A2(n_201), .B1(n_360), .B2(n_426), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_171), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_172), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_173), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_178), .B(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g616 ( .A1(n_179), .A2(n_219), .B1(n_265), .B2(n_498), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g539 ( .A1(n_181), .A2(n_212), .B1(n_457), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_184), .A2(n_218), .B1(n_444), .B2(n_446), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_185), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_187), .B(n_373), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_189), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_191), .A2(n_197), .B1(n_686), .B2(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g666 ( .A(n_194), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_195), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_196), .A2(n_220), .B1(n_527), .B2(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_199), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_203), .Y(n_523) );
INVx1_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g645 ( .A(n_211), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_213), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_214), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_217), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_221), .B(n_349), .Y(n_529) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_226), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_227), .A2(n_661), .B(n_697), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_488), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_231) );
INVx1_ASAP7_75t_L g656 ( .A(n_232), .Y(n_656) );
AOI22xp5_ASAP7_75t_SL g232 ( .A1(n_233), .A2(n_395), .B1(n_396), .B2(n_487), .Y(n_232) );
INVx1_ASAP7_75t_L g487 ( .A(n_233), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_332), .B2(n_333), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g331 ( .A(n_237), .Y(n_331) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_294), .Y(n_237) );
NOR2xp33_ASAP7_75t_SL g238 ( .A(n_239), .B(n_273), .Y(n_238) );
OAI221xp5_ASAP7_75t_SL g239 ( .A1(n_240), .A2(n_256), .B1(n_257), .B2(n_261), .C(n_262), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_240), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_240), .A2(n_462), .B1(n_644), .B2(n_645), .Y(n_643) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_SL g579 ( .A(n_241), .Y(n_579) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_251), .Y(n_242) );
INVx2_ASAP7_75t_L g300 ( .A(n_243), .Y(n_300) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_249), .Y(n_243) );
AND2x2_ASAP7_75t_L g260 ( .A(n_244), .B(n_249), .Y(n_260) );
AND2x2_ASAP7_75t_L g305 ( .A(n_244), .B(n_279), .Y(n_305) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g268 ( .A(n_245), .B(n_255), .Y(n_268) );
AND2x2_ASAP7_75t_L g272 ( .A(n_245), .B(n_249), .Y(n_272) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g250 ( .A(n_248), .Y(n_250) );
INVx1_ASAP7_75t_L g267 ( .A(n_249), .Y(n_267) );
INVx2_ASAP7_75t_L g279 ( .A(n_249), .Y(n_279) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_252), .B(n_260), .Y(n_259) );
AND2x4_ASAP7_75t_L g304 ( .A(n_252), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g351 ( .A(n_252), .B(n_300), .Y(n_351) );
AND2x6_ASAP7_75t_L g374 ( .A(n_252), .B(n_260), .Y(n_374) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g271 ( .A(n_253), .Y(n_271) );
INVx1_ASAP7_75t_L g278 ( .A(n_253), .Y(n_278) );
INVx1_ASAP7_75t_L g286 ( .A(n_253), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_253), .B(n_255), .Y(n_314) );
AND2x2_ASAP7_75t_L g285 ( .A(n_254), .B(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g311 ( .A(n_255), .B(n_271), .Y(n_311) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g462 ( .A(n_258), .Y(n_462) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx3_ASAP7_75t_L g347 ( .A(n_259), .Y(n_347) );
AND2x2_ASAP7_75t_L g310 ( .A(n_260), .B(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_L g322 ( .A(n_260), .B(n_285), .Y(n_322) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
BUFx3_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
BUFx2_ASAP7_75t_L g560 ( .A(n_265), .Y(n_560) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x6_ASAP7_75t_L g313 ( .A(n_267), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g276 ( .A(n_268), .B(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g291 ( .A(n_268), .B(n_292), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g476 ( .A(n_268), .B(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_SL g393 ( .A(n_269), .Y(n_393) );
BUFx3_ASAP7_75t_L g414 ( .A(n_269), .Y(n_414) );
BUFx6f_ASAP7_75t_L g561 ( .A(n_269), .Y(n_561) );
BUFx2_ASAP7_75t_SL g612 ( .A(n_269), .Y(n_612) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
INVx1_ASAP7_75t_L g483 ( .A(n_270), .Y(n_483) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x6_ASAP7_75t_L g284 ( .A(n_272), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g482 ( .A(n_272), .Y(n_482) );
OAI222xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_280), .B1(n_281), .B2(n_287), .C1(n_288), .C2(n_293), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_275), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_276), .Y(n_363) );
BUFx4f_ASAP7_75t_SL g498 ( .A(n_276), .Y(n_498) );
BUFx2_ASAP7_75t_L g566 ( .A(n_276), .Y(n_566) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_276), .Y(n_705) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g292 ( .A(n_278), .Y(n_292) );
INVx1_ASAP7_75t_L g477 ( .A(n_279), .Y(n_477) );
OAI221xp5_ASAP7_75t_SL g583 ( .A1(n_281), .A2(n_464), .B1(n_584), .B2(n_585), .C(n_586), .Y(n_583) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx4_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g563 ( .A(n_283), .Y(n_563) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_284), .Y(n_392) );
BUFx3_ASAP7_75t_L g495 ( .A(n_284), .Y(n_495) );
INVx2_ASAP7_75t_L g609 ( .A(n_284), .Y(n_609) );
AND2x6_ASAP7_75t_L g299 ( .A(n_285), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g319 ( .A(n_285), .B(n_305), .Y(n_319) );
OAI222xp33_ASAP7_75t_L g646 ( .A1(n_288), .A2(n_466), .B1(n_647), .B2(n_648), .C1(n_649), .C2(n_650), .Y(n_646) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx4f_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g365 ( .A(n_290), .Y(n_365) );
BUFx12f_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_291), .Y(n_431) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_291), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_315), .Y(n_294) );
OAI221xp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_301), .B1(n_302), .B2(n_306), .C(n_307), .Y(n_295) );
OAI221xp5_ASAP7_75t_SL g447 ( .A1(n_296), .A2(n_448), .B1(n_449), .B2(n_452), .C(n_453), .Y(n_447) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
INVx4_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_SL g359 ( .A(n_298), .Y(n_359) );
INVx2_ASAP7_75t_L g553 ( .A(n_298), .Y(n_553) );
INVx1_ASAP7_75t_L g686 ( .A(n_298), .Y(n_686) );
INVx11_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx11_ASAP7_75t_L g387 ( .A(n_299), .Y(n_387) );
INVx3_ASAP7_75t_L g403 ( .A(n_302), .Y(n_403) );
INVx4_ASAP7_75t_L g555 ( .A(n_302), .Y(n_555) );
INVx4_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g357 ( .A(n_304), .Y(n_357) );
INVx2_ASAP7_75t_L g381 ( .A(n_304), .Y(n_381) );
BUFx3_ASAP7_75t_L g451 ( .A(n_304), .Y(n_451) );
BUFx3_ASAP7_75t_L g514 ( .A(n_304), .Y(n_514) );
AND2x2_ASAP7_75t_L g326 ( .A(n_305), .B(n_311), .Y(n_326) );
AND2x4_ASAP7_75t_L g328 ( .A(n_305), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_305), .B(n_311), .Y(n_420) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g390 ( .A(n_309), .Y(n_390) );
BUFx3_ASAP7_75t_L g406 ( .A(n_309), .Y(n_406) );
INVx5_ASAP7_75t_L g445 ( .A(n_309), .Y(n_445) );
INVx4_ASAP7_75t_L g548 ( .A(n_309), .Y(n_548) );
INVx1_ASAP7_75t_L g714 ( .A(n_309), .Y(n_714) );
INVx8_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx6_ASAP7_75t_SL g343 ( .A(n_313), .Y(n_343) );
INVx1_ASAP7_75t_L g329 ( .A(n_314), .Y(n_329) );
NAND2xp33_ASAP7_75t_SL g315 ( .A(n_316), .B(n_323), .Y(n_315) );
BUFx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g454 ( .A(n_318), .Y(n_454) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_318), .Y(n_552) );
INVx3_ASAP7_75t_L g631 ( .A(n_318), .Y(n_631) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_SL g356 ( .A(n_319), .Y(n_356) );
BUFx2_ASAP7_75t_SL g402 ( .A(n_319), .Y(n_402) );
INVx2_ASAP7_75t_L g513 ( .A(n_319), .Y(n_513) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx3_ASAP7_75t_L g429 ( .A(n_321), .Y(n_429) );
INVx2_ASAP7_75t_L g638 ( .A(n_321), .Y(n_638) );
INVx2_ASAP7_75t_L g687 ( .A(n_321), .Y(n_687) );
INVx6_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
BUFx3_ASAP7_75t_L g388 ( .A(n_322), .Y(n_388) );
BUFx3_ASAP7_75t_L g457 ( .A(n_322), .Y(n_457) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g339 ( .A(n_326), .Y(n_339) );
BUFx3_ASAP7_75t_L g378 ( .A(n_326), .Y(n_378) );
BUFx3_ASAP7_75t_L g537 ( .A(n_326), .Y(n_537) );
INVx2_ASAP7_75t_L g441 ( .A(n_327), .Y(n_441) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_327), .Y(n_635) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g340 ( .A(n_328), .Y(n_340) );
INVx1_ASAP7_75t_L g383 ( .A(n_328), .Y(n_383) );
BUFx2_ASAP7_75t_L g506 ( .A(n_328), .Y(n_506) );
BUFx2_ASAP7_75t_SL g538 ( .A(n_328), .Y(n_538) );
BUFx2_ASAP7_75t_SL g556 ( .A(n_328), .Y(n_556) );
BUFx3_ASAP7_75t_L g717 ( .A(n_328), .Y(n_717) );
AND2x2_ASAP7_75t_L g508 ( .A(n_329), .B(n_477), .Y(n_508) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_SL g333 ( .A1(n_334), .A2(n_335), .B1(n_367), .B2(n_394), .Y(n_333) );
INVx3_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
XOR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_366), .Y(n_335) );
NAND4xp75_ASAP7_75t_L g336 ( .A(n_337), .B(n_344), .C(n_354), .D(n_361), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_341), .Y(n_337) );
INVxp67_ASAP7_75t_L g421 ( .A(n_340), .Y(n_421) );
BUFx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g407 ( .A(n_343), .Y(n_407) );
BUFx2_ASAP7_75t_L g446 ( .A(n_343), .Y(n_446) );
BUFx2_ASAP7_75t_L g549 ( .A(n_343), .Y(n_549) );
OA211x2_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B(n_348), .C(n_352), .Y(n_344) );
OA211x2_ASAP7_75t_L g408 ( .A1(n_346), .A2(n_409), .B(n_410), .C(n_413), .Y(n_408) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g582 ( .A(n_347), .Y(n_582) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_349), .Y(n_681) );
INVx5_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
INVx2_ASAP7_75t_L g412 ( .A(n_350), .Y(n_412) );
INVx4_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
INVx2_ASAP7_75t_SL g464 ( .A(n_362), .Y(n_464) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
NAND4xp75_ASAP7_75t_L g369 ( .A(n_370), .B(n_376), .C(n_384), .D(n_391), .Y(n_369) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_371), .B(n_375), .Y(n_370) );
BUFx4f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g528 ( .A(n_374), .Y(n_528) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g600 ( .A(n_378), .Y(n_600) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
INVx4_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx3_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
INVx2_ASAP7_75t_SL g540 ( .A(n_387), .Y(n_540) );
INVx2_ASAP7_75t_L g466 ( .A(n_392), .Y(n_466) );
INVx2_ASAP7_75t_SL g522 ( .A(n_392), .Y(n_522) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_433), .B1(n_434), .B2(n_486), .Y(n_396) );
INVx1_ASAP7_75t_SL g486 ( .A(n_397), .Y(n_486) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
XOR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_432), .Y(n_398) );
NAND4xp75_ASAP7_75t_L g399 ( .A(n_400), .B(n_408), .C(n_415), .D(n_430), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .Y(n_400) );
INVx3_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_416), .B(n_423), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_421), .B2(n_422), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g636 ( .A1(n_418), .A2(n_637), .B1(n_639), .B2(n_640), .C(n_641), .Y(n_636) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g439 ( .A(n_419), .Y(n_439) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_427), .B2(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_458), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_447), .Y(n_437) );
OAI221xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_438) );
BUFx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_445), .Y(n_534) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_449), .A2(n_631), .B1(n_632), .B2(n_633), .C(n_634), .Y(n_630) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_463), .C(n_472), .Y(n_458) );
OAI222xp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_466), .B2(n_467), .C1(n_468), .C2(n_471), .Y(n_463) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_478), .B2(n_479), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_474), .A2(n_479), .B1(n_652), .B2(n_653), .Y(n_651) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx3_ASAP7_75t_L g589 ( .A(n_476), .Y(n_589) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g591 ( .A(n_480), .Y(n_591) );
CKINVDCx16_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g657 ( .A(n_488), .Y(n_657) );
XOR2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_570), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_516), .B1(n_517), .B2(n_569), .Y(n_489) );
INVx3_ASAP7_75t_SL g569 ( .A(n_490), .Y(n_569) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_515), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_492), .B(n_503), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .Y(n_492) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B(n_497), .Y(n_493) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g647 ( .A(n_498), .Y(n_647) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .C(n_502), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
INVx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g712 ( .A(n_513), .Y(n_712) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_541), .B1(n_542), .B2(n_568), .Y(n_517) );
INVx1_ASAP7_75t_L g568 ( .A(n_518), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_531), .C(n_535), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g521 ( .A1(n_522), .A2(n_523), .B(n_524), .Y(n_521) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .C(n_530), .Y(n_525) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_539), .Y(n_535) );
INVx2_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_567), .Y(n_542) );
NOR4xp75_ASAP7_75t_L g543 ( .A(n_544), .B(n_550), .C(n_557), .D(n_562), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_545), .B(n_546), .Y(n_544) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NAND2x1_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OAI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_564), .B(n_565), .Y(n_562) );
XNOR2xp5_ASAP7_75t_SL g570 ( .A(n_571), .B(n_627), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_602), .B2(n_625), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_592), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g576 ( .A(n_577), .B(n_583), .C(n_587), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B1(n_580), .B2(n_581), .Y(n_577) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_590), .B2(n_591), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g626 ( .A(n_605), .Y(n_626) );
XOR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_624), .Y(n_605) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_617), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_613), .Y(n_607) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
OAI21xp5_ASAP7_75t_SL g702 ( .A1(n_609), .A2(n_703), .B(n_704), .Y(n_702) );
NAND3xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .C(n_616), .Y(n_613) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_621), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g655 ( .A(n_628), .Y(n_655) );
AND2x2_ASAP7_75t_SL g628 ( .A(n_629), .B(n_642), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_636), .Y(n_629) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .C(n_651), .Y(n_642) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_660), .B(n_664), .Y(n_659) );
OR2x2_ASAP7_75t_SL g721 ( .A(n_660), .B(n_665), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_662), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_662), .B(n_694), .Y(n_697) );
CKINVDCx16_ASAP7_75t_R g694 ( .A(n_663), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
OAI322xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_690), .A3(n_691), .B1(n_695), .B2(n_698), .C1(n_699), .C2(n_719), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_674), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND4xp75_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .C(n_683), .D(n_688), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_680), .B(n_682), .Y(n_679) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
XOR2x2_ASAP7_75t_L g699 ( .A(n_698), .B(n_700), .Y(n_699) );
NAND3x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_710), .C(n_715), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .Y(n_701) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .C(n_709), .Y(n_706) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_713), .Y(n_710) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
endmodule