module real_aes_9195_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_602;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g549 ( .A1(n_0), .A2(n_156), .B(n_550), .C(n_553), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_1), .B(n_494), .Y(n_554) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
INVx1_ASAP7_75t_L g190 ( .A(n_3), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_4), .B(n_148), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_5), .A2(n_463), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_6), .A2(n_133), .B(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_7), .A2(n_35), .B1(n_142), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_8), .B(n_133), .Y(n_159) );
AND2x6_ASAP7_75t_L g157 ( .A(n_9), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_10), .A2(n_157), .B(n_453), .C(n_455), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_11), .B(n_36), .Y(n_111) );
INVx1_ASAP7_75t_L g138 ( .A(n_12), .Y(n_138) );
INVx1_ASAP7_75t_L g183 ( .A(n_13), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_14), .B(n_146), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_15), .B(n_148), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_16), .B(n_134), .Y(n_195) );
AO32x2_ASAP7_75t_L g217 ( .A1(n_17), .A2(n_133), .A3(n_163), .B1(n_174), .B2(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_18), .B(n_142), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_19), .B(n_134), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_20), .A2(n_52), .B1(n_142), .B2(n_220), .Y(n_221) );
AOI22xp33_ASAP7_75t_SL g242 ( .A1(n_21), .A2(n_79), .B1(n_142), .B2(n_146), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_22), .B(n_142), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_23), .A2(n_174), .B(n_453), .C(n_514), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_24), .A2(n_174), .B(n_453), .C(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_25), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_26), .B(n_176), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_27), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_28), .A2(n_463), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_29), .B(n_176), .Y(n_214) );
INVx2_ASAP7_75t_L g144 ( .A(n_30), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_31), .A2(n_465), .B(n_473), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_32), .B(n_142), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_33), .B(n_176), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_34), .B(n_228), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_37), .B(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_38), .Y(n_459) );
AOI222xp33_ASAP7_75t_SL g121 ( .A1(n_39), .A2(n_77), .B1(n_122), .B2(n_728), .C1(n_729), .C2(n_733), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g728 ( .A(n_39), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_40), .B(n_148), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_41), .B(n_463), .Y(n_480) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_42), .A2(n_76), .B1(n_436), .B2(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_42), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_43), .A2(n_465), .B(n_467), .C(n_473), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_44), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g551 ( .A(n_45), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_46), .A2(n_89), .B1(n_220), .B2(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g468 ( .A(n_47), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_48), .B(n_142), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_49), .B(n_142), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_50), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_51), .B(n_154), .Y(n_153) );
AOI22xp33_ASAP7_75t_SL g199 ( .A1(n_53), .A2(n_57), .B1(n_142), .B2(n_146), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_54), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_55), .B(n_142), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_56), .B(n_142), .Y(n_225) );
INVx1_ASAP7_75t_L g158 ( .A(n_58), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_59), .B(n_463), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_60), .B(n_494), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_61), .A2(n_154), .B(n_186), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_62), .B(n_142), .Y(n_191) );
INVx1_ASAP7_75t_L g137 ( .A(n_63), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_65), .B(n_148), .Y(n_504) );
AO32x2_ASAP7_75t_L g238 ( .A1(n_66), .A2(n_133), .A3(n_174), .B1(n_239), .B2(n_243), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_67), .B(n_149), .Y(n_456) );
INVx1_ASAP7_75t_L g169 ( .A(n_68), .Y(n_169) );
INVx1_ASAP7_75t_L g209 ( .A(n_69), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_70), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_71), .B(n_470), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_72), .A2(n_453), .B(n_473), .C(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_73), .B(n_146), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g489 ( .A(n_74), .Y(n_489) );
INVx1_ASAP7_75t_L g105 ( .A(n_75), .Y(n_105) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_76), .A2(n_125), .B1(n_435), .B2(n_436), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_76), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_78), .B(n_469), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_80), .B(n_220), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_81), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_82), .B(n_146), .Y(n_213) );
INVx2_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_84), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_85), .A2(n_101), .B1(n_112), .B2(n_747), .Y(n_100) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_86), .B(n_173), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_87), .B(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g107 ( .A(n_88), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g439 ( .A(n_88), .B(n_109), .Y(n_439) );
INVx2_ASAP7_75t_L g727 ( .A(n_88), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_90), .A2(n_99), .B1(n_146), .B2(n_147), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_91), .B(n_463), .Y(n_500) );
INVx1_ASAP7_75t_L g503 ( .A(n_92), .Y(n_503) );
INVxp67_ASAP7_75t_L g492 ( .A(n_93), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_94), .B(n_146), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_95), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g449 ( .A(n_96), .Y(n_449) );
INVx1_ASAP7_75t_L g527 ( .A(n_97), .Y(n_527) );
AND2x2_ASAP7_75t_L g475 ( .A(n_98), .B(n_176), .Y(n_475) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g748 ( .A(n_102), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_107), .Y(n_119) );
INVx1_ASAP7_75t_SL g746 ( .A(n_107), .Y(n_746) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_108), .B(n_727), .Y(n_735) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g726 ( .A(n_109), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AOI22x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_121), .B1(n_736), .B2(n_737), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g736 ( .A(n_116), .Y(n_736) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_118), .A2(n_738), .B(n_745), .Y(n_737) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_437), .B1(n_440), .B2(n_724), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_124), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
INVx2_ASAP7_75t_L g435 ( .A(n_125), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_125), .A2(n_435), .B1(n_742), .B2(n_743), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g125 ( .A(n_126), .B(n_359), .Y(n_125) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_317), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_257), .C(n_293), .D(n_307), .Y(n_127) );
OAI221xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_201), .B1(n_233), .B2(n_244), .C(n_248), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_129), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_177), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_160), .Y(n_131) );
AND2x2_ASAP7_75t_L g254 ( .A(n_132), .B(n_161), .Y(n_254) );
INVx3_ASAP7_75t_L g262 ( .A(n_132), .Y(n_262) );
AND2x2_ASAP7_75t_L g316 ( .A(n_132), .B(n_180), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_132), .B(n_179), .Y(n_352) );
AND2x2_ASAP7_75t_L g410 ( .A(n_132), .B(n_272), .Y(n_410) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_139), .B(n_159), .Y(n_132) );
INVx4_ASAP7_75t_L g200 ( .A(n_133), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_133), .A2(n_480), .B(n_481), .Y(n_479) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_133), .Y(n_486) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_135), .B(n_136), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
OAI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_151), .B(n_157), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_145), .B(n_148), .Y(n_140) );
INVx3_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_142), .Y(n_529) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
BUFx3_ASAP7_75t_L g241 ( .A(n_143), .Y(n_241) );
AND2x6_ASAP7_75t_L g453 ( .A(n_143), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx1_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
INVx2_ASAP7_75t_L g184 ( .A(n_146), .Y(n_184) );
INVx3_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g156 ( .A(n_148), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_148), .A2(n_166), .B(n_167), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_SL g207 ( .A1(n_148), .A2(n_208), .B(n_209), .C(n_210), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_148), .B(n_492), .Y(n_491) );
INVx5_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OAI22xp5_ASAP7_75t_SL g239 ( .A1(n_149), .A2(n_173), .B1(n_240), .B2(n_242), .Y(n_239) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
INVx1_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
AND2x2_ASAP7_75t_L g451 ( .A(n_150), .B(n_155), .Y(n_451) );
INVx1_ASAP7_75t_L g454 ( .A(n_150), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_156), .Y(n_151) );
INVx2_ASAP7_75t_L g170 ( .A(n_154), .Y(n_170) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_156), .A2(n_170), .B(n_190), .C(n_191), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_156), .A2(n_173), .B1(n_198), .B2(n_199), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_156), .A2(n_173), .B1(n_219), .B2(n_221), .Y(n_218) );
BUFx3_ASAP7_75t_L g174 ( .A(n_157), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g181 ( .A1(n_157), .A2(n_182), .B(n_189), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_157), .A2(n_207), .B(n_211), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_157), .A2(n_224), .B(n_229), .Y(n_223) );
NAND2x1p5_ASAP7_75t_L g450 ( .A(n_157), .B(n_451), .Y(n_450) );
AND2x4_ASAP7_75t_L g463 ( .A(n_157), .B(n_451), .Y(n_463) );
INVx4_ASAP7_75t_SL g474 ( .A(n_157), .Y(n_474) );
AND2x2_ASAP7_75t_L g245 ( .A(n_160), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g259 ( .A(n_160), .B(n_180), .Y(n_259) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_161), .B(n_180), .Y(n_274) );
AND2x2_ASAP7_75t_L g286 ( .A(n_161), .B(n_262), .Y(n_286) );
OR2x2_ASAP7_75t_L g288 ( .A(n_161), .B(n_246), .Y(n_288) );
AND2x2_ASAP7_75t_L g323 ( .A(n_161), .B(n_246), .Y(n_323) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_161), .Y(n_368) );
INVx1_ASAP7_75t_L g376 ( .A(n_161), .Y(n_376) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_175), .Y(n_161) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_162), .A2(n_181), .B(n_192), .Y(n_180) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_163), .B(n_459), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_174), .Y(n_164) );
O2A1O1Ixp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_172), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_170), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_172), .A2(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g552 ( .A(n_173), .Y(n_552) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_174), .B(n_197), .C(n_200), .Y(n_196) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_176), .A2(n_206), .B(n_214), .Y(n_205) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_176), .A2(n_223), .B(n_232), .Y(n_222) );
INVx2_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_176), .A2(n_462), .B(n_464), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_176), .A2(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g520 ( .A(n_176), .Y(n_520) );
OAI221xp5_ASAP7_75t_L g293 ( .A1(n_177), .A2(n_294), .B1(n_298), .B2(n_302), .C(n_303), .Y(n_293) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g253 ( .A(n_178), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_193), .Y(n_178) );
INVx2_ASAP7_75t_L g252 ( .A(n_179), .Y(n_252) );
AND2x2_ASAP7_75t_L g305 ( .A(n_179), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_179), .B(n_262), .Y(n_324) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g387 ( .A(n_180), .B(n_262), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_186), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g455 ( .A1(n_184), .A2(n_456), .B(n_457), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_184), .A2(n_483), .B(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_186), .A2(n_527), .B(n_528), .C(n_529), .Y(n_526) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_187), .A2(n_212), .B(n_213), .Y(n_211) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g470 ( .A(n_188), .Y(n_470) );
AND2x2_ASAP7_75t_L g309 ( .A(n_193), .B(n_254), .Y(n_309) );
OAI322xp33_ASAP7_75t_L g377 ( .A1(n_193), .A2(n_333), .A3(n_378), .B1(n_380), .B2(n_383), .C1(n_385), .C2(n_389), .Y(n_377) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2x1_ASAP7_75t_L g260 ( .A(n_194), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g273 ( .A(n_194), .Y(n_273) );
AND2x2_ASAP7_75t_L g382 ( .A(n_194), .B(n_262), .Y(n_382) );
AND2x2_ASAP7_75t_L g414 ( .A(n_194), .B(n_286), .Y(n_414) );
OR2x2_ASAP7_75t_L g417 ( .A(n_194), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g247 ( .A(n_195), .Y(n_247) );
AO21x1_ASAP7_75t_L g246 ( .A1(n_197), .A2(n_200), .B(n_247), .Y(n_246) );
AO21x2_ASAP7_75t_L g447 ( .A1(n_200), .A2(n_448), .B(n_458), .Y(n_447) );
INVx3_ASAP7_75t_L g494 ( .A(n_200), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_200), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_200), .A2(n_524), .B(n_531), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_200), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_215), .Y(n_202) );
INVx1_ASAP7_75t_L g430 ( .A(n_203), .Y(n_430) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g235 ( .A(n_204), .B(n_222), .Y(n_235) );
INVx2_ASAP7_75t_L g270 ( .A(n_204), .Y(n_270) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g292 ( .A(n_205), .Y(n_292) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_205), .Y(n_300) );
OR2x2_ASAP7_75t_L g424 ( .A(n_205), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g249 ( .A(n_215), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g289 ( .A(n_215), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g341 ( .A(n_215), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
AND2x2_ASAP7_75t_L g236 ( .A(n_216), .B(n_237), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g296 ( .A(n_216), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g350 ( .A(n_216), .B(n_238), .Y(n_350) );
OR2x2_ASAP7_75t_L g358 ( .A(n_216), .B(n_292), .Y(n_358) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
BUFx2_ASAP7_75t_L g267 ( .A(n_217), .Y(n_267) );
AND2x2_ASAP7_75t_L g277 ( .A(n_217), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g301 ( .A(n_217), .B(n_222), .Y(n_301) );
AND2x2_ASAP7_75t_L g365 ( .A(n_217), .B(n_238), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_222), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_222), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g278 ( .A(n_222), .Y(n_278) );
INVx1_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
AND2x2_ASAP7_75t_L g295 ( .A(n_222), .B(n_296), .Y(n_295) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_222), .Y(n_373) );
INVx1_ASAP7_75t_L g425 ( .A(n_222), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g402 ( .A(n_234), .B(n_311), .Y(n_402) );
INVx2_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g329 ( .A(n_236), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g428 ( .A(n_236), .B(n_363), .Y(n_428) );
INVx1_ASAP7_75t_L g250 ( .A(n_237), .Y(n_250) );
AND2x2_ASAP7_75t_L g276 ( .A(n_237), .B(n_270), .Y(n_276) );
BUFx2_ASAP7_75t_L g335 ( .A(n_237), .Y(n_335) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_238), .Y(n_256) );
INVx1_ASAP7_75t_L g266 ( .A(n_238), .Y(n_266) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_241), .Y(n_472) );
INVx2_ASAP7_75t_L g553 ( .A(n_241), .Y(n_553) );
INVx1_ASAP7_75t_L g517 ( .A(n_243), .Y(n_517) );
NOR2xp67_ASAP7_75t_L g404 ( .A(n_244), .B(n_251), .Y(n_404) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AOI32xp33_ASAP7_75t_L g248 ( .A1(n_245), .A2(n_249), .A3(n_251), .B1(n_253), .B2(n_255), .Y(n_248) );
AND2x2_ASAP7_75t_L g388 ( .A(n_245), .B(n_261), .Y(n_388) );
AND2x2_ASAP7_75t_L g426 ( .A(n_245), .B(n_324), .Y(n_426) );
INVx1_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_250), .B(n_312), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_251), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_251), .B(n_254), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_251), .B(n_323), .Y(n_405) );
OR2x2_ASAP7_75t_L g419 ( .A(n_251), .B(n_288), .Y(n_419) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g346 ( .A(n_252), .B(n_254), .Y(n_346) );
OR2x2_ASAP7_75t_L g355 ( .A(n_252), .B(n_342), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_254), .B(n_305), .Y(n_327) );
INVx2_ASAP7_75t_L g342 ( .A(n_256), .Y(n_342) );
OR2x2_ASAP7_75t_L g357 ( .A(n_256), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g372 ( .A(n_256), .B(n_373), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_256), .A2(n_349), .B(n_430), .C(n_431), .Y(n_429) );
OAI321xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_263), .A3(n_268), .B1(n_271), .B2(n_275), .C(n_279), .Y(n_257) );
INVx1_ASAP7_75t_L g370 ( .A(n_258), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g381 ( .A(n_259), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_262), .B(n_376), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_263), .A2(n_401), .B1(n_403), .B2(n_405), .C(n_406), .Y(n_400) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
AND2x2_ASAP7_75t_L g338 ( .A(n_265), .B(n_312), .Y(n_338) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_266), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g311 ( .A(n_267), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_268), .A2(n_309), .B(n_354), .C(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g320 ( .A(n_270), .B(n_277), .Y(n_320) );
BUFx2_ASAP7_75t_L g330 ( .A(n_270), .Y(n_330) );
INVx1_ASAP7_75t_L g345 ( .A(n_270), .Y(n_345) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR2x2_ASAP7_75t_L g351 ( .A(n_273), .B(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g434 ( .A(n_273), .Y(n_434) );
INVx1_ASAP7_75t_L g427 ( .A(n_274), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g280 ( .A(n_276), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g384 ( .A(n_276), .B(n_301), .Y(n_384) );
INVx1_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_284), .B1(n_287), .B2(n_289), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_281), .B(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g349 ( .A(n_282), .B(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_283), .B(n_292), .Y(n_312) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g304 ( .A(n_286), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g314 ( .A(n_288), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_291), .A2(n_409), .B1(n_411), .B2(n_412), .C(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g297 ( .A(n_292), .Y(n_297) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_292), .Y(n_363) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_295), .B(n_414), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_296), .A2(n_301), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_299), .B(n_309), .Y(n_406) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g375 ( .A(n_300), .Y(n_375) );
AND2x2_ASAP7_75t_L g334 ( .A(n_301), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g423 ( .A(n_301), .Y(n_423) );
INVx1_ASAP7_75t_L g339 ( .A(n_304), .Y(n_339) );
INVx1_ASAP7_75t_L g394 ( .A(n_305), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_310), .B1(n_313), .B2(n_314), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_311), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g379 ( .A(n_312), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_312), .B(n_350), .Y(n_416) );
OR2x2_ASAP7_75t_L g389 ( .A(n_313), .B(n_342), .Y(n_389) );
INVx1_ASAP7_75t_L g328 ( .A(n_314), .Y(n_328) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_316), .B(n_367), .Y(n_366) );
NOR3xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_336), .C(n_347), .Y(n_317) );
OAI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_325), .C(n_331), .Y(n_318) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_320), .A2(n_391), .B1(n_395), .B2(n_398), .C(n_400), .Y(n_390) );
INVx1_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g332 ( .A(n_323), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g386 ( .A(n_323), .B(n_387), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_324), .A2(n_372), .B(n_374), .C(n_376), .Y(n_371) );
INVx2_ASAP7_75t_L g418 ( .A(n_324), .Y(n_418) );
OAI21xp5_ASAP7_75t_SL g325 ( .A1(n_326), .A2(n_328), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g397 ( .A(n_330), .B(n_350), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
OAI21xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B(n_340), .Y(n_336) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI21xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_343), .B(n_346), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_341), .B(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_346), .B(n_433), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_351), .B(n_353), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g374 ( .A(n_350), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND4x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_390), .C(n_407), .D(n_429), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_377), .Y(n_360) );
OAI211xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_366), .B(n_369), .C(n_371), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_365), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_376), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_388), .Y(n_385) );
INVx1_ASAP7_75t_L g411 ( .A(n_386), .Y(n_411) );
INVx2_ASAP7_75t_SL g399 ( .A(n_387), .Y(n_399) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g412 ( .A(n_397), .Y(n_412) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_SL g407 ( .A(n_408), .B(n_415), .Y(n_407) );
INVx1_ASAP7_75t_SL g409 ( .A(n_410), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_417), .B1(n_419), .B2(n_420), .C(n_421), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g730 ( .A(n_438), .Y(n_730) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g731 ( .A(n_440), .Y(n_731) );
OR3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_622), .C(n_687), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g441 ( .A(n_442), .B(n_563), .C(n_589), .D(n_612), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_495), .B1(n_533), .B2(n_540), .C(n_555), .Y(n_442) );
CKINVDCx14_ASAP7_75t_R g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_444), .A2(n_556), .B1(n_580), .B2(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_476), .Y(n_444) );
INVx1_ASAP7_75t_SL g616 ( .A(n_445), .Y(n_616) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_460), .Y(n_445) );
OR2x2_ASAP7_75t_L g538 ( .A(n_446), .B(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g558 ( .A(n_446), .B(n_477), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_446), .B(n_485), .Y(n_571) );
AND2x2_ASAP7_75t_L g588 ( .A(n_446), .B(n_460), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_446), .B(n_536), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_446), .B(n_587), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_446), .B(n_476), .Y(n_709) );
AOI211xp5_ASAP7_75t_SL g720 ( .A1(n_446), .A2(n_626), .B(n_721), .C(n_722), .Y(n_720) );
INVx5_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_447), .B(n_477), .Y(n_592) );
AND2x2_ASAP7_75t_L g595 ( .A(n_447), .B(n_478), .Y(n_595) );
OR2x2_ASAP7_75t_L g640 ( .A(n_447), .B(n_477), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_447), .B(n_485), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B(n_452), .Y(n_448) );
INVx5_ASAP7_75t_L g466 ( .A(n_453), .Y(n_466) );
INVx5_ASAP7_75t_SL g539 ( .A(n_460), .Y(n_539) );
AND2x2_ASAP7_75t_L g557 ( .A(n_460), .B(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_460), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g643 ( .A(n_460), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g675 ( .A(n_460), .B(n_485), .Y(n_675) );
OR2x2_ASAP7_75t_L g681 ( .A(n_460), .B(n_571), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_460), .B(n_631), .Y(n_690) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_475), .Y(n_460) );
BUFx2_ASAP7_75t_L g512 ( .A(n_463), .Y(n_512) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_466), .A2(n_474), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g547 ( .A1(n_466), .A2(n_474), .B(n_548), .C(n_549), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B(n_471), .C(n_472), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_469), .A2(n_472), .B(n_503), .C(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_485), .Y(n_476) );
AND2x2_ASAP7_75t_L g572 ( .A(n_477), .B(n_539), .Y(n_572) );
INVx1_ASAP7_75t_SL g585 ( .A(n_477), .Y(n_585) );
OR2x2_ASAP7_75t_L g620 ( .A(n_477), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g626 ( .A(n_477), .B(n_485), .Y(n_626) );
AND2x2_ASAP7_75t_L g684 ( .A(n_477), .B(n_536), .Y(n_684) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_478), .B(n_539), .Y(n_611) );
INVx3_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
OR2x2_ASAP7_75t_L g577 ( .A(n_485), .B(n_539), .Y(n_577) );
AND2x2_ASAP7_75t_L g587 ( .A(n_485), .B(n_585), .Y(n_587) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_485), .Y(n_635) );
AND2x2_ASAP7_75t_L g644 ( .A(n_485), .B(n_558), .Y(n_644) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_493), .Y(n_485) );
OA21x2_ASAP7_75t_L g545 ( .A1(n_494), .A2(n_546), .B(n_554), .Y(n_545) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_495), .A2(n_661), .B1(n_663), .B2(n_665), .C(n_668), .Y(n_660) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
AND2x2_ASAP7_75t_L g634 ( .A(n_497), .B(n_615), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_497), .B(n_693), .Y(n_697) );
OR2x2_ASAP7_75t_L g718 ( .A(n_497), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_497), .B(n_723), .Y(n_722) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx5_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
AND2x2_ASAP7_75t_L g642 ( .A(n_498), .B(n_509), .Y(n_642) );
AND2x2_ASAP7_75t_L g703 ( .A(n_498), .B(n_582), .Y(n_703) );
AND2x2_ASAP7_75t_L g716 ( .A(n_498), .B(n_536), .Y(n_716) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_521), .Y(n_507) );
AND2x4_ASAP7_75t_L g543 ( .A(n_508), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g561 ( .A(n_508), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
AND2x2_ASAP7_75t_L g637 ( .A(n_508), .B(n_615), .Y(n_637) );
AND2x2_ASAP7_75t_L g647 ( .A(n_508), .B(n_565), .Y(n_647) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_508), .Y(n_655) );
AND2x2_ASAP7_75t_L g667 ( .A(n_508), .B(n_545), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_508), .B(n_599), .Y(n_671) );
AND2x2_ASAP7_75t_L g708 ( .A(n_508), .B(n_703), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_508), .B(n_582), .Y(n_719) );
OR2x2_ASAP7_75t_L g721 ( .A(n_508), .B(n_657), .Y(n_721) );
INVx5_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g607 ( .A(n_509), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g617 ( .A(n_509), .B(n_562), .Y(n_617) );
AND2x2_ASAP7_75t_L g629 ( .A(n_509), .B(n_545), .Y(n_629) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_509), .Y(n_659) );
AND2x4_ASAP7_75t_L g693 ( .A(n_509), .B(n_544), .Y(n_693) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_518), .Y(n_509) );
AOI21xp5_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_513), .B(n_517), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
BUFx2_ASAP7_75t_L g542 ( .A(n_521), .Y(n_542) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g582 ( .A(n_522), .Y(n_582) );
AND2x2_ASAP7_75t_L g615 ( .A(n_522), .B(n_545), .Y(n_615) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g562 ( .A(n_523), .B(n_545), .Y(n_562) );
BUFx2_ASAP7_75t_L g608 ( .A(n_523), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_535), .B(n_616), .Y(n_695) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_536), .B(n_558), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_536), .B(n_539), .Y(n_597) );
AND2x2_ASAP7_75t_L g652 ( .A(n_536), .B(n_588), .Y(n_652) );
AOI221xp5_ASAP7_75t_SL g589 ( .A1(n_537), .A2(n_590), .B1(n_598), .B2(n_600), .C(n_604), .Y(n_589) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x2_ASAP7_75t_L g584 ( .A(n_538), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g625 ( .A(n_538), .B(n_626), .Y(n_625) );
OAI321xp33_ASAP7_75t_L g632 ( .A1(n_538), .A2(n_591), .A3(n_633), .B1(n_635), .B2(n_636), .C(n_638), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_539), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_542), .B(n_693), .Y(n_711) );
AND2x2_ASAP7_75t_L g598 ( .A(n_543), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_543), .B(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_544), .Y(n_574) );
AND2x2_ASAP7_75t_L g581 ( .A(n_544), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_544), .B(n_656), .Y(n_686) );
INVx1_ASAP7_75t_L g723 ( .A(n_544), .Y(n_723) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B(n_560), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_557), .A2(n_667), .B(n_716), .C(n_717), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_558), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_558), .B(n_596), .Y(n_662) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g605 ( .A(n_562), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_562), .B(n_565), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_562), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_562), .B(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_566), .B1(n_578), .B2(n_583), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g579 ( .A(n_565), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g602 ( .A(n_565), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g614 ( .A(n_565), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_565), .B(n_608), .Y(n_650) );
OR2x2_ASAP7_75t_L g657 ( .A(n_565), .B(n_582), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_565), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g707 ( .A(n_565), .B(n_693), .Y(n_707) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_569), .B1(n_573), .B2(n_575), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g613 ( .A(n_568), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g653 ( .A1(n_571), .A2(n_586), .B1(n_654), .B2(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g701 ( .A(n_572), .Y(n_701) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_576), .A2(n_613), .B1(n_616), .B2(n_617), .C(n_618), .Y(n_612) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g591 ( .A(n_577), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_581), .B(n_647), .Y(n_679) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_582), .Y(n_599) );
INVx1_ASAP7_75t_L g603 ( .A(n_582), .Y(n_603) );
NAND2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx1_ASAP7_75t_L g621 ( .A(n_588), .Y(n_621) );
AND2x2_ASAP7_75t_L g630 ( .A(n_588), .B(n_631), .Y(n_630) );
NAND2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AND2x2_ASAP7_75t_L g674 ( .A(n_595), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_624), .B1(n_627), .B2(n_630), .C(n_632), .Y(n_623) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_602), .B(n_659), .Y(n_658) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_606), .B(n_609), .Y(n_604) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
CKINVDCx16_ASAP7_75t_R g706 ( .A(n_609), .Y(n_706) );
OR2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g648 ( .A(n_611), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g669 ( .A(n_614), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_614), .B(n_674), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_617), .B(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g622 ( .A(n_623), .B(n_641), .C(n_660), .D(n_673), .Y(n_622) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g631 ( .A(n_626), .Y(n_631) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g664 ( .A(n_635), .B(n_640), .Y(n_664) );
INVxp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B(n_645), .C(n_653), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g712 ( .A1(n_643), .A2(n_685), .B(n_713), .C(n_720), .Y(n_712) );
INVx1_ASAP7_75t_SL g672 ( .A(n_644), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_648), .B1(n_650), .B2(n_651), .Y(n_645) );
INVx1_ASAP7_75t_L g676 ( .A(n_650), .Y(n_676) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_656), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_656), .B(n_667), .Y(n_700) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g677 ( .A(n_667), .Y(n_677) );
AOI21xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_672), .Y(n_668) );
INVxp33_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
AOI322xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_676), .A3(n_677), .B1(n_678), .B2(n_680), .C1(n_682), .C2(n_685), .Y(n_673) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
NAND3xp33_ASAP7_75t_SL g687 ( .A(n_688), .B(n_705), .C(n_712), .Y(n_687) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B1(n_694), .B2(n_696), .C(n_698), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g704 ( .A(n_693), .Y(n_704) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_701), .B2(n_702), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_707), .B1(n_708), .B2(n_709), .C(n_710), .Y(n_705) );
NAND2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g732 ( .A(n_725), .Y(n_732) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx3_ASAP7_75t_SL g734 ( .A(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
endmodule