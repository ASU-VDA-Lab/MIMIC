module fake_jpeg_27633_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_36),
.B(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_45),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_17),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_19),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_18),
.B1(n_19),
.B2(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_19),
.B1(n_34),
.B2(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_38),
.B1(n_46),
.B2(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_36),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_23),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_32),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_17),
.B1(n_22),
.B2(n_30),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_38),
.B(n_21),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_81),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_66),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_83),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_30),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_87),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_39),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_28),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_25),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_65),
.B1(n_55),
.B2(n_49),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_51),
.A2(n_23),
.B(n_40),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_39),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_99),
.Y(n_120)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_70),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_115),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_74),
.A2(n_54),
.B1(n_65),
.B2(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_116),
.B1(n_109),
.B2(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_58),
.B1(n_60),
.B2(n_27),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_84),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_58),
.B1(n_40),
.B2(n_20),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_27),
.B1(n_61),
.B2(n_70),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_26),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_26),
.C(n_27),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_76),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_43),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_134),
.B1(n_106),
.B2(n_113),
.Y(n_146)
);

A2O1A1O1Ixp25_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_73),
.B(n_92),
.C(n_26),
.D(n_24),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_93),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_137),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_130),
.B(n_135),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_75),
.B1(n_94),
.B2(n_79),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_33),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_75),
.B1(n_79),
.B2(n_61),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_91),
.C(n_43),
.Y(n_137)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_41),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_118),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_98),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_91),
.C(n_43),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_107),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_141),
.B(n_96),
.Y(n_143)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_127),
.B1(n_16),
.B2(n_15),
.C(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_154),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_124),
.B1(n_138),
.B2(n_125),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_152),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_150),
.A2(n_155),
.B(n_157),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_124),
.B1(n_126),
.B2(n_121),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_105),
.B1(n_24),
.B2(n_6),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_101),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_133),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_156),
.C(n_154),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_174),
.C(n_143),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_172),
.B1(n_160),
.B2(n_161),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_147),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_144),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_152),
.B1(n_145),
.B2(n_163),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_132),
.C(n_140),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_129),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_159),
.B(n_157),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_178),
.B(n_182),
.Y(n_197)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_16),
.C(n_13),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_1),
.B(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_3),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_191),
.B1(n_198),
.B2(n_178),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_195),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_188),
.B(n_193),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_148),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_196),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_175),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_172),
.A2(n_149),
.B1(n_162),
.B2(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_201),
.C(n_202),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_166),
.Y(n_198)
);

BUFx12f_ASAP7_75t_SL g199 ( 
.A(n_166),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_200),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_4),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_4),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_4),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_205),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_192),
.B(n_167),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_174),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_168),
.C(n_171),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_169),
.C(n_187),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_185),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_173),
.C(n_171),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_214),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_215),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_199),
.B1(n_197),
.B2(n_198),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_217),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_197),
.B(n_176),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_223),
.C(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_224),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_7),
.C(n_8),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_222),
.A2(n_203),
.B1(n_206),
.B2(n_210),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_221),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_229),
.A2(n_232),
.B(n_225),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_225),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_223),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g233 ( 
.A(n_227),
.B(n_219),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_SL g240 ( 
.A(n_233),
.B(n_237),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_236),
.Y(n_239)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_236),
.A2(n_231),
.B(n_235),
.C(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_205),
.B(n_9),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_8),
.C(n_9),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_10),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_240),
.B1(n_239),
.B2(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_244),
.B(n_245),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_11),
.Y(n_247)
);


endmodule