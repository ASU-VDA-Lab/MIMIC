module fake_jpeg_5778_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_24),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_42),
.A2(n_50),
.B1(n_26),
.B2(n_18),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_30),
.B1(n_18),
.B2(n_27),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_35),
.B1(n_34),
.B2(n_37),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

NAND2xp67_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_25),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_68),
.Y(n_96)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_79),
.B1(n_55),
.B2(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_71),
.Y(n_98)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_31),
.B1(n_38),
.B2(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_77),
.Y(n_103)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_35),
.B(n_34),
.C(n_40),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_45),
.C(n_47),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_94),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_93),
.B1(n_108),
.B2(n_32),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_52),
.B1(n_49),
.B2(n_37),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_37),
.B1(n_46),
.B2(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_107),
.B1(n_67),
.B2(n_85),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_104),
.B(n_113),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_37),
.B1(n_55),
.B2(n_40),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_36),
.C(n_53),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_36),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_35),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_78),
.B(n_35),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_28),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_84),
.A2(n_29),
.B(n_16),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_22),
.B(n_16),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_131),
.B(n_143),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_121),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_123),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_125),
.B1(n_130),
.B2(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_25),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_53),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_129),
.Y(n_147)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_115),
.C(n_17),
.Y(n_160)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_67),
.B1(n_39),
.B2(n_27),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_89),
.B(n_36),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_39),
.B1(n_32),
.B2(n_28),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_141),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_39),
.B1(n_32),
.B2(n_28),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_138),
.B1(n_107),
.B2(n_111),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_17),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_71),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_28),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_104),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_109),
.A2(n_53),
.B(n_28),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_128),
.C(n_141),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_152),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_158),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_164),
.B1(n_133),
.B2(n_132),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_156),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_90),
.Y(n_156)
);

OAI22x1_ASAP7_75t_L g157 ( 
.A1(n_131),
.A2(n_102),
.B1(n_105),
.B2(n_98),
.Y(n_157)
);

AOI22x1_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_134),
.B1(n_130),
.B2(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_99),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_170),
.B(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_99),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_166),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_17),
.B(n_25),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_165),
.Y(n_179)
);

CKINVDCx12_ASAP7_75t_R g168 ( 
.A(n_117),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_1),
.Y(n_170)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_1),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_127),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_157),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_176),
.B(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_160),
.B(n_166),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_187),
.B(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_188),
.A2(n_167),
.B1(n_152),
.B2(n_146),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_15),
.B1(n_14),
.B2(n_12),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_193),
.A2(n_194),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_144),
.A2(n_15),
.B1(n_12),
.B2(n_3),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_198),
.A2(n_205),
.B1(n_179),
.B2(n_182),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_167),
.C(n_156),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_212),
.C(n_174),
.Y(n_230)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_206),
.Y(n_226)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_154),
.B(n_172),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_185),
.A2(n_155),
.B(n_161),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_180),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_214),
.Y(n_229)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_171),
.C(n_4),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_2),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_194),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_208),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_230),
.C(n_231),
.Y(n_245)
);

NOR2xp67_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_184),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_234),
.B(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_173),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_178),
.Y(n_232)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_181),
.B1(n_173),
.B2(n_7),
.Y(n_233)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_5),
.C(n_6),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_222),
.A2(n_216),
.B(n_201),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_236),
.A2(n_207),
.B(n_213),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_217),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_220),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_219),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_206),
.B1(n_202),
.B2(n_200),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_202),
.B1(n_205),
.B2(n_227),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_223),
.C(n_228),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_251),
.B(n_252),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_203),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_253),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_211),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_243),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_257),
.B(n_260),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_238),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_235),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_8),
.C(n_9),
.Y(n_269)
);

OAI21x1_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_245),
.B(n_213),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_254),
.A3(n_241),
.B1(n_245),
.B2(n_251),
.C1(n_230),
.C2(n_239),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_261),
.B1(n_263),
.B2(n_268),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_263),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_258),
.C(n_9),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_271),
.C(n_269),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_8),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_271),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_8),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_10),
.Y(n_278)
);


endmodule