module real_jpeg_14573_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_54;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_50;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_47;
wire n_11;
wire n_14;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_12),
.B1(n_13),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_4),
.A2(n_12),
.B1(n_13),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_5),
.B(n_13),
.C(n_31),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_5),
.A2(n_17),
.B1(n_41),
.B2(n_47),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_6),
.A2(n_21),
.B1(n_41),
.B2(n_47),
.Y(n_49)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_36),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_25),
.B(n_35),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_19),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_16),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_13),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_18),
.A2(n_20),
.B1(n_22),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_23),
.A2(n_24),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_32),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_27),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_SL g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_31),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_55),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_50),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_50),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);


endmodule