module fake_jpeg_16061_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_3),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_14),
.B1(n_24),
.B2(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_50),
.B1(n_26),
.B2(n_14),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_14),
.B1(n_26),
.B2(n_16),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_36),
.C(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_59),
.B1(n_44),
.B2(n_45),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

AO22x2_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_36),
.B1(n_29),
.B2(n_32),
.Y(n_55)
);

AO22x1_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_44),
.B1(n_46),
.B2(n_42),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_26),
.B1(n_22),
.B2(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_61),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_22),
.B1(n_34),
.B2(n_30),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_67),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_13),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_23),
.A3(n_20),
.B1(n_16),
.B2(n_13),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_23),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_84),
.B1(n_55),
.B2(n_60),
.Y(n_93)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_45),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_60),
.B1(n_43),
.B2(n_45),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_56),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_44),
.B1(n_47),
.B2(n_36),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_66),
.B(n_47),
.C(n_43),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_74),
.B(n_55),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_91),
.B(n_99),
.Y(n_118)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_55),
.B(n_53),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_102),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_95),
.B1(n_100),
.B2(n_103),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_57),
.B1(n_52),
.B2(n_60),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_87),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_53),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_72),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_43),
.B1(n_64),
.B2(n_22),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_63),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_106),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_22),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

O2A1O1Ixp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_78),
.B(n_87),
.C(n_73),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_120),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_87),
.B1(n_79),
.B2(n_82),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_124),
.B1(n_91),
.B2(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_87),
.B1(n_82),
.B2(n_70),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_77),
.Y(n_126)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_70),
.B1(n_80),
.B2(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_124),
.B1(n_126),
.B2(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_135),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_134),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_142),
.C(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_105),
.B(n_88),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_41),
.B(n_15),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_104),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_72),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_95),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_113),
.B1(n_109),
.B2(n_107),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_119),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_100),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_149),
.C(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_148),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_99),
.C(n_96),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_151),
.A2(n_162),
.B1(n_172),
.B2(n_17),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_127),
.B1(n_112),
.B2(n_115),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_157),
.B1(n_147),
.B2(n_130),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_144),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_128),
.B1(n_139),
.B2(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_111),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_150),
.A2(n_110),
.B1(n_70),
.B2(n_90),
.Y(n_162)
);

XNOR2x1_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_72),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_169),
.Y(n_192)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_168),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_110),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_41),
.B1(n_96),
.B2(n_83),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_173),
.A2(n_17),
.B(n_15),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_147),
.C(n_141),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_177),
.C(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_151),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_135),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_56),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_181),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_71),
.B1(n_54),
.B2(n_2),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_184),
.A2(n_193),
.B1(n_15),
.B2(n_17),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_25),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_10),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_10),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_12),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_196),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_170),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_190),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_173),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_210),
.C(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_180),
.B(n_152),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_152),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_168),
.B1(n_159),
.B2(n_171),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_177),
.C(n_178),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_224),
.C(n_205),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_199),
.B1(n_200),
.B2(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_202),
.A2(n_167),
.B1(n_187),
.B2(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_210),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_166),
.C(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_172),
.C(n_184),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_71),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_231),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_228),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_208),
.C(n_196),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_19),
.C(n_25),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_214),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_215),
.B1(n_213),
.B2(n_225),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_236),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_226),
.A2(n_20),
.B1(n_19),
.B2(n_3),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_20),
.B1(n_19),
.B2(n_4),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_217),
.B(n_19),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_238),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_234),
.A2(n_218),
.B(n_1),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_249),
.B(n_231),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_247),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_248),
.A2(n_241),
.B1(n_246),
.B2(n_243),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_4),
.B(n_6),
.Y(n_262)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_241),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_254),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_227),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_256),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_242),
.A2(n_235),
.B(n_233),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_244),
.B(n_5),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_233),
.B1(n_5),
.B2(n_6),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_25),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_261),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_252),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_260),
.A2(n_250),
.B(n_254),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_259),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_6),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_7),
.B(n_8),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_7),
.B(n_8),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_8),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_266),
.C(n_8),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_9),
.Y(n_273)
);


endmodule