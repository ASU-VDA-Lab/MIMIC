module fake_netlist_6_1485_n_65 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_65);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_65;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_21;
wire n_18;
wire n_24;
wire n_37;
wire n_33;
wire n_54;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_36;
wire n_22;
wire n_26;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_20;
wire n_50;
wire n_49;
wire n_30;
wire n_64;
wire n_43;
wire n_19;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_25;
wire n_40;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_4),
.B(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx6p67_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AND2x4_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_12),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

OA21x2_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_18),
.B(n_25),
.Y(n_40)
);

OAI21x1_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_20),
.B(n_24),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_30),
.B(n_22),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_38),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_31),
.B1(n_34),
.B2(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_31),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_52),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_55),
.Y(n_59)
);

XOR2x2_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_53),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_50),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI21x1_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_25),
.B(n_39),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_62),
.C(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_36),
.Y(n_65)
);


endmodule