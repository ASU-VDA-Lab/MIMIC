module fake_jpeg_13291_n_132 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_132);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_63),
.Y(n_79)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_54),
.B1(n_50),
.B2(n_49),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_46),
.B1(n_51),
.B2(n_55),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_77),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_40),
.B(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_50),
.B1(n_52),
.B2(n_44),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_80),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

XOR2x2_ASAP7_75t_SL g95 ( 
.A(n_83),
.B(n_89),
.Y(n_95)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_0),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_2),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_94),
.B(n_6),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx5_ASAP7_75t_SL g106 ( 
.A(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_3),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_39),
.B1(n_9),
.B2(n_13),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_4),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_108),
.Y(n_114)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_26),
.B(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_103),
.B(n_99),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_109),
.B(n_102),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_8),
.B(n_18),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_117),
.B(n_119),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_19),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_106),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_109),
.B1(n_100),
.B2(n_104),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_118),
.B1(n_110),
.B2(n_114),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_125),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_29),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_31),
.C(n_33),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_35),
.B(n_36),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_38),
.Y(n_132)
);


endmodule