module fake_jpeg_4446_n_280 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_34),
.Y(n_66)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_30),
.Y(n_55)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_48),
.Y(n_79)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g85 ( 
.A(n_49),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_33),
.A2(n_18),
.B1(n_29),
.B2(n_16),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_50),
.A2(n_41),
.B1(n_53),
.B2(n_29),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_31),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_21),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_28),
.Y(n_84)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_22),
.B1(n_20),
.B2(n_18),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_40),
.B1(n_20),
.B2(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_18),
.B(n_29),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_68),
.B(n_66),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_69),
.A2(n_68),
.B1(n_67),
.B2(n_61),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVxp67_ASAP7_75t_SL g93 ( 
.A(n_71),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_58),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_40),
.B1(n_38),
.B2(n_32),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_53),
.B1(n_44),
.B2(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_86),
.B(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_28),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_52),
.C(n_64),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_87),
.C(n_73),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_95),
.B1(n_47),
.B2(n_44),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_55),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_56),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_57),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_110),
.B(n_80),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_59),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_100),
.A2(n_76),
.B(n_79),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_107),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_48),
.B1(n_53),
.B2(n_40),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_76),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_84),
.B1(n_70),
.B2(n_86),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_109),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_126),
.B1(n_131),
.B2(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_96),
.B(n_70),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_118),
.C(n_88),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_117),
.A2(n_17),
.B(n_26),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_84),
.C(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_123),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_77),
.B1(n_84),
.B2(n_69),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_93),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_130),
.A2(n_89),
.B1(n_88),
.B2(n_72),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_77),
.B1(n_44),
.B2(n_47),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_30),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_19),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_124),
.A2(n_90),
.B1(n_102),
.B2(n_110),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_133),
.B(n_122),
.Y(n_164)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_141),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_98),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_17),
.B(n_23),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_103),
.C(n_98),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_114),
.B1(n_113),
.B2(n_118),
.Y(n_161)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_144),
.B(n_151),
.Y(n_180)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_153),
.C(n_105),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_32),
.B1(n_38),
.B2(n_17),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_99),
.B1(n_72),
.B2(n_42),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_156),
.B1(n_78),
.B2(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_150),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_8),
.C(n_14),
.Y(n_150)
);

BUFx24_ASAP7_75t_SL g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_116),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_42),
.C(n_105),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_42),
.B1(n_78),
.B2(n_92),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_105),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_112),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_26),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_117),
.CI(n_111),
.CON(n_160),
.SN(n_160)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_161),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_120),
.B1(n_131),
.B2(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_173),
.C(n_183),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_158),
.B(n_109),
.C(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_121),
.B(n_101),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_172),
.B(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_181),
.B1(n_152),
.B2(n_145),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_139),
.A2(n_112),
.B1(n_38),
.B2(n_49),
.Y(n_177)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_112),
.B1(n_49),
.B2(n_26),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_156),
.B1(n_147),
.B2(n_148),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_141),
.C(n_143),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_186),
.A2(n_188),
.B(n_190),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_191),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_146),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_167),
.B(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_198),
.B1(n_204),
.B2(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_153),
.C(n_143),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_199),
.B(n_161),
.C(n_164),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_202),
.B1(n_163),
.B2(n_182),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_206),
.C(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_172),
.C(n_160),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_25),
.B(n_23),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_187),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_160),
.C(n_170),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_214),
.C(n_219),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_165),
.B1(n_169),
.B2(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_184),
.B1(n_201),
.B2(n_195),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_193),
.B(n_169),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_171),
.B1(n_167),
.B2(n_182),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_216),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_138),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_217),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_27),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_26),
.C(n_25),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_27),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_202),
.B1(n_194),
.B2(n_185),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_224),
.B1(n_230),
.B2(n_0),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_194),
.B1(n_188),
.B2(n_201),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_201),
.B1(n_27),
.B2(n_25),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_8),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_27),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_25),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_7),
.B(n_12),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_236),
.B(n_214),
.C(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_23),
.C(n_17),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_220),
.C(n_221),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_232),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_211),
.C(n_206),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_240),
.C(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_249),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_11),
.C(n_10),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_11),
.C(n_10),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_245),
.C(n_246),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_11),
.C(n_10),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_8),
.C(n_6),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_23),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_248),
.A2(n_250),
.B1(n_228),
.B2(n_232),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_259),
.C(n_260),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_226),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_1),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_223),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_234),
.B(n_6),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_0),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_1),
.Y(n_262)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_1),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_265),
.A2(n_258),
.B(n_4),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_267)
);

OAI321xp33_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_251),
.C(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_5),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_269),
.B(n_271),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_3),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_273),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

OAI21x1_ASAP7_75t_SL g277 ( 
.A1(n_275),
.A2(n_264),
.B(n_272),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_274),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_276),
.C(n_5),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_5),
.Y(n_280)
);


endmodule