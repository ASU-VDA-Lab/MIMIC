module fake_jpeg_10689_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_38),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_40),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_17),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_47),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_49),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_19),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_54),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_16),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_33),
.A2(n_19),
.B1(n_20),
.B2(n_13),
.Y(n_54)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_57),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_64),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_16),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_67),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_13),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_68),
.B1(n_45),
.B2(n_60),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_50),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_41),
.B1(n_32),
.B2(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_54),
.B1(n_47),
.B2(n_38),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_85),
.B1(n_74),
.B2(n_86),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_56),
.A2(n_42),
.B1(n_38),
.B2(n_30),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_69),
.B1(n_59),
.B2(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_23),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_42),
.B1(n_34),
.B2(n_19),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_19),
.B(n_23),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_68),
.B(n_66),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g88 ( 
.A(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_91),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_56),
.B1(n_65),
.B2(n_55),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_90),
.A2(n_98),
.B1(n_80),
.B2(n_76),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_94),
.Y(n_110)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_72),
.C(n_58),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_57),
.C(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_71),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_71),
.B(n_24),
.Y(n_106)
);

OAI22x1_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_75),
.B1(n_77),
.B2(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_106),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_83),
.B(n_76),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_22),
.B(n_18),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_96),
.B1(n_97),
.B2(n_95),
.Y(n_113)
);

OAI321xp33_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_90),
.A3(n_96),
.B1(n_89),
.B2(n_91),
.C(n_98),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_93),
.C(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_107),
.C(n_103),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_101),
.Y(n_123)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_25),
.B1(n_22),
.B2(n_18),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_110),
.Y(n_119)
);

NAND4xp25_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_115),
.C(n_118),
.D(n_18),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_124),
.B1(n_8),
.B2(n_12),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_109),
.B1(n_25),
.B2(n_5),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_125),
.A2(n_119),
.B(n_18),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_121),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_122),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_125),
.A2(n_122),
.B1(n_120),
.B2(n_123),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_127),
.B(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_9),
.B1(n_10),
.B2(n_4),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_133),
.Y(n_135)
);


endmodule