module real_jpeg_25781_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_300;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_297;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_269;
wire n_96;
wire n_273;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_0),
.A2(n_64),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_0),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_0),
.A2(n_19),
.B1(n_22),
.B2(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_0),
.A2(n_45),
.B1(n_46),
.B2(n_133),
.Y(n_241)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_5),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_5),
.A2(n_21),
.B1(n_64),
.B2(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_5),
.A2(n_21),
.B1(n_45),
.B2(n_46),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_7),
.A2(n_19),
.B1(n_22),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_7),
.A2(n_35),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_7),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_8),
.A2(n_40),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_8),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_19),
.B1(n_22),
.B2(n_40),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_8),
.A2(n_62),
.B(n_63),
.C(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_8),
.B(n_65),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_22),
.B(n_25),
.C(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_44),
.C(n_45),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_8),
.B(n_23),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_8),
.B(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_8),
.B(n_42),
.Y(n_257)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_112),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_111),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_15),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_15),
.B(n_300),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_15),
.B(n_300),
.Y(n_301)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_53),
.CI(n_80),
.CON(n_15),
.SN(n_15)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_16),
.A2(n_17),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_36),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_23),
.B(n_31),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_18),
.A2(n_73),
.B(n_74),
.Y(n_72)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_22),
.B1(n_25),
.B2(n_30),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_19),
.A2(n_22),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g189 ( 
.A1(n_22),
.A2(n_40),
.B(n_61),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_23),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_24),
.B(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_24),
.B(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_24),
.A2(n_32),
.B(n_102),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_24)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_27),
.A2(n_30),
.B(n_40),
.Y(n_212)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_28),
.B(n_229),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_31),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_31),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_32),
.B(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_48),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_37),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_38),
.A2(n_41),
.B(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_39),
.B(n_50),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_41),
.A2(n_49),
.B(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_42),
.B(n_216),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_45),
.B(n_253),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_49),
.B(n_226),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_50),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_70),
.B1(n_78),
.B2(n_79),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_54),
.A2(n_78),
.B1(n_97),
.B2(n_109),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_72),
.C(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_66),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_55),
.B(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_56),
.B(n_65),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_58),
.Y(n_135)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_59),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_59),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_65),
.B(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_66),
.B(n_131),
.Y(n_184)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_73),
.B(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_74),
.B(n_182),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_76),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_75),
.B(n_171),
.C(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_75),
.A2(n_76),
.B1(n_173),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_86),
.B(n_90),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_81),
.A2(n_87),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_81),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_81),
.B(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_81),
.A2(n_142),
.B1(n_211),
.B2(n_269),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_82),
.A2(n_147),
.B(n_148),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_82),
.B(n_85),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_82),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_125),
.Y(n_149)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_83),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_86),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_89),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_89),
.B(n_215),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_110),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_101),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_298),
.B(n_301),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_163),
.B(n_297),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_155),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_116),
.B(n_155),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_140),
.C(n_143),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_117),
.B(n_140),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_127),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_128),
.C(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_119),
.B(n_126),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_120),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_122),
.A2(n_124),
.B(n_147),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_124),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_136),
.B2(n_137),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_139),
.B(n_175),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_143),
.B(n_295),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_152),
.C(n_153),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_144),
.A2(n_145),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_150),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_149),
.B(n_239),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_151),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_152),
.A2(n_153),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_152),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_153),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_162),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_157),
.B(n_161),
.C(n_162),
.Y(n_300)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_292),
.B(n_296),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_204),
.B(n_278),
.C(n_291),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_192),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_166),
.B(n_192),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_179),
.B2(n_191),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_177),
.B2(n_178),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_169),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_169),
.B(n_178),
.C(n_191),
.Y(n_279)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_172),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_176),
.Y(n_183)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_181),
.B(n_186),
.C(n_187),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_184),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_190),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_198),
.C(n_199),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_194),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_202),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_203),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_277),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_220),
.B(n_276),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_207),
.B(n_217),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_213),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_210),
.B(n_213),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_211),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_271),
.B(n_275),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_262),
.B(n_270),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_243),
.B(n_261),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_224),
.B(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_242),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_233),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_236),
.C(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_234),
.Y(n_236)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_237),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_250),
.B(n_260),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_245),
.B(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_256),
.B(n_259),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_264),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_267),
.C(n_268),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_290),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_288),
.B2(n_289),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_289),
.C(n_290),
.Y(n_293)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);


endmodule