module fake_jpeg_3917_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_28),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_18),
.B1(n_26),
.B2(n_30),
.Y(n_56)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_49),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_48),
.B1(n_28),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_20),
.B1(n_18),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_37),
.B1(n_31),
.B2(n_27),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_23),
.B(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_66),
.B1(n_33),
.B2(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_0),
.Y(n_92)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_26),
.B1(n_23),
.B2(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_39),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_73),
.B1(n_79),
.B2(n_62),
.Y(n_109)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_85),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_81),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_38),
.B1(n_17),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_83),
.B1(n_87),
.B2(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_38),
.C(n_37),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_48),
.C(n_47),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_17),
.B1(n_34),
.B2(n_40),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_19),
.B(n_37),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_60),
.B(n_31),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_58),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_51),
.B1(n_41),
.B2(n_58),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_55),
.B(n_37),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_41),
.B(n_42),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_107),
.B1(n_109),
.B2(n_87),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_73),
.B(n_70),
.Y(n_120)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_98),
.Y(n_125)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_84),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_41),
.C(n_40),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_90),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_40),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_102),
.B(n_103),
.CI(n_83),
.CON(n_132),
.SN(n_132)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_42),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_114),
.B(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_71),
.A2(n_62),
.B1(n_51),
.B2(n_42),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_72),
.B1(n_75),
.B2(n_69),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_117),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_0),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_76),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_81),
.A2(n_31),
.B(n_27),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_87),
.A2(n_31),
.B1(n_27),
.B2(n_21),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_118),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_27),
.B1(n_21),
.B2(n_58),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_70),
.B(n_77),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_124),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_120),
.A2(n_92),
.B(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_129),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_127),
.B1(n_101),
.B2(n_110),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_85),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_113),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_72),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_139),
.B1(n_106),
.B2(n_97),
.Y(n_145)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_94),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_85),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_142),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_78),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_145),
.A2(n_171),
.B1(n_160),
.B2(n_151),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_162),
.C(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_144),
.B1(n_93),
.B2(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_143),
.B1(n_121),
.B2(n_122),
.Y(n_188)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_156),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_100),
.B1(n_114),
.B2(n_111),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_172),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_120),
.B(n_140),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_107),
.C(n_68),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_99),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_129),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_134),
.B(n_68),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_99),
.B1(n_86),
.B2(n_69),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_132),
.Y(n_172)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_133),
.B(n_131),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_186),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_131),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_170),
.B(n_167),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_154),
.B(n_132),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_194),
.C(n_146),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_138),
.B(n_121),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_192),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_80),
.B(n_86),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_191),
.A2(n_149),
.B1(n_153),
.B2(n_147),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_148),
.A2(n_86),
.B1(n_21),
.B2(n_14),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_169),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_165),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_195),
.Y(n_206)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_156),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_161),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.C(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_162),
.C(n_154),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_208),
.B(n_191),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_216),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_210),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_213),
.Y(n_224)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_150),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_190),
.B(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_207),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_211),
.B(n_178),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_220),
.C(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_178),
.C(n_203),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_228),
.Y(n_239)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_189),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_180),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_187),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_174),
.C(n_196),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_232),
.C(n_215),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_193),
.B(n_173),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_184),
.C(n_188),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_192),
.Y(n_233)
);

OAI22x1_ASAP7_75t_L g238 ( 
.A1(n_233),
.A2(n_216),
.B1(n_184),
.B2(n_198),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_240),
.C(n_221),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_206),
.B1(n_199),
.B2(n_212),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_2),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_224),
.B1(n_223),
.B2(n_222),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_204),
.C(n_198),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_233),
.A2(n_200),
.B1(n_215),
.B2(n_209),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_13),
.Y(n_250)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_223),
.B1(n_182),
.B2(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_176),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_252),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_250),
.B(n_3),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_13),
.C(n_2),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_1),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_1),
.C(n_2),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_255),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_258),
.B(n_259),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_262),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_234),
.B(n_243),
.Y(n_264)
);

AOI322xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_267),
.A3(n_257),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_242),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_265),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_266),
.B1(n_257),
.B2(n_265),
.Y(n_269)
);

O2A1O1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_271),
.B(n_272),
.C(n_7),
.Y(n_273)
);

O2A1O1Ixp33_ASAP7_75t_R g272 ( 
.A1(n_264),
.A2(n_4),
.B(n_6),
.C(n_7),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_274),
.C(n_10),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_10),
.C(n_11),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_10),
.CI(n_11),
.CON(n_276),
.SN(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_12),
.Y(n_277)
);


endmodule