module real_jpeg_20055_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_0),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_0),
.A2(n_29),
.B1(n_32),
.B2(n_46),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_29),
.B1(n_32),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_1),
.A2(n_37),
.B1(n_72),
.B2(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_37),
.B1(n_40),
.B2(n_45),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_2),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_2),
.A2(n_14),
.B(n_29),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_2),
.A2(n_40),
.B1(n_45),
.B2(n_98),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_28),
.B1(n_157),
.B2(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_2),
.B(n_73),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g188 ( 
.A1(n_2),
.A2(n_73),
.B(n_184),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_3),
.A2(n_69),
.B1(n_75),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_72),
.B1(n_73),
.B2(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_3),
.A2(n_29),
.B1(n_32),
.B2(n_78),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_3),
.A2(n_40),
.B1(n_45),
.B2(n_78),
.Y(n_192)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_69),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_5),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_72),
.B1(n_73),
.B2(n_76),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_5),
.A2(n_29),
.B1(n_32),
.B2(n_76),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_5),
.A2(n_40),
.B1(n_45),
.B2(n_76),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_6),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_33),
.B1(n_40),
.B2(n_45),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_33),
.B1(n_72),
.B2(n_73),
.Y(n_91)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_7),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_7),
.A2(n_27),
.B(n_101),
.Y(n_205)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_9),
.A2(n_40),
.B1(n_45),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_29),
.B1(n_32),
.B2(n_48),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_11),
.A2(n_69),
.B1(n_75),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_11),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_40),
.B1(n_45),
.B2(n_111),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_111),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_11),
.A2(n_72),
.B1(n_73),
.B2(n_111),
.Y(n_189)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_13),
.A2(n_68),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_40),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_14),
.A2(n_29),
.B1(n_32),
.B2(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_113),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_93),
.B2(n_112),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_49),
.B2(n_50),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_34),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_28),
.A2(n_59),
.B(n_60),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_28),
.A2(n_59),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_28),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_28),
.A2(n_102),
.B1(n_143),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_28),
.A2(n_34),
.B(n_145),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_31),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_32),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_35),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_140)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_35),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_36),
.A2(n_61),
.B(n_141),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_39),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_39),
.A2(n_42),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_39),
.A2(n_42),
.B1(n_153),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_39),
.A2(n_42),
.B1(n_175),
.B2(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_39),
.A2(n_192),
.B(n_212),
.Y(n_211)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_45),
.B1(n_84),
.B2(n_85),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_40),
.A2(n_72),
.A3(n_85),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_44),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_42),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_42),
.B(n_98),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_43),
.A2(n_45),
.B(n_98),
.C(n_149),
.Y(n_148)
);

NAND2xp33_ASAP7_75t_SL g185 ( 
.A(n_45),
.B(n_84),
.Y(n_185)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_62),
.B1(n_63),
.B2(n_92),
.Y(n_50)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_57),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_52),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_55),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_80),
.B2(n_81),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_74),
.B1(n_79),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_71),
.B1(n_97),
.B2(n_110),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.C(n_71),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_73),
.Y(n_96)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_98),
.CON(n_97),
.SN(n_97)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_72),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_84),
.B(n_86),
.C(n_87),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_79),
.B(n_98),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_88),
.B(n_90),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_104),
.B(n_106),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_83),
.A2(n_87),
.B1(n_105),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_83),
.A2(n_87),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_83),
.A2(n_87),
.B1(n_128),
.B2(n_189),
.Y(n_202)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_107),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_95),
.B(n_99),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_102),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_119),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_114),
.A2(n_115),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_118),
.B(n_119),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_129),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_123),
.B(n_125),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_129),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_230),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_225),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_214),
.B(n_224),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_197),
.B(n_213),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_178),
.B(n_196),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_166),
.B(n_177),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_154),
.B(n_165),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_146),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_150),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_159),
.B(n_164),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_158),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_168),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_174),
.C(n_176),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B1(n_194),
.B2(n_195),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_193),
.C(n_194),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_199),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_208),
.B2(n_209),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_210),
.C(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_204),
.C(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.C(n_222),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);


endmodule