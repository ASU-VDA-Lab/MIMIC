module fake_jpeg_28642_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_1),
.Y(n_51)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_40),
.B1(n_35),
.B2(n_37),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_35),
.B1(n_41),
.B2(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_43),
.B1(n_2),
.B2(n_4),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_66),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_83)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_6),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_8),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_85),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_73),
.Y(n_91)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_13),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_72),
.B(n_80),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_93),
.B(n_87),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_95),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_81),
.C(n_76),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_86),
.C(n_83),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_97),
.C(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_90),
.C(n_89),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_20),
.Y(n_103)
);

AOI211xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_21),
.B(n_22),
.C(n_24),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_105)
);

XNOR2x2_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_30),
.Y(n_106)
);


endmodule