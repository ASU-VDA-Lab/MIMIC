module fake_jpeg_17042_n_383 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_383);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_383;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_38),
.B(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_20),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_64),
.Y(n_75)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_58),
.Y(n_80)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_1),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_19),
.Y(n_101)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_24),
.B(n_1),
.Y(n_62)
);

OR2x4_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_32),
.Y(n_72)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_20),
.B(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_39),
.A2(n_22),
.B1(n_34),
.B2(n_17),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_74),
.B1(n_90),
.B2(n_96),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_71),
.B(n_83),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_99),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_84),
.B1(n_95),
.B2(n_10),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_46),
.B(n_29),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_86),
.B(n_114),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_29),
.B1(n_23),
.B2(n_31),
.Y(n_90)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_37),
.B1(n_26),
.B2(n_32),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_26),
.B1(n_37),
.B2(n_19),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_97),
.A2(n_98),
.B1(n_105),
.B2(n_109),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_52),
.A2(n_59),
.B1(n_61),
.B2(n_54),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_25),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_16),
.Y(n_102)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_115),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_48),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_30),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_48),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_110),
.A2(n_113),
.B1(n_82),
.B2(n_89),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_45),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_16),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g115 ( 
.A(n_55),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_72),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_143),
.B1(n_116),
.B2(n_117),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_73),
.Y(n_127)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_24),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_78),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_92),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_99),
.B(n_100),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_138),
.B(n_141),
.C(n_155),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_81),
.B(n_80),
.Y(n_141)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_88),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_146),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_105),
.A2(n_24),
.B(n_25),
.C(n_12),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_145),
.A2(n_153),
.B(n_160),
.C(n_142),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_92),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_147),
.B(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_87),
.B(n_75),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_100),
.A2(n_25),
.B(n_11),
.C(n_12),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_154),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_75),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_155),
.B(n_163),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_25),
.B1(n_11),
.B2(n_12),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_156),
.A2(n_157),
.B1(n_164),
.B2(n_165),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_10),
.B1(n_13),
.B2(n_25),
.Y(n_157)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_158),
.A2(n_160),
.B1(n_129),
.B2(n_151),
.Y(n_197)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_69),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_69),
.B(n_10),
.Y(n_161)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_13),
.Y(n_162)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_91),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_93),
.A2(n_108),
.B1(n_110),
.B2(n_107),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_79),
.A2(n_82),
.B1(n_89),
.B2(n_108),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_85),
.B1(n_67),
.B2(n_104),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_169),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_172),
.A2(n_173),
.B1(n_178),
.B2(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_138),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_193),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_175),
.A2(n_181),
.B1(n_182),
.B2(n_191),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_119),
.A2(n_143),
.B1(n_164),
.B2(n_118),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_180),
.A2(n_192),
.B1(n_198),
.B2(n_205),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_140),
.B1(n_138),
.B2(n_133),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_139),
.A2(n_145),
.B1(n_128),
.B2(n_131),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_141),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_216),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_153),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_124),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_190),
.Y(n_220)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_126),
.B(n_157),
.CI(n_123),
.CON(n_189),
.SN(n_189)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_189),
.B(n_210),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_121),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_152),
.B1(n_130),
.B2(n_166),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_159),
.B1(n_134),
.B2(n_135),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_SL g193 ( 
.A(n_134),
.B(n_135),
.C(n_169),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_194),
.A2(n_207),
.B(n_179),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_129),
.A2(n_144),
.B1(n_142),
.B2(n_148),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_204),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_136),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_132),
.A2(n_71),
.B1(n_72),
.B2(n_164),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_136),
.B(n_148),
.Y(n_207)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_138),
.B(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_189),
.Y(n_241)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_218),
.A2(n_244),
.B(n_233),
.Y(n_286)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_224),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_170),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_196),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_228),
.Y(n_265)
);

AO22x1_ASAP7_75t_SL g227 ( 
.A1(n_194),
.A2(n_178),
.B1(n_182),
.B2(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_227),
.A2(n_229),
.B1(n_234),
.B2(n_238),
.Y(n_275)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_179),
.A2(n_212),
.B1(n_173),
.B2(n_181),
.Y(n_229)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_232),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_183),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_233),
.B(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_174),
.A2(n_216),
.B1(n_175),
.B2(n_186),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_215),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_246),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_171),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_248),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_193),
.A2(n_189),
.B(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_204),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_199),
.B(n_191),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_249),
.B(n_255),
.Y(n_290)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_207),
.B(n_188),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_258),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_200),
.A2(n_203),
.B1(n_176),
.B2(n_207),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_254),
.A2(n_225),
.B1(n_253),
.B2(n_228),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_195),
.B(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_177),
.B(n_170),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_212),
.B(n_173),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_229),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_270),
.C(n_289),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_220),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_260),
.A2(n_283),
.B(n_285),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_262),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_235),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_268),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_251),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_249),
.B(n_220),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_280),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_258),
.C(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_231),
.B(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_278),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_279),
.A2(n_282),
.B1(n_272),
.B2(n_265),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_239),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_235),
.A2(n_231),
.B(n_219),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_218),
.A2(n_238),
.B(n_222),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_273),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_222),
.B(n_227),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_256),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_230),
.B(n_227),
.C(n_252),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_236),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_291),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_230),
.B(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_292),
.Y(n_313)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_274),
.Y(n_294)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_292),
.A2(n_232),
.B1(n_237),
.B2(n_221),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_295),
.A2(n_298),
.B1(n_315),
.B2(n_307),
.Y(n_331)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_278),
.A2(n_265),
.B(n_267),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_300),
.B(n_305),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_264),
.A2(n_279),
.B1(n_260),
.B2(n_287),
.Y(n_298)
);

FAx1_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_264),
.CI(n_285),
.CON(n_300),
.SN(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_302),
.B(n_303),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_304),
.B(n_277),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_314),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_260),
.B1(n_267),
.B2(n_263),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_289),
.A2(n_275),
.B1(n_263),
.B2(n_284),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_311),
.A2(n_307),
.B1(n_304),
.B2(n_310),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_270),
.C(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_312),
.B(n_299),
.C(n_298),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_271),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_269),
.A2(n_276),
.B1(n_273),
.B2(n_260),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_316),
.Y(n_326)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_281),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_317),
.Y(n_334)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_271),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_320),
.A2(n_329),
.B(n_338),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_290),
.B(n_276),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_321),
.A2(n_327),
.B(n_297),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_313),
.A2(n_290),
.B1(n_268),
.B2(n_280),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_323),
.B1(n_328),
.B2(n_332),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_313),
.A2(n_284),
.B1(n_283),
.B2(n_272),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_336),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_261),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_272),
.B1(n_261),
.B2(n_277),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_310),
.A2(n_266),
.B(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_309),
.B(n_293),
.Y(n_335)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_335),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_305),
.A2(n_300),
.B1(n_303),
.B2(n_309),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g351 ( 
.A1(n_337),
.A2(n_339),
.B(n_295),
.C(n_315),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_302),
.B1(n_297),
.B2(n_319),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_340),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_326),
.A2(n_317),
.B1(n_316),
.B2(n_318),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_345),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_299),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_322),
.Y(n_347)
);

INVx11_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_335),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_348),
.A2(n_350),
.B(n_351),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_349),
.A2(n_352),
.B1(n_334),
.B2(n_326),
.Y(n_356)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_325),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_312),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_354),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_356),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_355),
.A2(n_337),
.B1(n_342),
.B2(n_349),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_357),
.A2(n_361),
.B1(n_344),
.B2(n_351),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_323),
.C(n_328),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_364),
.C(n_365),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_320),
.C(n_331),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_330),
.C(n_334),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_366),
.B(n_367),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_343),
.C(n_355),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_343),
.C(n_344),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_370),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_346),
.C(n_341),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_365),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_375),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_369),
.B(n_362),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_374),
.Y(n_376)
);

OAI21x1_ASAP7_75t_L g378 ( 
.A1(n_376),
.A2(n_372),
.B(n_360),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_378),
.Y(n_379)
);

OAI21x1_ASAP7_75t_SL g380 ( 
.A1(n_379),
.A2(n_377),
.B(n_373),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_359),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_381),
.A2(n_360),
.B(n_362),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_356),
.Y(n_383)
);


endmodule