module fake_jpeg_31803_n_33 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_33);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_33;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_6),
.A2(n_1),
.B1(n_9),
.B2(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

AOI21xp33_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_0),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_19),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_3),
.Y(n_21)
);

NAND3xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_17),
.C(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_19),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_26),
.B(n_14),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_17),
.B1(n_14),
.B2(n_12),
.Y(n_25)
);

A2O1A1O1Ixp25_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_16),
.B(n_5),
.C(n_7),
.D(n_8),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_22),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_23),
.A3(n_30),
.B1(n_25),
.B2(n_4),
.C1(n_10),
.C2(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_33)
);


endmodule