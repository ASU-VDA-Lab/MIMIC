module fake_jpeg_29714_n_283 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx24_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_17),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_43),
.Y(n_80)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_0),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_48),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

CKINVDCx6p67_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_28),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_33),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_25),
.B(n_0),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx2_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_63),
.Y(n_122)
);

NAND2x1_ASAP7_75t_SL g64 ( 
.A(n_52),
.B(n_39),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_66),
.Y(n_132)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_79),
.Y(n_105)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_19),
.B1(n_38),
.B2(n_37),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_81),
.B1(n_32),
.B2(n_23),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_39),
.B1(n_28),
.B2(n_29),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_100),
.B1(n_103),
.B2(n_32),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_29),
.C(n_31),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_36),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_24),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_86),
.B(n_23),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_42),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_45),
.B(n_20),
.CON(n_92),
.SN(n_92)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_24),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_98),
.Y(n_117)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_36),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_44),
.A2(n_1),
.B(n_2),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_1),
.C(n_2),
.Y(n_112)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_24),
.B1(n_20),
.B2(n_35),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_48),
.C(n_47),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_106),
.B(n_109),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_99),
.B1(n_89),
.B2(n_68),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_134),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_46),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_114),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_76),
.B(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_66),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_59),
.B1(n_20),
.B2(n_3),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_63),
.B1(n_64),
.B2(n_90),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_75),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_108),
.B1(n_131),
.B2(n_117),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_80),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_17),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_80),
.B(n_65),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g194 ( 
.A1(n_137),
.A2(n_127),
.B(n_9),
.Y(n_194)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

AO22x2_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_90),
.B1(n_62),
.B2(n_72),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g191 ( 
.A1(n_139),
.A2(n_149),
.B(n_154),
.C(n_144),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_91),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_141),
.B(n_145),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_62),
.B1(n_72),
.B2(n_103),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_160),
.B1(n_104),
.B2(n_124),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_74),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_147),
.A2(n_153),
.B1(n_154),
.B2(n_157),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_111),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_116),
.A2(n_90),
.B(n_74),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_119),
.B(n_111),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_163),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_109),
.A2(n_89),
.B1(n_82),
.B2(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_87),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_155),
.B(n_161),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_82),
.B1(n_83),
.B2(n_66),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_83),
.B1(n_6),
.B2(n_7),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_5),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_106),
.B(n_6),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_118),
.B(n_15),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_8),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_176),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_175),
.B(n_180),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_174),
.B(n_181),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_119),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_132),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_189),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_159),
.A2(n_115),
.B1(n_107),
.B2(n_125),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_SL g180 ( 
.A(n_158),
.B(n_104),
.C(n_9),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_107),
.B(n_115),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_182),
.B(n_183),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_124),
.B(n_104),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_194),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_129),
.B1(n_127),
.B2(n_10),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_136),
.B(n_129),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_127),
.B1(n_9),
.B2(n_12),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_192),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_209),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_169),
.A2(n_137),
.B1(n_147),
.B2(n_139),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_181),
.B1(n_191),
.B2(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_157),
.A3(n_160),
.B1(n_158),
.B2(n_148),
.C1(n_142),
.C2(n_139),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_215),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_142),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_139),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_210),
.B(n_214),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_139),
.C(n_151),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_172),
.C(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_212),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_151),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_182),
.B(n_152),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_168),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_218),
.B(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_197),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_230),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_211),
.B(n_215),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_210),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_190),
.B1(n_185),
.B2(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_193),
.B(n_183),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_194),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_233),
.C(n_225),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_193),
.C(n_191),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_226),
.B(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_237),
.A2(n_240),
.B1(n_232),
.B2(n_196),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_197),
.B1(n_202),
.B2(n_200),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_198),
.C(n_213),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_246),
.C(n_230),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_204),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_214),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_247),
.B(n_252),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_244),
.A2(n_219),
.B1(n_233),
.B2(n_191),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_257),
.B1(n_240),
.B2(n_235),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_235),
.B1(n_216),
.B2(n_246),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_217),
.B(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_251),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_256),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.C(n_236),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_224),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_223),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_237),
.A2(n_208),
.B1(n_216),
.B2(n_195),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_263),
.A3(n_258),
.B1(n_262),
.B2(n_260),
.C1(n_251),
.C2(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_265),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_243),
.B1(n_195),
.B2(n_201),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_255),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_236),
.C(n_207),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_270),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_268),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_271),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_248),
.B(n_206),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_170),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_266),
.B(n_264),
.C(n_265),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_171),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_270),
.A2(n_212),
.B(n_171),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_276),
.A2(n_187),
.B(n_186),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_278),
.B1(n_276),
.B2(n_164),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_272),
.C(n_275),
.Y(n_280)
);

OAI221xp5_ASAP7_75t_SL g282 ( 
.A1(n_280),
.A2(n_281),
.B1(n_138),
.B2(n_13),
.C(n_14),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_8),
.C(n_15),
.Y(n_283)
);


endmodule