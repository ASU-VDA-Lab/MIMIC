module fake_aes_3514_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
NOR2xp33_ASAP7_75t_R g11 ( .A(n_7), .B(n_1), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_8), .B(n_2), .Y(n_13) );
INVxp33_ASAP7_75t_SL g14 ( .A(n_2), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_15), .B(n_0), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_12), .B(n_0), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_10), .B(n_3), .Y(n_18) );
INVxp67_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
OAI21x1_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_15), .B(n_13), .Y(n_20) );
BUFx3_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NAND3xp33_ASAP7_75t_L g24 ( .A(n_21), .B(n_19), .C(n_18), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_22), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
NOR2xp33_ASAP7_75t_L g28 ( .A(n_26), .B(n_14), .Y(n_28) );
NOR3xp33_ASAP7_75t_L g29 ( .A(n_28), .B(n_14), .C(n_26), .Y(n_29) );
INVx3_ASAP7_75t_SL g30 ( .A(n_27), .Y(n_30) );
INVx2_ASAP7_75t_SL g31 ( .A(n_27), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_30), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AOI322xp5_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_33), .A3(n_29), .B1(n_11), .B2(n_3), .C1(n_5), .C2(n_4), .Y(n_35) );
endmodule