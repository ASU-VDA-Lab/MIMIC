module fake_jpeg_23954_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_46),
.Y(n_62)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_45),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_8),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_0),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_32),
.B1(n_27),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_59),
.B1(n_21),
.B2(n_34),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_30),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_29),
.B1(n_38),
.B2(n_37),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_57),
.A2(n_64),
.B(n_75),
.Y(n_113)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_32),
.B1(n_27),
.B2(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_68),
.Y(n_100)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_79),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_20),
.B1(n_38),
.B2(n_32),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g97 ( 
.A(n_72),
.B(n_80),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_38),
.B1(n_18),
.B2(n_20),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_25),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_18),
.B1(n_24),
.B2(n_33),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_83),
.B1(n_31),
.B2(n_35),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_24),
.B1(n_34),
.B2(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_2),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_54),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_85),
.B(n_91),
.Y(n_156)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_86),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_65),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_87),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_39),
.B(n_46),
.C(n_47),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_88),
.A2(n_98),
.B(n_11),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_48),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_47),
.C(n_43),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_43),
.C(n_74),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_96),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_35),
.B(n_28),
.C(n_43),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_101),
.B1(n_109),
.B2(n_114),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_28),
.B1(n_24),
.B2(n_31),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_116),
.B1(n_119),
.B2(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_69),
.B1(n_52),
.B2(n_66),
.Y(n_139)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_43),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_82),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_115),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_80),
.B(n_21),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_22),
.B1(n_26),
.B2(n_23),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_122),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_23),
.C(n_26),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_138),
.B(n_152),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_70),
.B1(n_73),
.B2(n_69),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_125),
.A2(n_139),
.B1(n_140),
.B2(n_151),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_126),
.B(n_92),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_90),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_58),
.B1(n_63),
.B2(n_67),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_137),
.B1(n_99),
.B2(n_114),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_142),
.C(n_143),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_62),
.B(n_23),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_89),
.B(n_103),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_95),
.B1(n_113),
.B2(n_100),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_2),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_93),
.A2(n_52),
.B1(n_26),
.B2(n_22),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_76),
.C(n_23),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_23),
.C(n_22),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_26),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_89),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_93),
.A2(n_22),
.B1(n_11),
.B2(n_4),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_96),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_96),
.B(n_115),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_96),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

OAI32xp33_ASAP7_75t_L g155 ( 
.A1(n_98),
.A2(n_12),
.A3(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_15),
.Y(n_177)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_160),
.A2(n_164),
.B(n_187),
.Y(n_206)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_163),
.B(n_170),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_167),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_178),
.B1(n_136),
.B2(n_123),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_103),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_173),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_105),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_130),
.Y(n_174)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_177),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_137),
.A2(n_108),
.B1(n_86),
.B2(n_92),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_182),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_106),
.C(n_87),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_136),
.C(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_2),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_189),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_3),
.B(n_5),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_152),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_138),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g190 ( 
.A(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_155),
.B1(n_141),
.B2(n_129),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_192),
.A2(n_208),
.B1(n_209),
.B2(n_214),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_212),
.C(n_165),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_195),
.A2(n_196),
.B1(n_204),
.B2(n_218),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_175),
.B1(n_179),
.B2(n_178),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_132),
.B1(n_144),
.B2(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_211),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_132),
.B1(n_148),
.B2(n_123),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_133),
.B1(n_118),
.B2(n_150),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_180),
.C(n_173),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_215),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_133),
.B1(n_118),
.B2(n_149),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_133),
.B(n_3),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_216),
.A2(n_220),
.B(n_182),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_104),
.B1(n_3),
.B2(n_10),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_164),
.B(n_6),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_183),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_183),
.B1(n_159),
.B2(n_166),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_216),
.B(n_217),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_225),
.B(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_232),
.C(n_235),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_184),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_238),
.Y(n_262)
);

HB1xp67_ASAP7_75t_SL g260 ( 
.A(n_231),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_158),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_206),
.A2(n_158),
.B(n_170),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_159),
.C(n_191),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_198),
.A2(n_177),
.B1(n_185),
.B2(n_166),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_197),
.A2(n_171),
.B(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_241),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_104),
.B(n_12),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_198),
.A2(n_217),
.B1(n_201),
.B2(n_192),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_196),
.B1(n_195),
.B2(n_218),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_213),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_199),
.A2(n_6),
.B1(n_13),
.B2(n_14),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_247),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_215),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_250),
.A2(n_229),
.B1(n_236),
.B2(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_232),
.B(n_193),
.C(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_235),
.C(n_237),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_214),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_231),
.Y(n_280)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_245),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_261),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_220),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_223),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_227),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_266),
.B(n_234),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_285),
.B1(n_249),
.B2(n_254),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_242),
.B1(n_224),
.B2(n_205),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_274),
.B1(n_278),
.B2(n_284),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_277),
.C(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_242),
.B1(n_229),
.B2(n_233),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_259),
.B(n_211),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_248),
.B(n_251),
.C(n_260),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_194),
.B1(n_219),
.B2(n_228),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_283),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_210),
.C(n_225),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_252),
.C(n_220),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_255),
.B(n_250),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_225),
.B1(n_230),
.B2(n_202),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_209),
.B1(n_230),
.B2(n_226),
.Y(n_285)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_284),
.A2(n_258),
.B(n_253),
.C(n_264),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_294),
.B(n_275),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_258),
.B1(n_267),
.B2(n_257),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_290),
.A2(n_298),
.B1(n_273),
.B2(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_230),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_295),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_283),
.A2(n_264),
.B(n_267),
.C(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_202),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_265),
.B(n_261),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_269),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_277),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_271),
.A2(n_252),
.B1(n_14),
.B2(n_15),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_272),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_200),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_13),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_13),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_289),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_294),
.C(n_289),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_299),
.B1(n_291),
.B2(n_294),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_287),
.B1(n_294),
.B2(n_289),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_292),
.C(n_297),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_318),
.B(n_319),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_308),
.B(n_299),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_314),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_322),
.B(n_315),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_321),
.C(n_317),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_328),
.A2(n_323),
.B(n_326),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_317),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_310),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_16),
.Y(n_332)
);


endmodule