module fake_jpeg_17933_n_343 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_343);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_343;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_48),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_0),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_23),
.B1(n_31),
.B2(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_55),
.B(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_20),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_31),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_23),
.B1(n_19),
.B2(n_26),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_90),
.Y(n_125)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_82),
.B(n_99),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_30),
.B(n_34),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_22),
.B(n_23),
.C(n_29),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_48),
.C(n_45),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_88),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_53),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_103),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_45),
.C(n_43),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_38),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_95),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_54),
.B(n_52),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_22),
.B(n_32),
.Y(n_115)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_35),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_53),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_104),
.Y(n_126)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_60),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_60),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_36),
.C(n_54),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_130),
.C(n_45),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_115),
.A2(n_119),
.B(n_124),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_83),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_137),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_70),
.B1(n_61),
.B2(n_40),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_128),
.B1(n_140),
.B2(n_78),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_24),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_70),
.B1(n_40),
.B2(n_50),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_93),
.A2(n_80),
.B(n_76),
.Y(n_130)
);

BUFx24_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_80),
.A2(n_50),
.B1(n_24),
.B2(n_37),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_103),
.B1(n_78),
.B2(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_101),
.B1(n_19),
.B2(n_26),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_92),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_143),
.B(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_88),
.B(n_27),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_124),
.B(n_129),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_146),
.A2(n_152),
.B1(n_120),
.B2(n_117),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_126),
.A2(n_108),
.B1(n_102),
.B2(n_77),
.Y(n_147)
);

OAI22x1_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_97),
.B1(n_135),
.B2(n_136),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_151),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_24),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_137),
.B(n_112),
.C(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_105),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_96),
.B1(n_105),
.B2(n_83),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_142),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_104),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_139),
.C(n_127),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_132),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_160),
.A2(n_112),
.B(n_125),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_170),
.B1(n_185),
.B2(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_177),
.C(n_181),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_172),
.B(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_114),
.B1(n_120),
.B2(n_124),
.Y(n_170)
);

XOR2x1_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_143),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_113),
.B(n_125),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_150),
.A2(n_113),
.B(n_140),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_179),
.B(n_180),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_121),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_126),
.B(n_120),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_139),
.B1(n_136),
.B2(n_106),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_127),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_186),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_162),
.A2(n_116),
.B(n_122),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_147),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_151),
.A2(n_152),
.B1(n_144),
.B2(n_149),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_156),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_79),
.B1(n_98),
.B2(n_33),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_26),
.B1(n_19),
.B2(n_165),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_213),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_158),
.C(n_154),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_206),
.C(n_212),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_198),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_182),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_208),
.B(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_205),
.A2(n_207),
.B1(n_22),
.B2(n_38),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_161),
.C(n_164),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_19),
.B1(n_141),
.B2(n_21),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_45),
.C(n_135),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_43),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_220),
.C(n_173),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_170),
.A2(n_84),
.B1(n_81),
.B2(n_51),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_219),
.A2(n_221),
.B1(n_190),
.B2(n_178),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_51),
.C(n_44),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_33),
.B1(n_32),
.B2(n_29),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_18),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_223),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_236),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_228),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_185),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_241),
.C(n_247),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_198),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_172),
.B(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_233),
.A2(n_239),
.B1(n_242),
.B2(n_244),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_209),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_202),
.A2(n_178),
.B1(n_190),
.B2(n_187),
.Y(n_239)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_188),
.B1(n_179),
.B2(n_168),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_171),
.B(n_192),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_246),
.B(n_195),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_134),
.C(n_123),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_134),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_252),
.B(n_15),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_223),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_206),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_257),
.C(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_204),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_211),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_202),
.B1(n_218),
.B2(n_208),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_262),
.B1(n_271),
.B2(n_38),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_234),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_261),
.B(n_268),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_212),
.B1(n_219),
.B2(n_210),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_221),
.C(n_134),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_269),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_34),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_267),
.C(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_123),
.C(n_30),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_123),
.C(n_30),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_15),
.B1(n_16),
.B2(n_13),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_269),
.A2(n_233),
.B(n_245),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_272),
.A2(n_273),
.B(n_275),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_249),
.A2(n_242),
.B(n_238),
.C(n_232),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_265),
.A2(n_224),
.B(n_244),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_240),
.B1(n_247),
.B2(n_37),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_281),
.B1(n_289),
.B2(n_35),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_277),
.B(n_288),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_281)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

INVx11_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

AO221x1_ASAP7_75t_L g284 ( 
.A1(n_263),
.A2(n_18),
.B1(n_30),
.B2(n_34),
.C(n_25),
.Y(n_284)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_25),
.C(n_18),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_255),
.C(n_25),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_20),
.B(n_35),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_255),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_266),
.B(n_257),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_291),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_294),
.C(n_287),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_293),
.A2(n_274),
.B(n_273),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_18),
.C(n_25),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_299),
.C(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_285),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_34),
.C(n_28),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_28),
.C(n_21),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_28),
.B1(n_21),
.B2(n_20),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_285),
.B1(n_279),
.B2(n_281),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_11),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_272),
.B(n_275),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_309),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_312),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_305),
.A2(n_273),
.B(n_279),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_316),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_296),
.A2(n_273),
.B1(n_290),
.B2(n_282),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_294),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_289),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_315),
.A2(n_300),
.B(n_296),
.Y(n_317)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_317),
.B(n_324),
.C(n_306),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_314),
.A2(n_295),
.B(n_301),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_318),
.B(n_323),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_311),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_302),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_316),
.A2(n_299),
.B(n_8),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_326),
.A2(n_329),
.B(n_322),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_320),
.C(n_6),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_313),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_328),
.B(n_330),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g329 ( 
.A1(n_320),
.A2(n_8),
.B(n_11),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_319),
.B(n_6),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_332),
.A2(n_6),
.B(n_10),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_333),
.A2(n_334),
.B(n_335),
.Y(n_338)
);

AOI31xp33_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_5),
.A3(n_9),
.B(n_10),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_5),
.B(n_9),
.C(n_3),
.D(n_1),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_337),
.C(n_9),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_338),
.C(n_2),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_1),
.B(n_2),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_3),
.B1(n_37),
.B2(n_309),
.Y(n_343)
);


endmodule