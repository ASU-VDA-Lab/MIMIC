module fake_jpeg_24739_n_108 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_20),
.B(n_21),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_18),
.B1(n_16),
.B2(n_15),
.Y(n_31)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_10),
.B1(n_12),
.B2(n_22),
.Y(n_33)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_39),
.Y(n_49)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_23),
.B1(n_20),
.B2(n_14),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_28),
.B2(n_33),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_20),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_17),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_41),
.B1(n_40),
.B2(n_29),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_40),
.B(n_27),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_44),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_61),
.B(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_59),
.B(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_44),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_56),
.B(n_52),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_66),
.B(n_36),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_48),
.C(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_73),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_44),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_38),
.B1(n_35),
.B2(n_32),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_63),
.B(n_55),
.Y(n_71)
);

XNOR2x1_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_19),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_72),
.A2(n_64),
.B1(n_38),
.B2(n_57),
.Y(n_77)
);

AO21x1_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_18),
.B(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_69),
.B1(n_74),
.B2(n_67),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_77),
.A2(n_82),
.B(n_76),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_64),
.B1(n_62),
.B2(n_14),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_17),
.B1(n_19),
.B2(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_81),
.B(n_1),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_89),
.B(n_79),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_19),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_87),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_2),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_81),
.B(n_78),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_83),
.B(n_80),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_77),
.B1(n_92),
.B2(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_2),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_87),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_3),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_96),
.B(n_99),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_103),
.A2(n_3),
.B(n_4),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_104),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_4),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_5),
.B(n_6),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_7),
.Y(n_108)
);


endmodule