module real_jpeg_33846_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_0),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_0),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_0),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_1),
.A2(n_269),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_1),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_1),
.A2(n_272),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_L g427 ( 
.A1(n_1),
.A2(n_272),
.B1(n_428),
.B2(n_430),
.Y(n_427)
);

OAI22xp33_ASAP7_75t_SL g459 ( 
.A1(n_1),
.A2(n_272),
.B1(n_460),
.B2(n_462),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_2),
.B(n_529),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_2),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_3),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_3),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_3),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_5),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_5),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_115),
.B1(n_121),
.B2(n_122),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_6),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_6),
.A2(n_121),
.B1(n_169),
.B2(n_173),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_6),
.A2(n_121),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_6),
.A2(n_121),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_7),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_8),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_8),
.A2(n_49),
.B1(n_104),
.B2(n_108),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_49),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_8),
.B(n_154),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g419 ( 
.A(n_8),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_8),
.B(n_25),
.Y(n_455)
);

OAI32xp33_ASAP7_75t_L g471 ( 
.A1(n_8),
.A2(n_472),
.A3(n_474),
.B1(n_475),
.B2(n_481),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_9),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_10),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_10),
.Y(n_134)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_11),
.Y(n_487)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_12),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_13),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_13),
.A2(n_57),
.B1(n_123),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_13),
.A2(n_57),
.B1(n_221),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_13),
.A2(n_57),
.B1(n_207),
.B2(n_259),
.Y(n_258)
);

OAI321xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_190),
.A3(n_528),
.B1(n_530),
.B2(n_531),
.C(n_533),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_15),
.B(n_532),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_189),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_179),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_18),
.B(n_179),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_151),
.C(n_163),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_19),
.A2(n_151),
.B1(n_165),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_19),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_112),
.B1(n_113),
.B2(n_150),
.Y(n_19)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_20),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_77),
.B2(n_111),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_22),
.Y(n_188)
);

NOR2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_24),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_25),
.B(n_52),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_25),
.A2(n_50),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_25),
.B(n_327),
.Y(n_369)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AO21x1_ASAP7_75t_L g184 ( 
.A1(n_26),
.A2(n_40),
.B(n_63),
.Y(n_184)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AO21x2_ASAP7_75t_L g63 ( 
.A1(n_27),
.A2(n_64),
.B(n_71),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_28),
.A2(n_94),
.B1(n_98),
.B2(n_101),
.Y(n_93)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_30),
.Y(n_429)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_38),
.Y(n_223)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2x1_ASAP7_75t_L g265 ( 
.A(n_40),
.B(n_63),
.Y(n_265)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AO22x2_ASAP7_75t_L g126 ( 
.A1(n_47),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_126)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_48),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_49),
.A2(n_157),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_49),
.B(n_160),
.Y(n_159)
);

AOI32xp33_ASAP7_75t_L g414 ( 
.A1(n_49),
.A2(n_415),
.A3(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_49),
.B(n_476),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_49),
.B(n_503),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_49),
.B(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_51),
.B(n_369),
.Y(n_368)
);

NAND2x1_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_54),
.Y(n_340)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_62),
.B(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_65),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_65),
.Y(n_417)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_67),
.Y(n_172)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_71),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_77),
.B(n_165),
.C(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_R g187 ( 
.A(n_77),
.B(n_112),
.C(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_77),
.A2(n_111),
.B1(n_167),
.B2(n_197),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_77),
.B(n_368),
.C(n_370),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_77),
.A2(n_111),
.B1(n_368),
.B2(n_380),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_92),
.B(n_103),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_78),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_78),
.B(n_103),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_78),
.B(n_220),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_78),
.B(n_427),
.Y(n_440)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_93),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_79),
.Y(n_503)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_85),
.Y(n_461)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_85),
.Y(n_464)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_88),
.Y(n_305)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_91),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_92),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_92),
.B(n_228),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_92),
.B(n_103),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_92),
.B(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_107),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_107),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_107),
.Y(n_432)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_110),
.Y(n_424)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_125),
.B(n_135),
.Y(n_113)
);

OAI21x1_ASAP7_75t_SL g181 ( 
.A1(n_114),
.A2(n_152),
.B(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_120),
.Y(n_347)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_125),
.B(n_182),
.Y(n_236)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2x1p5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_126),
.B(n_268),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_128),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_128),
.Y(n_352)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_130),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_136),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_139),
.A2(n_143),
.B1(n_145),
.B2(n_148),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_140),
.Y(n_271)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_140),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_141),
.B(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_151),
.A2(n_165),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_153),
.B(n_267),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_154),
.B(n_156),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_155),
.B(n_311),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_156),
.B(n_236),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_159),
.Y(n_357)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_164),
.B(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_176),
.B(n_177),
.Y(n_167)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_177),
.B(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_178),
.B(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_181),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g317 ( 
.A(n_184),
.B(n_310),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_185),
.B(n_298),
.C(n_310),
.Y(n_297)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_190),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_285),
.B(n_524),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_244),
.B1(n_248),
.B2(n_281),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2x1_ASAP7_75t_L g525 ( 
.A(n_193),
.B(n_245),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_193),
.B(n_245),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.C(n_237),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_194),
.A2(n_237),
.B1(n_238),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_198),
.B(n_283),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_217),
.B(n_234),
.Y(n_198)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_199),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_199),
.B(n_235),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_199),
.A2(n_218),
.B1(n_233),
.B2(n_296),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_199),
.B(n_414),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_199),
.A2(n_233),
.B1(n_414),
.B2(n_446),
.Y(n_445)
);

AO21x2_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_203),
.B(n_210),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_200),
.A2(n_257),
.B(n_303),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_202),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_203),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_204),
.B(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_204),
.B(n_211),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_204),
.B(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx8_ASAP7_75t_L g498 ( 
.A(n_206),
.Y(n_498)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_207),
.Y(n_473)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_255),
.Y(n_254)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_217),
.B(n_280),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_233),
.Y(n_217)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_218),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_226),
.B(n_227),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_223),
.Y(n_474)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_227),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_227),
.B(n_426),
.Y(n_453)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

XOR2x2_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_241),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_242),
.B(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_243),
.B(n_252),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_243),
.B(n_440),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_249),
.B(n_282),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_277),
.C(n_278),
.Y(n_249)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_250),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.C(n_266),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_251),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_253),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g457 ( 
.A(n_254),
.B(n_458),
.Y(n_457)
);

BUFx4f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_257),
.B(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_265),
.Y(n_443)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

NAND2x1_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_277),
.B(n_279),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2x1p5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_405),
.Y(n_285)
);

OAI21x1_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_358),
.B(n_399),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_313),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_297),
.B2(n_312),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_290),
.B(n_297),
.Y(n_398)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_291),
.B(n_312),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_292),
.B(n_295),
.C(n_297),
.Y(n_401)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22x1_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_299),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_301),
.B(n_440),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_306),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_306),
.B(n_458),
.Y(n_504)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

AOI21x1_ASAP7_75t_L g396 ( 
.A1(n_313),
.A2(n_397),
.B(n_398),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.C(n_322),
.Y(n_313)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_320),
.Y(n_362)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_333),
.B(n_335),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_324),
.A2(n_334),
.B(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_325),
.A2(n_333),
.B1(n_334),
.B2(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_325),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_337),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

HAxp5_ASAP7_75t_SL g392 ( 
.A(n_338),
.B(n_339),
.CON(n_392),
.SN(n_392)
);

OAI31xp33_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_341),
.A3(n_344),
.B(n_348),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_353),
.B(n_357),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_374),
.B(n_396),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

NAND2x1p5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_363),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.C(n_371),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_372),
.Y(n_395)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_368),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_369),
.B(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_375),
.B(n_522),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_394),
.Y(n_376)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_377),
.B(n_394),
.Y(n_522)
);

OAI21xp33_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_381),
.B(n_393),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_378),
.B(n_434),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_391),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_382),
.B(n_391),
.Y(n_393)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_383),
.B(n_392),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.C(n_387),
.Y(n_383)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_385),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.Y(n_411)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NOR2x1_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_389),
.Y(n_507)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_392),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_396),
.B(n_400),
.C(n_521),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_401),
.B(n_402),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_520),
.B(n_523),
.Y(n_405)
);

AO21x1_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_435),
.B(n_519),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_433),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_408),
.B(n_433),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_412),
.C(n_425),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_409),
.B(n_448),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_425),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_449),
.B(n_518),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_447),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_447),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_441),
.C(n_444),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_438),
.A2(n_439),
.B1(n_441),
.B2(n_442),
.Y(n_466)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_466),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_467),
.B(n_517),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_465),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_465),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_454),
.C(n_456),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_453),
.A2(n_454),
.B1(n_455),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_457),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_497),
.Y(n_496)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx12f_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_468),
.A2(n_493),
.B(n_516),
.Y(n_467)
);

NOR2x1_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_490),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_469),
.B(n_490),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_488),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_470),
.A2(n_471),
.B1(n_488),
.B2(n_489),
.Y(n_499)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_472),
.Y(n_509)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx4_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_494),
.A2(n_500),
.B(n_515),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_499),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_SL g515 ( 
.A(n_495),
.B(n_499),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_507),
.Y(n_506)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_501),
.A2(n_505),
.B(n_514),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_504),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_504),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_508),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_510),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_525),
.A2(n_526),
.B(n_527),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_528),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_534),
.Y(n_533)
);


endmodule