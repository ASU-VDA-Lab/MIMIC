module fake_jpeg_8926_n_78 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_46),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_54),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_41),
.B1(n_38),
.B2(n_20),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_31),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_30),
.B1(n_15),
.B2(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_13),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_17),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g67 ( 
.A1(n_61),
.A2(n_63),
.A3(n_64),
.B1(n_24),
.B2(n_25),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_59),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_65),
.C(n_66),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_56),
.C(n_69),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_57),
.C(n_58),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_26),
.B(n_27),
.C(n_63),
.D(n_68),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_62),
.Y(n_78)
);


endmodule