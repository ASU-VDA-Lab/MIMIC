module fake_jpeg_21886_n_107 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_107);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_107;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_23),
.Y(n_32)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_25),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_31),
.B1(n_25),
.B2(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_21),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_11),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_23),
.B(n_21),
.C(n_24),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_42),
.B1(n_28),
.B2(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_21),
.C(n_24),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_32),
.Y(n_47)
);

AOI32xp33_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_32),
.A3(n_28),
.B1(n_30),
.B2(n_14),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_38),
.B(n_3),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_50),
.B1(n_43),
.B2(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_51),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_13),
.B1(n_18),
.B2(n_9),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_18),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_55),
.B(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_2),
.C(n_5),
.Y(n_74)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_44),
.A3(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

OAI21x1_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_58),
.B(n_65),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_59),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_81),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_55),
.B1(n_56),
.B2(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

A2O1A1O1Ixp25_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_67),
.B(n_66),
.C(n_68),
.D(n_75),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_76),
.B(n_69),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_85),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_77),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_81),
.B1(n_78),
.B2(n_60),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_53),
.C(n_57),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_36),
.C(n_5),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_6),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_97),
.C(n_6),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_2),
.B(n_5),
.Y(n_97)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_101),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_6),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_103),
.C(n_7),
.Y(n_105)
);

BUFx24_ASAP7_75t_SL g106 ( 
.A(n_105),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_7),
.Y(n_107)
);


endmodule