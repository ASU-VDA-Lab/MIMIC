module fake_jpeg_12370_n_192 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_192);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_32),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_4),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_87),
.Y(n_98)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_52),
.B(n_1),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_52),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_103),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_69),
.B1(n_78),
.B2(n_59),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_61),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_78),
.B1(n_69),
.B2(n_76),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_60),
.B1(n_68),
.B2(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_117),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_121),
.B1(n_129),
.B2(n_2),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_118),
.Y(n_135)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_64),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_63),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_123),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_86),
.B1(n_75),
.B2(n_79),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_94),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_72),
.A3(n_56),
.B1(n_80),
.B2(n_71),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_8),
.Y(n_150)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_60),
.B1(n_68),
.B2(n_77),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_127),
.A2(n_81),
.B1(n_74),
.B2(n_66),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_17),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_53),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_2),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_134),
.B1(n_143),
.B2(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_62),
.B1(n_57),
.B2(n_82),
.Y(n_134)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_18),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_150),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_3),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_11),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_114),
.B(n_21),
.Y(n_149)
);

AO22x2_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_24),
.B1(n_46),
.B2(n_43),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_151),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_9),
.B(n_10),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_158),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_20),
.C(n_12),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_167),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_164),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_166),
.B(n_145),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_29),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_152),
.B1(n_141),
.B2(n_151),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_178),
.B(n_163),
.Y(n_180)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_145),
.B(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_160),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_149),
.B(n_13),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_179),
.A2(n_180),
.B(n_182),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_155),
.B(n_161),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_176),
.C(n_173),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_165),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_157),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_184),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_172),
.B(n_162),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_162),
.A3(n_169),
.B1(n_155),
.B2(n_11),
.C1(n_19),
.C2(n_31),
.Y(n_190)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.C(n_33),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_34),
.Y(n_192)
);


endmodule