module real_jpeg_8712_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_1),
.A2(n_42),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_1),
.A2(n_10),
.B1(n_42),
.B2(n_65),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_22),
.B1(n_26),
.B2(n_42),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_2),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_2),
.A2(n_9),
.B(n_57),
.Y(n_88)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_5),
.A2(n_22),
.B1(n_26),
.B2(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_38),
.B(n_44),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_5),
.B(n_38),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_5),
.A2(n_9),
.B(n_22),
.Y(n_116)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_8),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_9),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_9),
.A2(n_33),
.B1(n_57),
.B2(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_9),
.A2(n_10),
.B1(n_33),
.B2(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_9),
.B(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_9),
.B(n_52),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_9),
.A2(n_54),
.B(n_58),
.C(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_10),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_67),
.B(n_68),
.C(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_68),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_33),
.B(n_68),
.C(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_107),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_105),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_14),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_15),
.B(n_91),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx24_ASAP7_75t_SL g167 ( 
.A(n_16),
.Y(n_167)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_50),
.CI(n_76),
.CON(n_16),
.SN(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_34),
.B2(n_35),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_27),
.B(n_29),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_27),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_26),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_27),
.B(n_33),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_28),
.A2(n_30),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_28),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_31),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_32),
.B(n_145),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_33),
.A2(n_39),
.B(n_45),
.C(n_116),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_33),
.B(n_44),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_33),
.A2(n_38),
.B(n_55),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_34),
.A2(n_35),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_34),
.A2(n_35),
.B1(n_51),
.B2(n_95),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_35),
.B(n_115),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_35),
.B(n_51),
.C(n_147),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_46),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_37),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_39),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_47),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_63),
.C(n_73),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_73),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_59),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_56),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_54),
.B(n_58),
.C(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_58),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_57),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_63),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_69),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_85),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_78),
.A2(n_79),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_102),
.C(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_123),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_89),
.A2(n_99),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_89),
.B(n_131),
.C(n_134),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_90),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_98),
.C(n_100),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_92),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_98),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_102),
.A2(n_103),
.B1(n_119),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_102),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_103),
.B(n_113),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_160),
.B(n_165),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_149),
.B(n_159),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_136),
.B(n_148),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_126),
.B(n_135),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_117),
.B(n_125),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_122),
.B(n_124),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_128),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_134),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_152),
.C(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_138),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_147),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_141),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_150),
.B(n_151),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);


endmodule