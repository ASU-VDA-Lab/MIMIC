module fake_netlist_1_2343_n_1097 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1097);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1097;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_801;
wire n_988;
wire n_1059;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_1022;
wire n_918;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_1042;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_529;
wire n_455;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_624;
wire n_426;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_459;
wire n_863;
wire n_322;
wire n_907;
wire n_708;
wire n_1062;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_1046;
wire n_460;
wire n_935;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_937;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_653;
wire n_357;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1088;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_1043;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_504;
wire n_581;
wire n_458;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_772;
wire n_405;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
INVx1_ASAP7_75t_L g316 ( .A(n_73), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_274), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_171), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_312), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_34), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_10), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_202), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_277), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_213), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_162), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_196), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_297), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_158), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_106), .Y(n_331) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_19), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_88), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_3), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_136), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_192), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_267), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_151), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_206), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_120), .Y(n_340) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_63), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_39), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_58), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_127), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_39), .Y(n_345) );
INVx4_ASAP7_75t_R g346 ( .A(n_308), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_293), .Y(n_347) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_52), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_257), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_4), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_222), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_285), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_218), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_301), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_184), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_278), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_219), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_187), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_70), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_269), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_265), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_180), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_76), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_156), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_10), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_71), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_131), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_64), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_155), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_84), .Y(n_372) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_310), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_106), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_35), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_96), .Y(n_376) );
CKINVDCx5p33_ASAP7_75t_R g377 ( .A(n_240), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_189), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_6), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_176), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_115), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_40), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_233), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_253), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_245), .Y(n_385) );
CKINVDCx16_ASAP7_75t_R g386 ( .A(n_255), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_242), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_289), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_35), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_307), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_95), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_304), .Y(n_392) );
BUFx5_ASAP7_75t_L g393 ( .A(n_247), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_313), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_309), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_168), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_103), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_256), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_135), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_250), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_47), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_67), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_169), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_263), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_100), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_153), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_74), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_121), .Y(n_408) );
INVxp33_ASAP7_75t_SL g409 ( .A(n_264), .Y(n_409) );
INVxp33_ASAP7_75t_SL g410 ( .A(n_251), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_64), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_214), .B(n_268), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_273), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_272), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_127), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_221), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_97), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_161), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_244), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_53), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_260), .Y(n_421) );
CKINVDCx14_ASAP7_75t_R g422 ( .A(n_63), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_243), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_150), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_305), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_111), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_296), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_0), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_284), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_75), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_182), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_303), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_258), .Y(n_433) );
CKINVDCx14_ASAP7_75t_R g434 ( .A(n_89), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_153), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_13), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_40), .Y(n_437) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_80), .Y(n_438) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_197), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_37), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_259), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_82), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_311), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_77), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_86), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_25), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_79), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_61), .Y(n_448) );
NOR2xp67_ASAP7_75t_L g449 ( .A(n_85), .B(n_190), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_238), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_11), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_116), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_280), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_72), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_266), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_74), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_330), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_400), .B(n_0), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_400), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_330), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_422), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_331), .Y(n_463) );
XOR2xp5_ASAP7_75t_L g464 ( .A(n_333), .B(n_1), .Y(n_464) );
NAND2xp33_ASAP7_75t_L g465 ( .A(n_393), .B(n_179), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_322), .B(n_1), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_331), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_341), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_350), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_390), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_393), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_422), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_390), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_350), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_379), .B(n_2), .Y(n_475) );
INVx2_ASAP7_75t_SL g476 ( .A(n_351), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_341), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_379), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_382), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_393), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_383), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_318), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_382), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_393), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_415), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_417), .B(n_3), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_393), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_460), .B(n_354), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_459), .B(n_458), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_459), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_460), .B(n_354), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_462), .B(n_434), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_462), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_471), .Y(n_494) );
INVx2_ASAP7_75t_SL g495 ( .A(n_459), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_458), .B(n_378), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_460), .B(n_378), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_481), .B(n_386), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_471), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_471), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_481), .B(n_385), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_458), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_472), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g504 ( .A(n_476), .B(n_336), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_458), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_480), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_476), .B(n_347), .Y(n_507) );
AND2x4_ASAP7_75t_L g508 ( .A(n_475), .B(n_415), .Y(n_508) );
INVx5_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
AND2x6_ASAP7_75t_SL g510 ( .A(n_486), .B(n_316), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_466), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_458), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_458), .B(n_385), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_480), .Y(n_514) );
NOR2xp33_ASAP7_75t_SL g515 ( .A(n_475), .B(n_432), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_475), .Y(n_516) );
INVx4_ASAP7_75t_L g517 ( .A(n_475), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_503), .B(n_486), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_492), .B(n_466), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_492), .B(n_476), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_493), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_490), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_492), .B(n_441), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_516), .A2(n_410), .B1(n_409), .B2(n_480), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_516), .B(n_457), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_498), .B(n_332), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_490), .B(n_484), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_508), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_490), .B(n_484), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_490), .B(n_484), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_501), .B(n_443), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_508), .Y(n_532) );
AO22x1_ASAP7_75t_L g533 ( .A1(n_498), .A2(n_410), .B1(n_409), .B2(n_335), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_516), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_502), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_516), .A2(n_487), .B1(n_319), .B2(n_334), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_501), .B(n_329), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_502), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_505), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_516), .A2(n_487), .B1(n_327), .B2(n_340), .Y(n_540) );
OAI21xp33_ASAP7_75t_L g541 ( .A1(n_515), .A2(n_342), .B(n_338), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_504), .B(n_329), .Y(n_542) );
AND2x6_ASAP7_75t_L g543 ( .A(n_508), .B(n_317), .Y(n_543) );
AOI21x1_ASAP7_75t_L g544 ( .A1(n_489), .A2(n_487), .B(n_323), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_508), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_495), .B(n_320), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_505), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_508), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_489), .A2(n_465), .B(n_421), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_505), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_517), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_358), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_517), .A2(n_344), .B1(n_365), .B2(n_345), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_507), .B(n_457), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_517), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_517), .A2(n_366), .B1(n_368), .B2(n_367), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_488), .Y(n_557) );
NAND2x1_ASAP7_75t_L g558 ( .A(n_495), .B(n_346), .Y(n_558) );
AND2x6_ASAP7_75t_L g559 ( .A(n_488), .B(n_324), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_491), .Y(n_560) );
AND2x4_ASAP7_75t_L g561 ( .A(n_511), .B(n_461), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_493), .B(n_515), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_491), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_497), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_512), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_497), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_494), .A2(n_343), .B1(n_361), .B2(n_321), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_510), .B(n_461), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_494), .B(n_384), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_509), .Y(n_570) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_510), .B(n_463), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_499), .B(n_388), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_513), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_500), .B(n_463), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_568), .A2(n_506), .B1(n_514), .B2(n_500), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_526), .B(n_464), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_521), .Y(n_578) );
OR2x6_ASAP7_75t_L g579 ( .A(n_533), .B(n_438), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_571), .B(n_388), .Y(n_580) );
INVx5_ASAP7_75t_L g581 ( .A(n_543), .Y(n_581) );
O2A1O1Ixp5_ASAP7_75t_L g582 ( .A1(n_554), .A2(n_496), .B(n_514), .C(n_512), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_522), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_557), .B(n_361), .Y(n_584) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_562), .B(n_369), .Y(n_585) );
INVx4_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_561), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_545), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_562), .A2(n_372), .B1(n_389), .B2(n_371), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_518), .B(n_523), .Y(n_590) );
BUFx6f_ASAP7_75t_L g591 ( .A(n_571), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_554), .A2(n_380), .B(n_376), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_560), .A2(n_391), .B1(n_405), .B2(n_374), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
AO31x2_ASAP7_75t_L g595 ( .A1(n_549), .A2(n_421), .A3(n_414), .B(n_326), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_572), .A2(n_430), .B1(n_440), .B2(n_405), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_534), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_563), .B(n_396), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_561), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_564), .B(n_399), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_566), .Y(n_601) );
INVx3_ASAP7_75t_L g602 ( .A(n_525), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_525), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_519), .B(n_399), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_541), .A2(n_408), .B1(n_420), .B2(n_411), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_531), .B(n_408), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_570), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_551), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_537), .B(n_394), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_528), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_532), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_548), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_574), .B(n_411), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_529), .A2(n_509), .B(n_439), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_530), .A2(n_328), .B(n_325), .Y(n_617) );
INVx4_ASAP7_75t_L g618 ( .A(n_543), .Y(n_618) );
AOI21x1_ASAP7_75t_L g619 ( .A1(n_544), .A2(n_339), .B(n_337), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_575), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_520), .B(n_435), .Y(n_621) );
NAND2x1_ASAP7_75t_SL g622 ( .A(n_567), .B(n_449), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_559), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_572), .B(n_348), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_553), .B(n_370), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_542), .B(n_444), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_530), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_552), .B(n_444), .Y(n_628) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_570), .Y(n_629) );
BUFx2_ASAP7_75t_L g630 ( .A(n_559), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_524), .A2(n_454), .B1(n_445), .B2(n_375), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_546), .A2(n_373), .B(n_509), .Y(n_632) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_546), .A2(n_381), .B(n_424), .C(n_401), .Y(n_633) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_536), .A2(n_402), .B(n_403), .C(n_397), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_569), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_570), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_556), .B(n_406), .Y(n_637) );
O2A1O1Ixp5_ASAP7_75t_SL g638 ( .A1(n_573), .A2(n_469), .B(n_474), .C(n_467), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_559), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
AND2x4_ASAP7_75t_L g641 ( .A(n_540), .B(n_407), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_558), .B(n_448), .C(n_445), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_535), .A2(n_428), .B1(n_436), .B2(n_426), .Y(n_643) );
INVx3_ASAP7_75t_L g644 ( .A(n_535), .Y(n_644) );
BUFx2_ASAP7_75t_SL g645 ( .A(n_538), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_538), .B(n_437), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_539), .A2(n_446), .B(n_447), .C(n_442), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_565), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_547), .B(n_451), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_550), .Y(n_650) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_565), .A2(n_456), .B(n_452), .C(n_467), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_557), .B(n_509), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_527), .A2(n_509), .B(n_349), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_557), .B(n_509), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_601), .B(n_418), .Y(n_655) );
OAI21x1_ASAP7_75t_L g656 ( .A1(n_619), .A2(n_414), .B(n_412), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_578), .Y(n_657) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_638), .A2(n_353), .B(n_352), .Y(n_658) );
OAI21x1_ASAP7_75t_L g659 ( .A1(n_653), .A2(n_356), .B(n_355), .Y(n_659) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_582), .A2(n_359), .B(n_357), .Y(n_660) );
OAI21x1_ASAP7_75t_L g661 ( .A1(n_653), .A2(n_362), .B(n_360), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_606), .A2(n_364), .B(n_363), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_607), .B(n_478), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_581), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_579), .A2(n_479), .B1(n_483), .B2(n_478), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_579), .A2(n_483), .B1(n_485), .B2(n_479), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_586), .Y(n_667) );
OAI21x1_ASAP7_75t_SL g668 ( .A1(n_618), .A2(n_392), .B(n_387), .Y(n_668) );
OAI21x1_ASAP7_75t_L g669 ( .A1(n_644), .A2(n_398), .B(n_395), .Y(n_669) );
AO31x2_ASAP7_75t_L g670 ( .A1(n_651), .A2(n_647), .A3(n_646), .B(n_643), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_635), .A2(n_590), .B(n_620), .C(n_633), .Y(n_671) );
AO32x2_ASAP7_75t_L g672 ( .A1(n_643), .A2(n_470), .A3(n_473), .B1(n_482), .B2(n_341), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_649), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_645), .A2(n_482), .B1(n_416), .B2(n_419), .Y(n_674) );
OAI21x1_ASAP7_75t_L g675 ( .A1(n_632), .A2(n_423), .B(n_413), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_609), .Y(n_676) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_648), .A2(n_427), .B(n_425), .Y(n_677) );
BUFx6f_ASAP7_75t_L g678 ( .A(n_608), .Y(n_678) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_608), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_585), .A2(n_393), .B1(n_433), .B2(n_404), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_592), .A2(n_482), .B1(n_429), .B2(n_431), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_652), .A2(n_654), .B(n_598), .Y(n_682) );
INVx3_ASAP7_75t_L g683 ( .A(n_586), .Y(n_683) );
AO22x2_ASAP7_75t_L g684 ( .A1(n_593), .A2(n_453), .B1(n_450), .B2(n_455), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_577), .B(n_377), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_652), .A2(n_654), .B(n_598), .Y(n_686) );
OA21x2_ASAP7_75t_L g687 ( .A1(n_617), .A2(n_393), .B(n_470), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_581), .B(n_4), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_611), .Y(n_689) );
BUFx4f_ASAP7_75t_L g690 ( .A(n_591), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_650), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_584), .A2(n_477), .B(n_468), .Y(n_692) );
OAI21x1_ASAP7_75t_L g693 ( .A1(n_616), .A2(n_473), .B(n_470), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_602), .Y(n_694) );
AOI22x1_ASAP7_75t_L g695 ( .A1(n_639), .A2(n_473), .B1(n_470), .B2(n_181), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_587), .Y(n_696) );
AO22x2_ASAP7_75t_L g697 ( .A1(n_623), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_606), .A2(n_473), .B(n_470), .C(n_8), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_583), .A2(n_473), .B(n_470), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_591), .Y(n_700) );
AO31x2_ASAP7_75t_L g701 ( .A1(n_634), .A2(n_8), .A3(n_5), .B(n_7), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_600), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_602), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_603), .Y(n_704) );
OAI21x1_ASAP7_75t_SL g705 ( .A1(n_600), .A2(n_9), .B(n_11), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_627), .A2(n_185), .B(n_183), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_615), .A2(n_9), .B(n_12), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g708 ( .A1(n_576), .A2(n_12), .B(n_14), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_612), .B(n_14), .Y(n_709) );
AO22x2_ASAP7_75t_L g710 ( .A1(n_599), .A2(n_17), .B1(n_15), .B2(n_16), .Y(n_710) );
OAI21x1_ASAP7_75t_L g711 ( .A1(n_594), .A2(n_188), .B(n_186), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_613), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_624), .B(n_18), .Y(n_713) );
OAI21x1_ASAP7_75t_L g714 ( .A1(n_594), .A2(n_597), .B(n_614), .Y(n_714) );
OA21x2_ASAP7_75t_L g715 ( .A1(n_622), .A2(n_193), .B(n_191), .Y(n_715) );
O2A1O1Ixp33_ASAP7_75t_L g716 ( .A1(n_604), .A2(n_21), .B(n_18), .C(n_20), .Y(n_716) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_597), .A2(n_195), .B(n_194), .Y(n_717) );
OAI21x1_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_199), .B(n_198), .Y(n_718) );
AND2x2_ASAP7_75t_L g719 ( .A(n_626), .B(n_20), .Y(n_719) );
O2A1O1Ixp33_ASAP7_75t_L g720 ( .A1(n_604), .A2(n_23), .B(n_21), .C(n_22), .Y(n_720) );
OAI21x1_ASAP7_75t_L g721 ( .A1(n_640), .A2(n_201), .B(n_200), .Y(n_721) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_630), .B(n_203), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_608), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_588), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_641), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_624), .A2(n_26), .B1(n_24), .B2(n_25), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_637), .B(n_24), .Y(n_727) );
INVx1_ASAP7_75t_SL g728 ( .A(n_629), .Y(n_728) );
BUFx2_ASAP7_75t_L g729 ( .A(n_625), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_637), .A2(n_26), .B(n_27), .Y(n_730) );
OA21x2_ASAP7_75t_L g731 ( .A1(n_595), .A2(n_205), .B(n_204), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_625), .B(n_28), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_621), .B(n_29), .Y(n_733) );
OR2x6_ASAP7_75t_L g734 ( .A(n_629), .B(n_30), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_589), .B(n_628), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g736 ( .A1(n_605), .A2(n_33), .B1(n_31), .B2(n_32), .Y(n_736) );
AOI21x1_ASAP7_75t_L g737 ( .A1(n_610), .A2(n_580), .B(n_595), .Y(n_737) );
OAI21x1_ASAP7_75t_L g738 ( .A1(n_595), .A2(n_208), .B(n_207), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_642), .B(n_32), .Y(n_739) );
OAI21x1_ASAP7_75t_L g740 ( .A1(n_636), .A2(n_210), .B(n_209), .Y(n_740) );
NOR2xp33_ASAP7_75t_SL g741 ( .A(n_636), .B(n_211), .Y(n_741) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_596), .A2(n_36), .B1(n_33), .B2(n_34), .Y(n_742) );
OAI21xp33_ASAP7_75t_SL g743 ( .A1(n_631), .A2(n_38), .B(n_41), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_665), .A2(n_44), .B1(n_42), .B2(n_43), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g745 ( .A1(n_666), .A2(n_46), .B1(n_44), .B2(n_45), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_666), .A2(n_729), .B1(n_680), .B2(n_702), .Y(n_746) );
OA21x2_ASAP7_75t_L g747 ( .A1(n_738), .A2(n_215), .B(n_212), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_710), .Y(n_748) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_735), .B(n_48), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_684), .A2(n_51), .B1(n_49), .B2(n_50), .Y(n_750) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_678), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_710), .Y(n_752) );
OR2x6_ASAP7_75t_L g753 ( .A(n_734), .B(n_51), .Y(n_753) );
OA21x2_ASAP7_75t_L g754 ( .A1(n_656), .A2(n_217), .B(n_216), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_657), .Y(n_755) );
AO31x2_ASAP7_75t_L g756 ( .A1(n_698), .A2(n_56), .A3(n_54), .B(n_55), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g757 ( .A1(n_743), .A2(n_57), .B(n_55), .C(n_56), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_684), .A2(n_61), .B1(n_59), .B2(n_60), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_671), .B(n_62), .Y(n_759) );
INVx1_ASAP7_75t_SL g760 ( .A(n_691), .Y(n_760) );
AOI222xp33_ASAP7_75t_L g761 ( .A1(n_742), .A2(n_65), .B1(n_66), .B2(n_67), .C1(n_68), .C2(n_69), .Y(n_761) );
AO31x2_ASAP7_75t_L g762 ( .A1(n_681), .A2(n_81), .A3(n_78), .B(n_79), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_719), .B(n_83), .Y(n_763) );
BUFx8_ASAP7_75t_L g764 ( .A(n_688), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_709), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_709), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_655), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_676), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_713), .A2(n_91), .B1(n_87), .B2(n_90), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_725), .B(n_92), .Y(n_770) );
OAI21x1_ASAP7_75t_L g771 ( .A1(n_699), .A2(n_223), .B(n_220), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_673), .A2(n_96), .B1(n_93), .B2(n_94), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_685), .B(n_97), .Y(n_773) );
OR2x6_ASAP7_75t_L g774 ( .A(n_734), .B(n_98), .Y(n_774) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_688), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_727), .A2(n_100), .B1(n_98), .B2(n_99), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_655), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_712), .Y(n_778) );
AND2x2_ASAP7_75t_L g779 ( .A(n_696), .B(n_99), .Y(n_779) );
AOI222xp33_ASAP7_75t_L g780 ( .A1(n_730), .A2(n_101), .B1(n_102), .B2(n_103), .C1(n_104), .C2(n_105), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_689), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_732), .Y(n_782) );
INVx5_ASAP7_75t_SL g783 ( .A(n_663), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_662), .B(n_107), .Y(n_784) );
AOI222xp33_ASAP7_75t_L g785 ( .A1(n_708), .A2(n_108), .B1(n_109), .B2(n_110), .C1(n_111), .C2(n_112), .Y(n_785) );
OAI221xp5_ASAP7_75t_SL g786 ( .A1(n_726), .A2(n_109), .B1(n_110), .B2(n_112), .C(n_113), .Y(n_786) );
OAI21xp5_ASAP7_75t_L g787 ( .A1(n_682), .A2(n_113), .B(n_114), .Y(n_787) );
OAI21xp5_ASAP7_75t_L g788 ( .A1(n_682), .A2(n_117), .B(n_118), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_686), .A2(n_122), .B1(n_119), .B2(n_121), .Y(n_789) );
AO21x2_ASAP7_75t_L g790 ( .A1(n_660), .A2(n_225), .B(n_224), .Y(n_790) );
OAI221xp5_ASAP7_75t_SL g791 ( .A1(n_736), .A2(n_122), .B1(n_123), .B2(n_124), .C(n_125), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_704), .Y(n_792) );
A2O1A1Ixp33_ASAP7_75t_L g793 ( .A1(n_707), .A2(n_129), .B(n_126), .C(n_128), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_701), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_690), .Y(n_795) );
BUFx8_ASAP7_75t_L g796 ( .A(n_700), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_733), .A2(n_133), .B1(n_130), .B2(n_132), .Y(n_797) );
OAI211xp5_ASAP7_75t_L g798 ( .A1(n_739), .A2(n_707), .B(n_720), .C(n_716), .Y(n_798) );
BUFx2_ASAP7_75t_L g799 ( .A(n_667), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g800 ( .A1(n_674), .A2(n_136), .B1(n_134), .B2(n_135), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_670), .B(n_137), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_674), .A2(n_138), .B1(n_139), .B2(n_140), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_701), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_724), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_663), .A2(n_141), .B1(n_142), .B2(n_143), .Y(n_805) );
OAI22xp5_ASAP7_75t_L g806 ( .A1(n_697), .A2(n_144), .B1(n_145), .B2(n_146), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_683), .Y(n_807) );
OAI21x1_ASAP7_75t_L g808 ( .A1(n_693), .A2(n_227), .B(n_226), .Y(n_808) );
OAI211xp5_ASAP7_75t_L g809 ( .A1(n_716), .A2(n_147), .B(n_148), .C(n_149), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_705), .Y(n_810) );
AND2x4_ASAP7_75t_L g811 ( .A(n_664), .B(n_152), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_670), .B(n_154), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_692), .A2(n_668), .B1(n_703), .B2(n_694), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_697), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_722), .A2(n_155), .B1(n_157), .B2(n_158), .Y(n_815) );
AO21x2_ASAP7_75t_L g816 ( .A1(n_658), .A2(n_229), .B(n_228), .Y(n_816) );
A2O1A1Ixp33_ASAP7_75t_L g817 ( .A1(n_720), .A2(n_159), .B(n_160), .C(n_161), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_670), .B(n_163), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_669), .B(n_164), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_675), .B(n_165), .Y(n_820) );
HB1xp67_ASAP7_75t_L g821 ( .A(n_760), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_794), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_768), .B(n_672), .Y(n_823) );
INVx2_ASAP7_75t_SL g824 ( .A(n_796), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_755), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_778), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_781), .Y(n_827) );
AND2x4_ASAP7_75t_L g828 ( .A(n_753), .B(n_723), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_808), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_749), .B(n_737), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_804), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_767), .B(n_672), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_751), .Y(n_833) );
INVx5_ASAP7_75t_L g834 ( .A(n_753), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_777), .B(n_715), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_803), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_782), .B(n_677), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_771), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_765), .Y(n_839) );
NAND3xp33_ASAP7_75t_L g840 ( .A(n_785), .B(n_731), .C(n_695), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_766), .B(n_687), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_792), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_780), .B(n_728), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_774), .B(n_714), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_747), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_774), .B(n_731), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_754), .Y(n_847) );
INVx2_ASAP7_75t_L g848 ( .A(n_754), .Y(n_848) );
BUFx2_ASAP7_75t_L g849 ( .A(n_775), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_801), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_812), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_818), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_748), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_811), .Y(n_854) );
OR2x2_ASAP7_75t_L g855 ( .A(n_752), .B(n_679), .Y(n_855) );
AND2x4_ASAP7_75t_L g856 ( .A(n_810), .B(n_679), .Y(n_856) );
INVx2_ASAP7_75t_SL g857 ( .A(n_764), .Y(n_857) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_820), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_816), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_756), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_787), .B(n_711), .Y(n_861) );
OR2x2_ASAP7_75t_L g862 ( .A(n_814), .B(n_659), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_756), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_783), .B(n_661), .Y(n_864) );
INVx2_ASAP7_75t_SL g865 ( .A(n_795), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_787), .B(n_717), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_779), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_756), .Y(n_868) );
AND2x4_ASAP7_75t_L g869 ( .A(n_799), .B(n_718), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_783), .B(n_166), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_762), .Y(n_871) );
BUFx2_ASAP7_75t_L g872 ( .A(n_807), .Y(n_872) );
INVx2_ASAP7_75t_L g873 ( .A(n_762), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_788), .B(n_721), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_750), .B(n_706), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_791), .A2(n_741), .B1(n_168), .B2(n_169), .C(n_170), .Y(n_876) );
OR2x6_ASAP7_75t_L g877 ( .A(n_806), .B(n_740), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_758), .B(n_167), .Y(n_878) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_763), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_761), .B(n_170), .Y(n_880) );
AND2x4_ASAP7_75t_L g881 ( .A(n_813), .B(n_790), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_759), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_746), .B(n_171), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_819), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_806), .Y(n_885) );
AO21x2_ASAP7_75t_L g886 ( .A1(n_798), .A2(n_172), .B(n_173), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_770), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_784), .Y(n_888) );
INVxp33_ASAP7_75t_L g889 ( .A(n_773), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_793), .B(n_174), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_815), .B(n_230), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_776), .B(n_175), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_744), .B(n_176), .Y(n_893) );
OR2x2_ASAP7_75t_L g894 ( .A(n_797), .B(n_177), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_817), .B(n_178), .Y(n_895) );
INVx4_ASAP7_75t_L g896 ( .A(n_745), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_800), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_802), .Y(n_898) );
OR2x2_ASAP7_75t_L g899 ( .A(n_786), .B(n_231), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_789), .B(n_232), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_809), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_889), .B(n_757), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_879), .B(n_805), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_821), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_825), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_826), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_827), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_839), .B(n_769), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_867), .B(n_772), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_831), .Y(n_910) );
AND2x2_ASAP7_75t_L g911 ( .A(n_880), .B(n_234), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_822), .Y(n_912) );
OAI33xp33_ASAP7_75t_L g913 ( .A1(n_883), .A2(n_235), .A3(n_236), .B1(n_237), .B2(n_239), .B3(n_241), .Y(n_913) );
INVx2_ASAP7_75t_SL g914 ( .A(n_834), .Y(n_914) );
INVx3_ASAP7_75t_L g915 ( .A(n_869), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_839), .B(n_842), .Y(n_916) );
INVxp67_ASAP7_75t_L g917 ( .A(n_872), .Y(n_917) );
OAI33xp33_ASAP7_75t_L g918 ( .A1(n_894), .A2(n_246), .A3(n_248), .B1(n_249), .B2(n_252), .B3(n_254), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_822), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_836), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_849), .B(n_314), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_841), .Y(n_922) );
INVx2_ASAP7_75t_L g923 ( .A(n_841), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_871), .Y(n_924) );
NOR2x1_ASAP7_75t_SL g925 ( .A(n_834), .B(n_261), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_853), .Y(n_926) );
AND2x4_ASAP7_75t_L g927 ( .A(n_844), .B(n_262), .Y(n_927) );
INVx4_ASAP7_75t_L g928 ( .A(n_834), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_853), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_873), .Y(n_930) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_896), .B(n_270), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_873), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_854), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_824), .B(n_271), .Y(n_934) );
AO21x2_ASAP7_75t_L g935 ( .A1(n_840), .A2(n_275), .B(n_276), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_888), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_870), .B(n_279), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_888), .Y(n_938) );
INVx4_ASAP7_75t_L g939 ( .A(n_834), .Y(n_939) );
AND2x4_ASAP7_75t_L g940 ( .A(n_844), .B(n_281), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_843), .A2(n_282), .B1(n_283), .B2(n_286), .Y(n_941) );
OR2x6_ASAP7_75t_L g942 ( .A(n_891), .B(n_287), .Y(n_942) );
OAI33xp33_ASAP7_75t_L g943 ( .A1(n_892), .A2(n_290), .A3(n_291), .B1(n_292), .B2(n_294), .B3(n_295), .Y(n_943) );
HB1xp67_ASAP7_75t_L g944 ( .A(n_855), .Y(n_944) );
INVx3_ASAP7_75t_L g945 ( .A(n_869), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_823), .Y(n_946) );
NOR4xp75_ASAP7_75t_L g947 ( .A(n_857), .B(n_298), .C(n_300), .D(n_302), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_855), .Y(n_948) );
INVx2_ASAP7_75t_L g949 ( .A(n_832), .Y(n_949) );
OA21x2_ASAP7_75t_L g950 ( .A1(n_847), .A2(n_848), .B(n_845), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_885), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_832), .Y(n_952) );
INVx2_ASAP7_75t_L g953 ( .A(n_860), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_885), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_862), .Y(n_955) );
AND2x6_ASAP7_75t_L g956 ( .A(n_846), .B(n_869), .Y(n_956) );
AND2x2_ASAP7_75t_L g957 ( .A(n_893), .B(n_878), .Y(n_957) );
BUFx2_ASAP7_75t_L g958 ( .A(n_828), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_887), .B(n_884), .Y(n_959) );
INVx3_ASAP7_75t_L g960 ( .A(n_856), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_860), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_837), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_863), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g964 ( .A(n_897), .B(n_898), .Y(n_964) );
NAND3xp33_ASAP7_75t_L g965 ( .A(n_902), .B(n_901), .C(n_876), .Y(n_965) );
INVx3_ASAP7_75t_L g966 ( .A(n_928), .Y(n_966) );
OR2x2_ASAP7_75t_L g967 ( .A(n_922), .B(n_850), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_922), .B(n_868), .Y(n_968) );
AND2x2_ASAP7_75t_L g969 ( .A(n_923), .B(n_868), .Y(n_969) );
AND2x2_ASAP7_75t_SL g970 ( .A(n_927), .B(n_891), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_905), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_906), .Y(n_972) );
INVx1_ASAP7_75t_L g973 ( .A(n_907), .Y(n_973) );
OR2x2_ASAP7_75t_L g974 ( .A(n_904), .B(n_851), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_910), .Y(n_975) );
INVx2_ASAP7_75t_SL g976 ( .A(n_928), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_916), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_923), .B(n_852), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_919), .Y(n_979) );
AND2x4_ASAP7_75t_L g980 ( .A(n_915), .B(n_881), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_912), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_920), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_944), .B(n_830), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_924), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_959), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_948), .B(n_864), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_933), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g988 ( .A1(n_942), .A2(n_899), .B1(n_890), .B2(n_895), .Y(n_988) );
OR2x2_ASAP7_75t_L g989 ( .A(n_917), .B(n_882), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_926), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_929), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_936), .Y(n_992) );
INVx2_ASAP7_75t_SL g993 ( .A(n_939), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_938), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_917), .B(n_858), .Y(n_995) );
OR2x2_ASAP7_75t_L g996 ( .A(n_964), .B(n_858), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_957), .B(n_833), .Y(n_997) );
INVx2_ASAP7_75t_SL g998 ( .A(n_939), .Y(n_998) );
AND2x4_ASAP7_75t_L g999 ( .A(n_945), .B(n_858), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_930), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_955), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_951), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_902), .A2(n_886), .B1(n_900), .B2(n_861), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_949), .B(n_835), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_954), .B(n_835), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_955), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_949), .B(n_858), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_952), .B(n_866), .Y(n_1008) );
INVx2_ASAP7_75t_L g1009 ( .A(n_932), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_903), .B(n_866), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_952), .B(n_877), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_909), .B(n_875), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_958), .B(n_865), .Y(n_1013) );
INVx2_ASAP7_75t_L g1014 ( .A(n_950), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_946), .B(n_877), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_950), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g1017 ( .A(n_942), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_980), .B(n_945), .Y(n_1018) );
INVx1_ASAP7_75t_L g1019 ( .A(n_971), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_972), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_977), .B(n_962), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_1010), .B(n_960), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_1008), .B(n_956), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_1011), .B(n_956), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_973), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_965), .B(n_931), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_975), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_985), .B(n_960), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_987), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1014), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1031 ( .A(n_983), .B(n_953), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_979), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_982), .Y(n_1033) );
NOR2x1_ASAP7_75t_R g1034 ( .A(n_1017), .B(n_911), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_967), .B(n_961), .Y(n_1035) );
INVx3_ASAP7_75t_L g1036 ( .A(n_966), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_970), .A2(n_941), .B1(n_921), .B2(n_937), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_997), .B(n_940), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_1012), .B(n_908), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1011), .B(n_961), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_978), .B(n_940), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_990), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_1015), .B(n_963), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_991), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_974), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1002), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1004), .B(n_859), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_986), .B(n_914), .Y(n_1048) );
INVx2_ASAP7_75t_L g1049 ( .A(n_1016), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1019), .Y(n_1050) );
AOI21xp33_ASAP7_75t_L g1051 ( .A1(n_1026), .A2(n_988), .B(n_1013), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1020), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1025), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_1039), .B(n_1006), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1027), .Y(n_1055) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_1037), .A2(n_1003), .B1(n_998), .B2(n_993), .Y(n_1056) );
NOR2xp33_ASAP7_75t_L g1057 ( .A(n_1034), .B(n_934), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_1045), .B(n_1001), .Y(n_1058) );
NAND2xp5_ASAP7_75t_SL g1059 ( .A(n_1036), .B(n_976), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1029), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1032), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_1033), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_1051), .A2(n_1044), .B1(n_1042), .B2(n_1046), .C(n_1021), .Y(n_1063) );
AND2x4_ASAP7_75t_L g1064 ( .A(n_1059), .B(n_1018), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1058), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_1050), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1052), .Y(n_1067) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_1053), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1055), .Y(n_1069) );
OAI322xp33_ASAP7_75t_L g1070 ( .A1(n_1056), .A2(n_1022), .A3(n_1028), .B1(n_1048), .B2(n_1031), .C1(n_1035), .C2(n_1041), .Y(n_1070) );
AOI22xp33_ASAP7_75t_SL g1071 ( .A1(n_1057), .A2(n_1023), .B1(n_1038), .B2(n_1024), .Y(n_1071) );
AOI221xp5_ASAP7_75t_L g1072 ( .A1(n_1070), .A2(n_1054), .B1(n_1062), .B2(n_1060), .C(n_1061), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1068), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_1071), .A2(n_1043), .B1(n_1040), .B2(n_989), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g1075 ( .A1(n_1063), .A2(n_1043), .B1(n_913), .B2(n_992), .C(n_994), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_1065), .B(n_1047), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_1072), .A2(n_1069), .B1(n_1067), .B2(n_1066), .C(n_1064), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1076), .Y(n_1078) );
NOR3xp33_ASAP7_75t_L g1079 ( .A(n_1075), .B(n_918), .C(n_943), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_1074), .A2(n_996), .B1(n_1005), .B2(n_995), .C(n_1030), .Y(n_1080) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_1073), .Y(n_1081) );
NAND2xp5_ASAP7_75t_L g1082 ( .A(n_1078), .B(n_1049), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1081), .Y(n_1083) );
NAND5xp2_ASAP7_75t_L g1084 ( .A(n_1077), .B(n_874), .C(n_947), .D(n_925), .E(n_1007), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1080), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1085), .B(n_1079), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1083), .Y(n_1087) );
NAND4xp25_ASAP7_75t_L g1088 ( .A(n_1084), .B(n_999), .C(n_1007), .D(n_968), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1087), .Y(n_1089) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_1088), .A2(n_1082), .B1(n_999), .B2(n_935), .Y(n_1090) );
OAI22xp33_ASAP7_75t_SL g1091 ( .A1(n_1086), .A2(n_981), .B1(n_1009), .B2(n_1000), .Y(n_1091) );
OAI21xp5_ASAP7_75t_L g1092 ( .A1(n_1089), .A2(n_829), .B(n_838), .Y(n_1092) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1091), .Y(n_1093) );
XOR2xp5_ASAP7_75t_L g1094 ( .A(n_1093), .B(n_1090), .Y(n_1094) );
OAI21xp5_ASAP7_75t_L g1095 ( .A1(n_1094), .A2(n_1092), .B(n_829), .Y(n_1095) );
BUFx3_ASAP7_75t_L g1096 ( .A(n_1095), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_1096), .A2(n_1004), .B1(n_969), .B2(n_984), .Y(n_1097) );
endmodule