module real_jpeg_32329_n_21 (n_17, n_8, n_0, n_157, n_2, n_10, n_9, n_12, n_154, n_156, n_152, n_6, n_159, n_153, n_151, n_161, n_11, n_14, n_160, n_7, n_18, n_3, n_5, n_4, n_1, n_20, n_19, n_158, n_16, n_15, n_13, n_155, n_21);

input n_17;
input n_8;
input n_0;
input n_157;
input n_2;
input n_10;
input n_9;
input n_12;
input n_154;
input n_156;
input n_152;
input n_6;
input n_159;
input n_153;
input n_151;
input n_161;
input n_11;
input n_14;
input n_160;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_20;
input n_19;
input n_158;
input n_16;
input n_15;
input n_13;
input n_155;

output n_21;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_0),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_0),
.B(n_75),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_1),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_1),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_2),
.A2(n_145),
.B1(n_146),
.B2(n_149),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_2),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_25),
.Y(n_24)
);

AOI221xp5_ASAP7_75t_L g91 ( 
.A1(n_5),
.A2(n_10),
.B1(n_92),
.B2(n_96),
.C(n_98),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_5),
.B(n_92),
.C(n_96),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_6),
.B(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_9),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_10),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_12),
.B(n_24),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_13),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_13),
.A2(n_61),
.A3(n_63),
.B1(n_68),
.B2(n_129),
.C1(n_131),
.C2(n_161),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_14),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_14),
.B(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_15),
.B(n_70),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_17),
.B(n_44),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_18),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_20),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_144),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B(n_143),
.Y(n_22)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_136),
.B(n_140),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_41),
.B(n_135),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_40),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_33),
.B(n_40),
.Y(n_135)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B(n_134),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI31xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_80),
.A3(n_117),
.B(n_124),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_67),
.C(n_74),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_53),
.A2(n_125),
.B(n_128),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR3xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_74),
.C(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_152),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

OA21x2_ASAP7_75t_SL g125 ( 
.A1(n_67),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_111),
.C(n_112),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_102),
.B(n_110),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_91),
.B1(n_100),
.B2(n_101),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_157),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_109),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_151),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_153),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_154),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_155),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_156),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_158),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_159),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_160),
.Y(n_120)
);


endmodule