module fake_jpeg_18735_n_225 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_26),
.Y(n_47)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_53),
.B(n_39),
.Y(n_60)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_1),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_35),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_64),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_21),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_43),
.B(n_49),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_41),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_28),
.B1(n_27),
.B2(n_32),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_73),
.A2(n_34),
.B1(n_25),
.B2(n_32),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_28),
.B1(n_36),
.B2(n_24),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_77),
.B1(n_25),
.B2(n_29),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_36),
.B1(n_23),
.B2(n_24),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_48),
.C(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_85),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_35),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_87),
.B(n_93),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_54),
.B1(n_58),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_88),
.A2(n_92),
.B1(n_96),
.B2(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_91),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_58),
.B1(n_47),
.B2(n_52),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_99),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_101),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_98),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_18),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_110),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_35),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_64),
.A2(n_82),
.B1(n_70),
.B2(n_69),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_76),
.A2(n_34),
.B1(n_37),
.B2(n_21),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_116),
.B1(n_82),
.B2(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_55),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_83),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_76),
.A2(n_55),
.B1(n_52),
.B2(n_42),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_109),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_124),
.B1(n_88),
.B2(n_91),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_62),
.B1(n_78),
.B2(n_44),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_83),
.B(n_78),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_109),
.B(n_90),
.Y(n_147)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_48),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_105),
.Y(n_141)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

BUFx2_ASAP7_75t_SL g139 ( 
.A(n_135),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_132),
.A2(n_98),
.B1(n_103),
.B2(n_86),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_140),
.B(n_149),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_132),
.A2(n_86),
.B1(n_97),
.B2(n_113),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_125),
.A2(n_97),
.B1(n_96),
.B2(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_125),
.A2(n_106),
.B1(n_104),
.B2(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_147),
.B1(n_126),
.B2(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_122),
.C(n_118),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_120),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_152),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_145),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_143),
.B1(n_142),
.B2(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_164),
.Y(n_174)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_138),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_163),
.B(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_173),
.B1(n_94),
.B2(n_62),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_126),
.C(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_102),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_171),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_147),
.B1(n_129),
.B2(n_122),
.C(n_141),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_163),
.B1(n_152),
.B2(n_156),
.C(n_154),
.Y(n_179)
);

XOR2x2_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_137),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_154),
.B(n_94),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_130),
.B1(n_131),
.B2(n_123),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_176),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_134),
.C(n_101),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_168),
.Y(n_189)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_158),
.CI(n_153),
.CON(n_178),
.SN(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_180),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_181),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_157),
.B(n_156),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_119),
.B(n_124),
.C(n_161),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_185),
.B1(n_59),
.B2(n_67),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_188),
.B1(n_166),
.B2(n_176),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_138),
.B1(n_135),
.B2(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_193),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_198),
.C(n_178),
.Y(n_203)
);

AO221x1_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_182),
.B1(n_188),
.B2(n_180),
.C(n_4),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_44),
.B(n_42),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_59),
.C(n_48),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_182),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_178),
.C(n_37),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_37),
.C(n_33),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

AOI321xp33_ASAP7_75t_L g206 ( 
.A1(n_200),
.A2(n_191),
.A3(n_192),
.B1(n_195),
.B2(n_197),
.C(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_79),
.Y(n_214)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_17),
.A3(n_16),
.B1(n_15),
.B2(n_13),
.C1(n_38),
.C2(n_33),
.Y(n_208)
);

AOI322xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_191),
.A3(n_17),
.B1(n_16),
.B2(n_38),
.C1(n_33),
.C2(n_7),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_7),
.C2(n_9),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_214),
.Y(n_217)
);

NOR2xp67_ASAP7_75t_SL g216 ( 
.A(n_209),
.B(n_213),
.Y(n_216)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_216),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_208),
.B(n_79),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_46),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_217),
.B(n_2),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_46),
.C1(n_215),
.C2(n_220),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_12),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_222),
.Y(n_225)
);


endmodule