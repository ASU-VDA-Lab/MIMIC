module fake_jpeg_13798_n_645 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_645);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_645;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx6p67_ASAP7_75t_R g165 ( 
.A(n_60),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_64),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_7),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_66),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_17),
.B(n_7),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_67),
.B(n_78),
.Y(n_156)
);

INVx11_ASAP7_75t_SL g68 ( 
.A(n_45),
.Y(n_68)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_75),
.Y(n_184)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_31),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_77),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_79),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_83),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_21),
.B(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_86),
.B(n_89),
.Y(n_183)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_88),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_9),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_9),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_92),
.B(n_95),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_26),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_59),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_37),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_97),
.B(n_98),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_26),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_100),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_101),
.Y(n_207)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_102),
.B(n_104),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_33),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_28),
.Y(n_108)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_6),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_116),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_38),
.Y(n_111)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_22),
.B(n_10),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_23),
.B(n_5),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_120),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_30),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_18),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_18),
.Y(n_125)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_122),
.A2(n_77),
.B1(n_79),
.B2(n_85),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_145),
.A2(n_174),
.B1(n_179),
.B2(n_125),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_60),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_152),
.B(n_182),
.Y(n_270)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_164),
.Y(n_209)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx2_ASAP7_75t_R g172 ( 
.A(n_83),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_172),
.B(n_178),
.Y(n_232)
);

AO22x2_ASAP7_75t_L g174 ( 
.A1(n_62),
.A2(n_57),
.B1(n_40),
.B2(n_50),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_63),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

AND2x4_ASAP7_75t_SL g178 ( 
.A(n_64),
.B(n_57),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_72),
.A2(n_27),
.B1(n_20),
.B2(n_58),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_180),
.Y(n_236)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_60),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_89),
.B(n_29),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_187),
.B(n_27),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_113),
.B(n_25),
.C(n_52),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_192),
.B(n_198),
.Y(n_247)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_108),
.Y(n_195)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_112),
.Y(n_201)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_68),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_205),
.Y(n_252)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_94),
.Y(n_204)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_94),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_211),
.B(n_263),
.Y(n_283)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_212),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_73),
.B1(n_75),
.B2(n_119),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_213),
.A2(n_239),
.B1(n_82),
.B2(n_193),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_46),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_214),
.B(n_219),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_215),
.A2(n_225),
.B1(n_245),
.B2(n_157),
.Y(n_284)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_197),
.Y(n_218)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_46),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_222),
.Y(n_304)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

BUFx24_ASAP7_75t_L g339 ( 
.A(n_223),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_188),
.A2(n_93),
.B1(n_114),
.B2(n_110),
.Y(n_225)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

INVx3_ASAP7_75t_SL g303 ( 
.A(n_226),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_229),
.Y(n_296)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_140),
.Y(n_231)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_127),
.A2(n_20),
.B1(n_123),
.B2(n_101),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_233),
.A2(n_248),
.B1(n_251),
.B2(n_259),
.Y(n_332)
);

BUFx16f_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_234),
.B(n_240),
.Y(n_294)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_143),
.Y(n_237)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_237),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_158),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_103),
.B1(n_99),
.B2(n_91),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_241),
.B(n_273),
.Y(n_328)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_146),
.Y(n_242)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_242),
.Y(n_298)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_156),
.Y(n_243)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_243),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_183),
.A2(n_81),
.B1(n_80),
.B2(n_74),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_177),
.A2(n_50),
.B1(n_47),
.B2(n_48),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_167),
.Y(n_249)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_250),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_128),
.A2(n_47),
.B1(n_48),
.B2(n_39),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_163),
.Y(n_254)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_142),
.Y(n_257)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_138),
.A2(n_47),
.B1(n_48),
.B2(n_39),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_189),
.Y(n_260)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_260),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_141),
.B(n_53),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_261),
.B(n_269),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_191),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_262),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_187),
.B(n_30),
.Y(n_263)
);

CKINVDCx9p33_ASAP7_75t_R g265 ( 
.A(n_169),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_265),
.B(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_130),
.Y(n_268)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_268),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_141),
.B(n_42),
.Y(n_269)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_142),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_272),
.B(n_280),
.Y(n_302)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_139),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_203),
.B(n_183),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_275),
.B(n_279),
.Y(n_293)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_148),
.Y(n_276)
);

INVx4_ASAP7_75t_SL g277 ( 
.A(n_169),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_278),
.Y(n_313)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_150),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_203),
.B(n_48),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_151),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_160),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_284),
.A2(n_287),
.B1(n_312),
.B2(n_323),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_213),
.A2(n_153),
.B1(n_179),
.B2(n_196),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_133),
.B(n_168),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_291),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_157),
.B1(n_166),
.B2(n_145),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g356 ( 
.A1(n_292),
.A2(n_320),
.B1(n_331),
.B2(n_235),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_306),
.A2(n_314),
.B1(n_315),
.B2(n_322),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_232),
.A2(n_133),
.B(n_178),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_318),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_247),
.A2(n_154),
.B1(n_136),
.B2(n_175),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_248),
.A2(n_199),
.B1(n_190),
.B2(n_132),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_233),
.A2(n_171),
.B1(n_147),
.B2(n_155),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_270),
.A2(n_58),
.B(n_51),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_237),
.A2(n_143),
.B1(n_147),
.B2(n_155),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_251),
.A2(n_199),
.B1(n_190),
.B2(n_131),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_226),
.A2(n_131),
.B1(n_185),
.B2(n_29),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_51),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_329),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_236),
.B(n_0),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_258),
.A2(n_135),
.B1(n_96),
.B2(n_165),
.Y(n_331)
);

AO21x2_ASAP7_75t_L g333 ( 
.A1(n_282),
.A2(n_96),
.B(n_134),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_333),
.A2(n_340),
.B1(n_217),
.B2(n_242),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_259),
.B(n_100),
.Y(n_337)
);

OAI21xp33_ASAP7_75t_L g380 ( 
.A1(n_337),
.A2(n_4),
.B(n_5),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_256),
.A2(n_47),
.B1(n_11),
.B2(n_3),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_264),
.B(n_0),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_0),
.Y(n_364)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_260),
.B1(n_250),
.B2(n_244),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_348),
.B1(n_352),
.B2(n_368),
.Y(n_391)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_342),
.Y(n_345)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_345),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_284),
.A2(n_267),
.B1(n_255),
.B2(n_224),
.Y(n_348)
);

INVx13_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_350),
.Y(n_398)
);

CKINVDCx10_ASAP7_75t_R g351 ( 
.A(n_339),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_351),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_314),
.A2(n_282),
.B1(n_253),
.B2(n_238),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_297),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_366),
.Y(n_396)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_356),
.B(n_361),
.Y(n_407)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_321),
.Y(n_357)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_357),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_249),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_364),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_338),
.B(n_209),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_360),
.B(n_362),
.Y(n_427)
);

INVx4_ASAP7_75t_SL g361 ( 
.A(n_339),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_208),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_296),
.B(n_220),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_363),
.B(n_371),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_220),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_367),
.Y(n_406)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_286),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_266),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_287),
.A2(n_231),
.B1(n_212),
.B2(n_271),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_327),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_373),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_283),
.B(n_266),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_372),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_1),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_308),
.B(n_12),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_376),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_316),
.B(n_302),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_334),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_377),
.A2(n_351),
.B1(n_309),
.B2(n_310),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_294),
.B(n_222),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_378),
.Y(n_409)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_383),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_4),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_381),
.A2(n_333),
.B1(n_303),
.B2(n_334),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_234),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_382),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_1),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_332),
.A2(n_257),
.B1(n_228),
.B2(n_227),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_384),
.A2(n_388),
.B1(n_286),
.B2(n_310),
.Y(n_402)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_312),
.B(n_277),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_305),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_324),
.B(n_1),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_386),
.B(n_387),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_300),
.B(n_227),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_291),
.A2(n_223),
.B1(n_5),
.B2(n_11),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_337),
.A2(n_4),
.B1(n_13),
.B2(n_16),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_389),
.A2(n_324),
.B1(n_333),
.B2(n_383),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_359),
.B(n_301),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_414),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_397),
.B(n_405),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_347),
.A2(n_346),
.B1(n_348),
.B2(n_370),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_400),
.B1(n_403),
.B2(n_415),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_347),
.A2(n_333),
.B1(n_340),
.B2(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_402),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_346),
.A2(n_333),
.B1(n_303),
.B2(n_336),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_404),
.A2(n_368),
.B1(n_358),
.B2(n_389),
.Y(n_452)
);

NOR2x1_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_286),
.Y(n_405)
);

INVx13_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_325),
.C(n_335),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_420),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_375),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_371),
.A2(n_336),
.B1(n_290),
.B2(n_311),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_419),
.A2(n_355),
.B(n_353),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_350),
.B(n_311),
.C(n_330),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_365),
.B(n_330),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_425),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_285),
.Y(n_425)
);

AO21x2_ASAP7_75t_SL g426 ( 
.A1(n_381),
.A2(n_295),
.B(n_304),
.Y(n_426)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_426),
.Y(n_436)
);

AOI21xp33_ASAP7_75t_L g448 ( 
.A1(n_429),
.A2(n_386),
.B(n_373),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_430),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_354),
.Y(n_434)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_409),
.B(n_374),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_435),
.B(n_448),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_405),
.A2(n_419),
.B(n_396),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_438),
.Y(n_491)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_395),
.Y(n_439)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_424),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_447),
.Y(n_469)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_425),
.Y(n_444)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_445),
.Y(n_495)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_446),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_411),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_451),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_399),
.A2(n_370),
.B1(n_385),
.B2(n_384),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_450),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_393),
.Y(n_451)
);

OAI22x1_ASAP7_75t_L g484 ( 
.A1(n_452),
.A2(n_402),
.B1(n_401),
.B2(n_398),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_427),
.B(n_345),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_453),
.B(n_413),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_422),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_454),
.B(n_455),
.Y(n_473)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_428),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_457),
.Y(n_489)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_428),
.Y(n_457)
);

NAND2x1_ASAP7_75t_SL g458 ( 
.A(n_398),
.B(n_361),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_458),
.A2(n_417),
.B(n_390),
.Y(n_468)
);

NOR2x1_ASAP7_75t_L g459 ( 
.A(n_394),
.B(n_369),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_459),
.A2(n_410),
.B(n_434),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_426),
.A2(n_358),
.B1(n_385),
.B2(n_356),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_462),
.Y(n_477)
);

INVx13_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_461),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_426),
.A2(n_356),
.B1(n_364),
.B2(n_377),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_400),
.A2(n_388),
.B1(n_356),
.B2(n_372),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_403),
.A2(n_379),
.B1(n_357),
.B2(n_343),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_407),
.A2(n_290),
.B1(n_295),
.B2(n_304),
.Y(n_465)
);

OAI32xp33_ASAP7_75t_L g466 ( 
.A1(n_406),
.A2(n_289),
.A3(n_285),
.B1(n_298),
.B2(n_299),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_460),
.Y(n_478)
);

XNOR2x1_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_414),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_467),
.B(n_479),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_468),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_412),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_470),
.B(n_474),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_392),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_410),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_482),
.Y(n_524)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_478),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_432),
.B(n_441),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_432),
.B(n_406),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_483),
.B(n_485),
.Y(n_512)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_484),
.Y(n_515)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_458),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_486),
.B(n_497),
.Y(n_501)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_394),
.B(n_407),
.C(n_423),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_459),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_422),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_401),
.Y(n_493)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_437),
.A2(n_426),
.B1(n_404),
.B2(n_416),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_496),
.A2(n_391),
.B1(n_443),
.B2(n_461),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_453),
.B(n_451),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_430),
.B(n_416),
.C(n_420),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_439),
.C(n_431),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g500 ( 
.A(n_435),
.B(n_413),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_500),
.B(n_423),
.Y(n_502)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_491),
.A2(n_437),
.B1(n_450),
.B2(n_440),
.Y(n_503)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_503),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_477),
.A2(n_440),
.B1(n_436),
.B2(n_447),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_504),
.A2(n_508),
.B1(n_487),
.B2(n_472),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_505),
.B(n_511),
.C(n_514),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_491),
.A2(n_452),
.B1(n_436),
.B2(n_462),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_506),
.A2(n_530),
.B1(n_468),
.B2(n_481),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_507),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_477),
.A2(n_431),
.B1(n_465),
.B2(n_443),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_493),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_509),
.B(n_522),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_445),
.C(n_446),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_470),
.B(n_407),
.C(n_455),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_478),
.A2(n_443),
.B(n_458),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_516),
.A2(n_489),
.B(n_472),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_466),
.Y(n_518)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_518),
.Y(n_541)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_471),
.Y(n_520)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_520),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_469),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_492),
.B(n_476),
.Y(n_523)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_523),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_471),
.B(n_449),
.Y(n_525)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_525),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_479),
.B(n_429),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_526),
.B(n_482),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_469),
.B(n_456),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_527),
.B(n_528),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_473),
.B(n_457),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_483),
.B(n_299),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_531),
.B(n_490),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_536),
.A2(n_521),
.B1(n_515),
.B2(n_504),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_555),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_475),
.C(n_467),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_539),
.B(n_542),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_521),
.A2(n_481),
.B(n_473),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_510),
.B(n_474),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_543),
.B(n_552),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_501),
.A2(n_480),
.B1(n_494),
.B2(n_495),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_545),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_501),
.B(n_494),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_546),
.B(n_549),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_484),
.C(n_496),
.Y(n_549)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_550),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_514),
.B(n_488),
.C(n_487),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_551),
.B(n_557),
.C(n_520),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_488),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_524),
.B(n_495),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_523),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g578 ( 
.A1(n_554),
.A2(n_556),
.B1(n_519),
.B2(n_509),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_508),
.A2(n_429),
.B1(n_461),
.B2(n_298),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_505),
.B(n_289),
.C(n_361),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_512),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_560),
.B(n_564),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_538),
.B(n_516),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_562),
.B(n_566),
.Y(n_583)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_535),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_563),
.B(n_576),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_552),
.B(n_529),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_534),
.A2(n_507),
.B(n_532),
.Y(n_566)
);

BUFx12_ASAP7_75t_L g567 ( 
.A(n_555),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_567),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_569),
.B(n_570),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_537),
.B(n_529),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_574),
.C(n_557),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_553),
.B(n_506),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_SL g585 ( 
.A(n_573),
.B(n_536),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_538),
.B(n_527),
.C(n_525),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_533),
.Y(n_575)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_575),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_502),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_547),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_578),
.A2(n_513),
.B1(n_548),
.B2(n_519),
.Y(n_591)
);

NOR2xp67_ASAP7_75t_SL g579 ( 
.A(n_539),
.B(n_526),
.Y(n_579)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_579),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_574),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_582),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_561),
.B(n_522),
.Y(n_581)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_581),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_568),
.A2(n_575),
.B1(n_541),
.B2(n_513),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_584),
.B(n_589),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_585),
.B(n_573),
.Y(n_609)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_591),
.Y(n_608)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_568),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_592),
.B(n_593),
.Y(n_603)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_569),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_572),
.B(n_549),
.C(n_554),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_595),
.B(n_559),
.C(n_571),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_558),
.B(n_540),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_596),
.B(n_562),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_565),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_599),
.B(n_601),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_594),
.B(n_559),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_592),
.A2(n_544),
.B1(n_535),
.B2(n_517),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_602),
.B(n_609),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_604),
.B(n_606),
.Y(n_613)
);

INVx13_ASAP7_75t_L g605 ( 
.A(n_581),
.Y(n_605)
);

AOI31xp67_ASAP7_75t_L g617 ( 
.A1(n_605),
.A2(n_567),
.A3(n_590),
.B(n_591),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_593),
.A2(n_515),
.B1(n_518),
.B2(n_517),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_610),
.A2(n_612),
.B1(n_590),
.B2(n_528),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_597),
.A2(n_542),
.B1(n_567),
.B2(n_560),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_611),
.A2(n_583),
.B(n_595),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_596),
.Y(n_612)
);

AOI21xp33_ASAP7_75t_L g629 ( 
.A1(n_614),
.A2(n_620),
.B(n_598),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_617),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_604),
.B(n_584),
.C(n_585),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_619),
.B(n_621),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_603),
.A2(n_588),
.B(n_586),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_607),
.A2(n_588),
.B1(n_586),
.B2(n_564),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_608),
.A2(n_530),
.B1(n_570),
.B2(n_556),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_622),
.B(n_609),
.Y(n_624)
);

NAND4xp25_ASAP7_75t_L g623 ( 
.A(n_600),
.B(n_349),
.C(n_319),
.D(n_309),
.Y(n_623)
);

INVx11_ASAP7_75t_L g628 ( 
.A(n_623),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_624),
.B(n_625),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_616),
.B(n_600),
.Y(n_625)
);

CKINVDCx14_ASAP7_75t_R g626 ( 
.A(n_613),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_618),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_629),
.A2(n_631),
.B(n_614),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_619),
.A2(n_598),
.B1(n_603),
.B2(n_606),
.Y(n_631)
);

NOR2x1_ASAP7_75t_L g632 ( 
.A(n_627),
.B(n_618),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_632),
.A2(n_633),
.B(n_634),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_630),
.A2(n_620),
.B(n_611),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_635),
.A2(n_628),
.B(n_605),
.Y(n_639)
);

OAI21xp33_ASAP7_75t_L g638 ( 
.A1(n_636),
.A2(n_628),
.B(n_630),
.Y(n_638)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_638),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_639),
.B(n_602),
.C(n_622),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_641),
.B(n_637),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_640),
.C(n_319),
.Y(n_643)
);

XNOR2xp5_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_223),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_13),
.B(n_16),
.Y(n_645)
);


endmodule