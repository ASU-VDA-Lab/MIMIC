module fake_jpeg_2739_n_96 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_96);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_96;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_29),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_34),
.C(n_31),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_32),
.B1(n_34),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_49),
.A2(n_35),
.B1(n_3),
.B2(n_4),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_29),
.Y(n_57)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_2),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_58),
.B(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_45),
.B1(n_43),
.B2(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_66),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_46),
.B1(n_35),
.B2(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_46),
.B1(n_35),
.B2(n_6),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_67),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_5),
.C(n_7),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_35),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_54),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_77),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_75),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_16),
.C(n_25),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_78),
.C(n_79),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_15),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_18),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_63),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_84),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_64),
.C(n_74),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_86),
.B1(n_65),
.B2(n_7),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_88),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_80),
.C(n_83),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_89),
.C(n_82),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_84),
.A3(n_88),
.B1(n_13),
.B2(n_14),
.C1(n_19),
.C2(n_20),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_11),
.C(n_21),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_22),
.B(n_24),
.C(n_26),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_10),
.Y(n_96)
);


endmodule