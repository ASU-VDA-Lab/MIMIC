module real_jpeg_14341_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_297, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_297;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_197;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_3),
.A2(n_22),
.B1(n_26),
.B2(n_99),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_3),
.A2(n_32),
.B1(n_36),
.B2(n_99),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_99),
.Y(n_175)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_32),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_6),
.A2(n_22),
.B1(n_26),
.B2(n_39),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_6),
.A2(n_39),
.B1(n_50),
.B2(n_51),
.Y(n_287)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_8),
.A2(n_32),
.B1(n_36),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_8),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_42),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_10),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_10),
.A2(n_27),
.B1(n_32),
.B2(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_10),
.A2(n_27),
.B1(n_56),
.B2(n_57),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_10),
.B(n_68),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_22),
.C(n_35),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_10),
.B(n_84),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_10),
.B(n_37),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_10),
.A2(n_57),
.B(n_70),
.C(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_10),
.B(n_55),
.Y(n_195)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_276),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_120),
.B(n_274),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_100),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_16),
.B(n_100),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_60),
.C(n_77),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_17),
.A2(n_18),
.B1(n_60),
.B2(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_43),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_19),
.A2(n_20),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_28),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_20),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_20),
.A2(n_44),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_20),
.B(n_178),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_20),
.A2(n_28),
.B1(n_44),
.B2(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_25),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_21),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_21),
.B(n_25),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_21),
.A2(n_209),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AO22x1_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_22),
.B(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_24),
.B(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_24),
.B(n_81),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_24),
.A2(n_80),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_27),
.A2(n_36),
.B(n_71),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_27),
.B(n_53),
.C(n_57),
.Y(n_207)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_28),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_38),
.B(n_40),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_29),
.A2(n_65),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_30),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_30),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_30),
.B(n_64),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_32),
.A2(n_36),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_32),
.B(n_145),
.Y(n_144)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_37),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_37),
.B(n_137),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_38),
.A2(n_62),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_40),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_40),
.B(n_148),
.Y(n_234)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_58),
.B(n_59),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_47),
.B(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_48),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_48),
.B(n_108),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_55),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_51),
.B(n_207),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_55),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_55),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_55),
.B(n_98),
.Y(n_215)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_58),
.A2(n_237),
.B(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_60),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_76),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_66),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_62),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_63),
.B(n_136),
.Y(n_185)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_72),
.Y(n_66)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_68),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_68),
.B(n_92),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_68),
.A2(n_91),
.B(n_92),
.Y(n_238)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_75),
.Y(n_88)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_72),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_72),
.B(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_73),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_103),
.B1(n_104),
.B2(n_119),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_76),
.B(n_101),
.C(n_103),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_77),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.C(n_93),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_78),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_79),
.B(n_85),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_80),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_87),
.A2(n_93),
.B1(n_94),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_87),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_88),
.B(n_191),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_90),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_97),
.B(n_107),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_111),
.B2(n_112),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_105),
.B(n_114),
.C(n_115),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_105),
.A2(n_106),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_110),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_118),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_113),
.A2(n_114),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_113),
.B(n_213),
.C(n_218),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_113),
.A2(n_114),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_115),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_268),
.B(n_273),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_255),
.B(n_267),
.Y(n_121)
);

AOI321xp33_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_221),
.A3(n_248),
.B1(n_253),
.B2(n_254),
.C(n_297),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_198),
.B(n_220),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_182),
.B(n_197),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_169),
.B(n_181),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_149),
.B(n_168),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_142),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_142),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B1(n_134),
.B2(n_141),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_139),
.C(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_162),
.B(n_167),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_157),
.B(n_161),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_156),
.B(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_160),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_165),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_171),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_196),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_196),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_187),
.C(n_189),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_194),
.C(n_195),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_200),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_211),
.B2(n_212),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_204),
.C(n_211),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_210),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_242),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_242),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_230),
.C(n_241),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.C(n_228),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_225),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_226),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_241),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_238),
.C(n_239),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_234),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_246),
.C(n_247),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_252),
.Y(n_253)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_257),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_264),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_264),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_294),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_279),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_288),
.B1(n_289),
.B2(n_293),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_286),
.Y(n_293)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);


endmodule