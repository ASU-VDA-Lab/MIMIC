module fake_jpeg_2699_n_236 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_236);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_235;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_60),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_86),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_79),
.B1(n_59),
.B2(n_61),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_66),
.B(n_76),
.C(n_57),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_70),
.B(n_68),
.C(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_58),
.B1(n_56),
.B2(n_78),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_102),
.B1(n_80),
.B2(n_85),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_72),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_59),
.B1(n_78),
.B2(n_55),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_96),
.B1(n_99),
.B2(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_80),
.B1(n_72),
.B2(n_73),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_79),
.B1(n_62),
.B2(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_71),
.B1(n_62),
.B2(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_119),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_81),
.B1(n_101),
.B2(n_75),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_116),
.B1(n_120),
.B2(n_83),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_114),
.Y(n_132)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_112),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_63),
.C(n_65),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_84),
.B1(n_83),
.B2(n_64),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_53),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_118),
.B(n_122),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_75),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_85),
.B1(n_84),
.B2(n_64),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_83),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_123),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_45),
.B1(n_44),
.B2(n_42),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_128),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_64),
.B1(n_22),
.B2(n_24),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_129),
.B1(n_130),
.B2(n_138),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_108),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_142),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_1),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_52),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_144),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_3),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_3),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_4),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_111),
.B(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_145),
.B(n_5),
.Y(n_151)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_146),
.B1(n_130),
.B2(n_132),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_149),
.A2(n_165),
.B(n_12),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_109),
.C(n_120),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_156),
.C(n_131),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_5),
.Y(n_154)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_6),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_26),
.C(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_140),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_160),
.A2(n_161),
.B(n_162),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_8),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_137),
.B(n_9),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_28),
.B1(n_48),
.B2(n_47),
.Y(n_165)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

AOI21x1_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_51),
.B(n_46),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_170),
.B(n_37),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_169),
.A2(n_171),
.B1(n_131),
.B2(n_10),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_182),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_127),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_181),
.C(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_177),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_36),
.B(n_35),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_167),
.B(n_156),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_30),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_9),
.B(n_12),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_20),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_192),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_13),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_194),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_147),
.A2(n_15),
.B(n_16),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_16),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_205),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_181),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_200),
.Y(n_208)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_152),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_212),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_173),
.C(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_189),
.C(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_194),
.C(n_184),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_163),
.B(n_196),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_185),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_206),
.B1(n_203),
.B2(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_220),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_198),
.B(n_161),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_214),
.C(n_191),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_165),
.B1(n_215),
.B2(n_208),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_195),
.B1(n_171),
.B2(n_217),
.Y(n_226)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_218),
.Y(n_229)
);

FAx1_ASAP7_75t_SL g230 ( 
.A(n_229),
.B(n_225),
.CI(n_224),
.CON(n_230),
.SN(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_230),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_232),
.A2(n_227),
.B(n_230),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_233),
.Y(n_234)
);

OAI321xp33_ASAP7_75t_L g235 ( 
.A1(n_234),
.A2(n_183),
.A3(n_221),
.B1(n_166),
.B2(n_19),
.C(n_17),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_235),
.B(n_17),
.Y(n_236)
);


endmodule