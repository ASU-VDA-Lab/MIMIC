module real_jpeg_18085_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_43;
wire n_8;
wire n_54;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_47;
wire n_51;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_18),
.Y(n_17)
);

AND2x2_ASAP7_75t_SL g34 ( 
.A(n_5),
.B(n_20),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_43),
.Y(n_6)
);

MAJIxp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_31),
.C(n_32),
.Y(n_7)
);

OAI21xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_16),
.B(n_26),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_9),
.A2(n_10),
.B1(n_36),
.B2(n_41),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_34),
.C(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_15),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_15),
.B(n_36),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_20),
.B(n_25),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_20),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);


endmodule