module fake_jpeg_27212_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_51),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_26),
.B(n_24),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_15),
.B(n_4),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_21),
.B(n_26),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_14),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_49),
.B(n_52),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_32),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_28),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_17),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_64),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_61),
.B(n_69),
.C(n_70),
.Y(n_94)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_14),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_72),
.Y(n_80)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_16),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_35),
.B1(n_36),
.B2(n_0),
.Y(n_69)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_1),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_15),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_10),
.B(n_11),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_91),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_57),
.C(n_41),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_92),
.C(n_71),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_57),
.C(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_9),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_70),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_72),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_104),
.C(n_105),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_79),
.C(n_65),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_10),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_94),
.B1(n_80),
.B2(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_114),
.B1(n_95),
.B2(n_102),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_89),
.C(n_86),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_69),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_76),
.B1(n_56),
.B2(n_42),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_100),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_117),
.B(n_63),
.CI(n_67),
.CON(n_123),
.SN(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_121),
.B(n_107),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_121),
.C(n_117),
.Y(n_125)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_110),
.B(n_59),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_125),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_120),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_121),
.B(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_89),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_125),
.C(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_128),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_130),
.B(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_56),
.Y(n_137)
);


endmodule