module real_jpeg_8897_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_326, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_326;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_1),
.A2(n_37),
.B1(n_67),
.B2(n_68),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_67),
.B1(n_68),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_2),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_141),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_141),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_141),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_3),
.A2(n_12),
.B(n_28),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_4),
.A2(n_67),
.B1(n_68),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_4),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_105),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_105),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_105),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_5),
.A2(n_61),
.B1(n_67),
.B2(n_68),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_61),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_61),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_9),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_27),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_67),
.B1(n_68),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_11),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_100),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_100),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_100),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_31),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_12),
.B(n_31),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_12),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_12),
.A2(n_27),
.B(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_12),
.B(n_27),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_12),
.B(n_52),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_125),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_13),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_13),
.A2(n_67),
.B1(n_68),
.B2(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_112),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_112),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_14),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_14),
.A2(n_67),
.B1(n_68),
.B2(n_80),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_80),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_16),
.A2(n_44),
.B1(n_67),
.B2(n_68),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_42),
.B1(n_43),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_17),
.A2(n_51),
.B1(n_67),
.B2(n_68),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_17),
.A2(n_31),
.B1(n_32),
.B2(n_51),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_86),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_72),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_53),
.B1(n_54),
.B2(n_71),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_34),
.B(n_35),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_25),
.A2(n_34),
.B1(n_85),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_26),
.A2(n_30),
.B1(n_57),
.B2(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_26),
.A2(n_30),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_26),
.A2(n_30),
.B1(n_151),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_26),
.A2(n_30),
.B1(n_167),
.B2(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_26),
.A2(n_30),
.B1(n_207),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_26),
.A2(n_30),
.B1(n_218),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_26),
.A2(n_30),
.B1(n_244),
.B2(n_262),
.Y(n_261)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_29),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_30),
.B(n_125),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_SL g63 ( 
.A1(n_31),
.A2(n_64),
.B(n_65),
.C(n_66),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_31),
.B(n_33),
.Y(n_155)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_32),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_46),
.B1(n_49),
.B2(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_47),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_43),
.A2(n_47),
.B(n_125),
.C(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_45),
.A2(n_52),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_49),
.B1(n_60),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_46),
.A2(n_49),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_46),
.A2(n_49),
.B1(n_222),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_46),
.A2(n_49),
.B1(n_247),
.B2(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_46),
.A2(n_49),
.B1(n_79),
.B2(n_265),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.C(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_62),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_66),
.B(n_70),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_66),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_63),
.A2(n_66),
.B1(n_111),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_63),
.A2(n_66),
.B1(n_138),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_63),
.A2(n_66),
.B1(n_147),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_63),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_63),
.A2(n_66),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_63),
.A2(n_66),
.B1(n_230),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_63),
.A2(n_66),
.B1(n_239),
.B2(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_66),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_67),
.B(n_69),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_67),
.B(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_68),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_70),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.C(n_81),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_310),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_78),
.C(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_78),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_78),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_81),
.B(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI321xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_307),
.A3(n_317),
.B1(n_322),
.B2(n_323),
.C(n_325),
.Y(n_88)
);

AOI321xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_255),
.A3(n_295),
.B1(n_301),
.B2(n_306),
.C(n_326),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_212),
.C(n_251),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_182),
.B(n_211),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_161),
.B(n_181),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_143),
.B(n_160),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_132),
.B(n_142),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_118),
.B(n_131),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_106),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_101),
.A2(n_102),
.B1(n_159),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_104),
.A2(n_122),
.B1(n_123),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_113),
.B2(n_117),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_126),
.B(n_130),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_124),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_123),
.B1(n_140),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_122),
.A2(n_123),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_122),
.A2(n_123),
.B1(n_193),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_122),
.A2(n_123),
.B1(n_227),
.B2(n_237),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_122),
.A2(n_123),
.B(n_237),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_134),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_137),
.C(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_144),
.B(n_145),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.CI(n_152),
.CON(n_145),
.SN(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_157),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_174),
.B2(n_175),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_177),
.C(n_179),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_173),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_166),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_171),
.C(n_173),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_176),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_183),
.B(n_184),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_197),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_186),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_186),
.B(n_196),
.C(n_197),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_187),
.B(n_191),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_194),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_208),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_205),
.B2(n_206),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_205),
.C(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_202),
.A2(n_204),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g302 ( 
.A1(n_213),
.A2(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_232),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_214),
.B(n_232),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_225),
.C(n_231),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_224),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_219),
.B1(n_220),
.B2(n_223),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_217),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_SL g249 ( 
.A(n_219),
.B(n_223),
.C(n_224),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_231),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_228),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_249),
.B2(n_250),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_235),
.B(n_240),
.C(n_250),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_238),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_245),
.C(n_248),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_245),
.B1(n_246),
.B2(n_248),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_243),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_253),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_274),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_256),
.B(n_274),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_267),
.C(n_273),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_258),
.B1(n_267),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_263),
.C(n_266),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_261),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_262),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_267),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_269),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_289),
.B(n_291),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_270),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_270),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_271),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_293),
.B2(n_294),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_286),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_286),
.C(n_294),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_282),
.B(n_284),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_282),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_284),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_284),
.A2(n_309),
.B1(n_313),
.B2(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_292),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_298),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_315),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_315),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_313),
.C(n_314),
.Y(n_308)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_309),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_319),
.Y(n_322)
);


endmodule