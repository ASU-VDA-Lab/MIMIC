module fake_jpeg_17098_n_185 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_35),
.B(n_37),
.Y(n_70)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_1),
.C(n_2),
.Y(n_39)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_39),
.B(n_4),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_46),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_17),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_47),
.B1(n_15),
.B2(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_1),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_33),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_58),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_33),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_66),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_26),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_77),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_67),
.B(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_37),
.B(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_25),
.C(n_31),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_83),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_66),
.A2(n_27),
.B1(n_22),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_82),
.A2(n_102),
.B1(n_12),
.B2(n_14),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_42),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_70),
.B(n_51),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_89),
.A2(n_96),
.B1(n_92),
.B2(n_100),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_61),
.Y(n_90)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_36),
.B1(n_29),
.B2(n_28),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_96),
.B1(n_78),
.B2(n_68),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_54),
.B(n_6),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_7),
.B(n_71),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_20),
.B1(n_31),
.B2(n_6),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_9),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_12),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_58),
.CI(n_54),
.CON(n_104),
.SN(n_104)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_112),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_74),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_114),
.B1(n_93),
.B2(n_100),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_62),
.B1(n_75),
.B2(n_52),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_77),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_84),
.B(n_52),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_69),
.C(n_75),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_114),
.C(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_69),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_117),
.B(n_118),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_133),
.B1(n_127),
.B2(n_131),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_84),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_131),
.C(n_134),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_91),
.B(n_97),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_97),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_104),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_101),
.CON(n_138),
.SN(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_110),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_138),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_152),
.B1(n_137),
.B2(n_129),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_110),
.B(n_105),
.C(n_122),
.D(n_84),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_127),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_121),
.A3(n_82),
.B1(n_86),
.B2(n_113),
.C1(n_90),
.C2(n_106),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_134),
.C(n_126),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_159),
.C(n_141),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_157),
.A2(n_143),
.B1(n_128),
.B2(n_141),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_160),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_133),
.C(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_130),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_106),
.C(n_144),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_160),
.A2(n_143),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_152),
.C(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_168),
.B(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_173),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_162),
.B1(n_161),
.B2(n_137),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_174),
.B1(n_173),
.B2(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_177),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_158),
.C(n_108),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_170),
.A2(n_149),
.B(n_153),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_111),
.A3(n_102),
.B1(n_94),
.B2(n_95),
.C1(n_98),
.C2(n_88),
.Y(n_180)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_111),
.B(n_115),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_95),
.C(n_98),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_181),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_184),
.B(n_183),
.Y(n_185)
);


endmodule