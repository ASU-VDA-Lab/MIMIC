module fake_jpeg_26312_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_23),
.B(n_30),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_30),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_23),
.B1(n_30),
.B2(n_25),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_39),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_54),
.Y(n_82)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_16),
.B1(n_24),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_44),
.B1(n_16),
.B2(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_43),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_16),
.B1(n_24),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_16),
.B1(n_44),
.B2(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_57),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_59),
.Y(n_74)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_38),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_70),
.B(n_71),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_78),
.B1(n_68),
.B2(n_46),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_18),
.B(n_33),
.C(n_25),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_75),
.A2(n_18),
.A3(n_33),
.B1(n_20),
.B2(n_32),
.Y(n_113)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_16),
.B1(n_37),
.B2(n_41),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_23),
.B(n_22),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_87),
.B1(n_98),
.B2(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_40),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_90),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_21),
.B1(n_19),
.B2(n_24),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_39),
.Y(n_118)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_51),
.B(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_95),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_92),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_24),
.B1(n_26),
.B2(n_21),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_45),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_40),
.C(n_38),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_94),
.B(n_39),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_32),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_102),
.Y(n_114)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_46),
.A2(n_27),
.B1(n_28),
.B2(n_20),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_110),
.B1(n_112),
.B2(n_93),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_71),
.A2(n_61),
.B1(n_50),
.B2(n_48),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_109),
.B1(n_78),
.B2(n_73),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_48),
.B1(n_67),
.B2(n_63),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_27),
.B1(n_28),
.B2(n_67),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_70),
.A2(n_27),
.B1(n_28),
.B2(n_19),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_125),
.Y(n_151)
);

NAND3xp33_ASAP7_75t_SL g115 ( 
.A(n_74),
.B(n_38),
.C(n_34),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_45),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_120),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_19),
.B1(n_21),
.B2(n_26),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_119),
.A2(n_84),
.B1(n_29),
.B2(n_89),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_20),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_33),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_26),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_27),
.B1(n_18),
.B2(n_25),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_126),
.A2(n_95),
.B1(n_90),
.B2(n_74),
.Y(n_136)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_99),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_72),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_132),
.B(n_29),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_136),
.B1(n_142),
.B2(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_134),
.B(n_140),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_107),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_138),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_121),
.B(n_80),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_139),
.A2(n_29),
.B(n_22),
.Y(n_184)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_153),
.Y(n_163)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_143),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_85),
.B1(n_94),
.B2(n_86),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_157),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_105),
.A2(n_75),
.A3(n_86),
.B1(n_77),
.B2(n_102),
.Y(n_146)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_150),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_107),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_149),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_122),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_75),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_77),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_159),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_103),
.A2(n_73),
.B1(n_96),
.B2(n_91),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_162),
.B1(n_22),
.B2(n_31),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_158),
.B1(n_124),
.B2(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_97),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_83),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_83),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_106),
.A2(n_83),
.B1(n_88),
.B2(n_22),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_107),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_167),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_120),
.C(n_106),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_177),
.C(n_182),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_126),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_133),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_178),
.B1(n_188),
.B2(n_195),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_117),
.C(n_113),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_146),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_117),
.C(n_124),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_161),
.A2(n_128),
.B1(n_22),
.B2(n_31),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_0),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_186),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_180),
.A2(n_152),
.B(n_134),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_144),
.C(n_139),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_187),
.B(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_0),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_1),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_22),
.B1(n_31),
.B2(n_9),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_196),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_139),
.B(n_31),
.C(n_8),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_151),
.C(n_131),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_1),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_141),
.Y(n_200)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_201),
.B(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_192),
.Y(n_202)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_209),
.Y(n_239)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_210),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_142),
.B(n_152),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_218),
.B(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_216),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_175),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_171),
.A2(n_153),
.B(n_154),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_223),
.B(n_194),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_162),
.B1(n_131),
.B2(n_143),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_181),
.B1(n_189),
.B2(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_145),
.C(n_143),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_182),
.C(n_176),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_171),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_187),
.A2(n_2),
.B(n_3),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_193),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_224),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_235),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_229),
.B(n_199),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_198),
.C(n_221),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_232),
.A2(n_243),
.B1(n_187),
.B2(n_194),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_163),
.C(n_173),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g269 ( 
.A(n_233),
.B(n_11),
.C(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_204),
.B1(n_205),
.B2(n_213),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_208),
.B1(n_210),
.B2(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_240),
.B(n_245),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_163),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_241),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_181),
.B1(n_168),
.B2(n_193),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_212),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_201),
.B(n_172),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_197),
.B1(n_168),
.B2(n_218),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_248),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_190),
.B(n_10),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_254),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_258),
.B1(n_261),
.B2(n_267),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_243),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_229),
.B(n_219),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_257),
.B1(n_268),
.B2(n_236),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_232),
.A2(n_203),
.B1(n_211),
.B2(n_207),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_207),
.B1(n_222),
.B2(n_198),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_269),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_172),
.B1(n_197),
.B2(n_191),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_199),
.C(n_180),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_264),
.C(n_239),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_180),
.C(n_223),
.Y(n_264)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_236),
.A2(n_190),
.B1(n_4),
.B2(n_5),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_247),
.A2(n_15),
.B1(n_13),
.B2(n_11),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_275),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_227),
.B(n_231),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_269),
.B(n_234),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_239),
.C(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_280),
.C(n_284),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_231),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_281),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_252),
.B1(n_267),
.B2(n_255),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_260),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_244),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_245),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_244),
.C(n_248),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_257),
.A2(n_228),
.B1(n_234),
.B2(n_226),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_266),
.B1(n_263),
.B2(n_250),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_292),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_274),
.A2(n_256),
.B1(n_254),
.B2(n_228),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_299),
.B(n_7),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_294),
.B(n_298),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_6),
.B(n_7),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_3),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_6),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_251),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_277),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_295),
.B(n_273),
.C(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_305),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_275),
.Y(n_303)
);

AOI31xp67_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_291),
.A3(n_293),
.B(n_294),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_3),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_287),
.C(n_290),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_306),
.B(n_308),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_6),
.Y(n_312)
);

NAND3xp33_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_298),
.C(n_292),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_318),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_317),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_306),
.C(n_305),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_307),
.C(n_301),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_286),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

AOI21x1_ASAP7_75t_SL g324 ( 
.A1(n_320),
.A2(n_321),
.B(n_323),
.Y(n_324)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_315),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_311),
.B(n_323),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_320),
.Y(n_327)
);

NOR3xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_325),
.C(n_316),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_322),
.Y(n_329)
);


endmodule