module fake_jpeg_16762_n_162 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_162);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_33),
.B(n_37),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_16),
.A2(n_15),
.B1(n_28),
.B2(n_22),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_36),
.A2(n_45),
.B1(n_31),
.B2(n_11),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_46),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_16),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_4),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_15),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_14),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_23),
.B(n_7),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_20),
.Y(n_55)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_82),
.B1(n_34),
.B2(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_63),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_29),
.C(n_14),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_12),
.C(n_64),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_73),
.B(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_31),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_31),
.B(n_10),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_38),
.C(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_8),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_67),
.B1(n_59),
.B2(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_8),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_57),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_89),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_95),
.C(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_94),
.B1(n_97),
.B2(n_102),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_51),
.B(n_34),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_94),
.B(n_54),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_99),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_93),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_54),
.A2(n_43),
.B1(n_51),
.B2(n_39),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_96),
.B1(n_102),
.B2(n_101),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_68),
.A2(n_80),
.B1(n_77),
.B2(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_95),
.B1(n_96),
.B2(n_87),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_56),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_101),
.Y(n_108)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_81),
.B1(n_78),
.B2(n_61),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_62),
.C(n_78),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_61),
.C(n_56),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_118),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_69),
.C(n_62),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_113),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_121),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_103),
.C(n_83),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_92),
.C(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_104),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_131),
.Y(n_137)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_90),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_115),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_139),
.C(n_128),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_111),
.C(n_121),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_118),
.B1(n_106),
.B2(n_105),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_140),
.A2(n_142),
.B1(n_137),
.B2(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_127),
.B1(n_124),
.B2(n_128),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_133),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_146),
.B(n_150),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_134),
.B(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_140),
.C(n_150),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_139),
.CI(n_136),
.CON(n_150),
.SN(n_150)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_145),
.B1(n_147),
.B2(n_151),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_155),
.B(n_152),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_153),
.B(n_158),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_157),
.Y(n_162)
);


endmodule