module real_jpeg_26096_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_1),
.A2(n_56),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_60),
.B1(n_65),
.B2(n_70),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_1),
.A2(n_36),
.B1(n_38),
.B2(n_70),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_1),
.A2(n_26),
.B1(n_30),
.B2(n_70),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_2),
.A2(n_54),
.B1(n_73),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_60),
.B1(n_65),
.B2(n_108),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_2),
.A2(n_36),
.B1(n_38),
.B2(n_108),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_108),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_73),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_3),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_3),
.B(n_59),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_3),
.B(n_36),
.C(n_80),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_3),
.A2(n_60),
.B1(n_65),
.B2(n_200),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_3),
.B(n_123),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_3),
.A2(n_36),
.B1(n_38),
.B2(n_200),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_3),
.B(n_26),
.C(n_41),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_3),
.A2(n_25),
.B(n_262),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_60),
.B1(n_65),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_7),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_7),
.A2(n_36),
.B1(n_38),
.B2(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_54),
.B1(n_55),
.B2(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_7),
.A2(n_26),
.B1(n_30),
.B2(n_84),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_36),
.B1(n_38),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_9),
.A2(n_46),
.B1(n_60),
.B2(n_65),
.Y(n_125)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_11),
.A2(n_56),
.B1(n_73),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_11),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_11),
.A2(n_60),
.B1(n_65),
.B2(n_145),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_11),
.A2(n_36),
.B1(n_38),
.B2(n_145),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_11),
.A2(n_26),
.B1(n_30),
.B2(n_145),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_12),
.A2(n_35),
.B1(n_60),
.B2(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_13),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_13),
.A2(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_57),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_13),
.A2(n_26),
.B1(n_30),
.B2(n_57),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_15),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_15),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_89)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_16),
.Y(n_174)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_16),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_16),
.A2(n_170),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_135),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_133),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_21),
.B(n_112),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_22),
.A2(n_75),
.B1(n_76),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_22),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_23),
.A2(n_24),
.B(n_50),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_24),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_24),
.A2(n_32),
.B1(n_33),
.B2(n_49),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_29),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_29),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_25),
.A2(n_27),
.B1(n_96),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_25),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_25),
.A2(n_172),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_25),
.B(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_25),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_30),
.B1(n_41),
.B2(n_43),
.Y(n_44)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_28),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_28),
.B(n_200),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_30),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_34),
.A2(n_39),
.B1(n_47),
.B2(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_36),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_36),
.A2(n_38),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_36),
.B(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_39),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_39),
.A2(n_47),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_39),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_39),
.A2(n_47),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.Y(n_39)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_44),
.A2(n_87),
.B1(n_102),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_44),
.A2(n_155),
.B(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_44),
.A2(n_193),
.B(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_44),
.B(n_200),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_47),
.B(n_194),
.Y(n_250)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B(n_66),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_52),
.A2(n_58),
.B1(n_109),
.B2(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI32xp33_ASAP7_75t_L g166 ( 
.A1(n_54),
.A2(n_63),
.A3(n_65),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_55),
.Y(n_199)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_68),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_58),
.A2(n_66),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_59),
.A2(n_71),
.B1(n_107),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_65),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_60),
.B(n_64),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_60),
.B(n_225),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_71),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_71),
.A2(n_111),
.B(n_196),
.Y(n_195)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_78),
.A2(n_162),
.B(n_164),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g238 ( 
.A1(n_78),
.A2(n_164),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_79),
.A2(n_104),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_79),
.A2(n_148),
.B(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_87),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_87),
.A2(n_250),
.B(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_89),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_91),
.A2(n_92),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.C(n_105),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_93),
.A2(n_94),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_95),
.Y(n_157)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_103),
.B(n_105),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_110),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_130),
.B2(n_132),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_122),
.A2(n_123),
.B1(n_163),
.B2(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_123),
.B(n_149),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_311),
.B(n_317),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_182),
.B(n_310),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_175),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_138),
.B(n_175),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_156),
.C(n_158),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_139),
.A2(n_140),
.B1(n_156),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_150),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_146),
.C(n_150),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_151),
.B(n_154),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_156),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_158),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_165),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_161),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_165),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_169),
.Y(n_202)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_174),
.A2(n_275),
.B(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_177),
.B(n_178),
.C(n_181),
.Y(n_316)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_217),
.B(n_304),
.C(n_309),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_211),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_211),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_202),
.C(n_203),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_185),
.A2(n_186),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_191),
.C(n_195),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_190),
.Y(n_205)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_200),
.B(n_201),
.Y(n_196)
);

INVx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_202),
.B(n_203),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_298),
.B(n_303),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_251),
.B(n_297),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_240),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_222),
.B(n_240),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.C(n_237),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_223),
.B(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_226),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B(n_231),
.Y(n_226)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_231),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_233),
.A2(n_237),
.B1(n_238),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_233),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_241),
.B(n_247),
.C(n_248),
.Y(n_302)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_291),
.B(n_296),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_271),
.B(n_290),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_265),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_259),
.C(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_269),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_279),
.B(n_289),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_284),
.B(n_288),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_295),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);


endmodule