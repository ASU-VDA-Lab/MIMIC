module fake_jpeg_7906_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_1),
.C(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_47),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_30),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_28),
.B1(n_29),
.B2(n_25),
.Y(n_58)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_46),
.B1(n_50),
.B2(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_32),
.A2(n_28),
.B1(n_29),
.B2(n_25),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_62),
.B1(n_72),
.B2(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_28),
.B1(n_23),
.B2(n_14),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_67),
.B1(n_15),
.B2(n_22),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_30),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_63),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_39),
.B1(n_34),
.B2(n_19),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_19),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_15),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_34),
.B(n_39),
.C(n_23),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_41),
.B1(n_55),
.B2(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_33),
.B1(n_32),
.B2(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_20),
.B1(n_17),
.B2(n_22),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_57),
.B1(n_60),
.B2(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_31),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_89),
.C(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_86),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_86),
.B1(n_89),
.B2(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_41),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_88),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_21),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_19),
.C(n_34),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_58),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_38),
.C(n_34),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_99),
.B(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_68),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_73),
.B(n_65),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_3),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_64),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_98),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_106),
.B1(n_77),
.B2(n_82),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_56),
.B1(n_33),
.B2(n_47),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_70),
.B1(n_49),
.B2(n_43),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_81),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_113),
.C(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_94),
.A2(n_84),
.B1(n_80),
.B2(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_4),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_121),
.C(n_4),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_118),
.B(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_99),
.B1(n_107),
.B2(n_105),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_106),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_21),
.B(n_5),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_126),
.B1(n_130),
.B2(n_132),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_129),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_92),
.B1(n_102),
.B2(n_96),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_115),
.C(n_92),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_120),
.C(n_116),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_104),
.B(n_96),
.C(n_76),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_139),
.C(n_127),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_131),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_143),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_134),
.B(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_137),
.B(n_142),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_113),
.C(n_116),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_126),
.B(n_113),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_127),
.CI(n_123),
.CON(n_146),
.SN(n_146)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_129),
.B(n_13),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_70),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_144),
.A2(n_69),
.B1(n_49),
.B2(n_7),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_148),
.C(n_144),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_146),
.A2(n_150),
.B1(n_6),
.B2(n_8),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_123),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_149),
.B(n_6),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_132),
.C(n_69),
.Y(n_148)
);

NAND4xp25_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_69),
.C(n_49),
.D(n_7),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_154),
.C(n_156),
.Y(n_160)
);

AOI31xp67_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_5),
.A3(n_6),
.B(n_7),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_8),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_49),
.Y(n_156)
);

NOR5xp2_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_158),
.C(n_8),
.D(n_9),
.E(n_11),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_152),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

AOI21x1_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_162),
.B(n_11),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_147),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_147),
.C(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_166),
.Y(n_167)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_159),
.B(n_146),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_160),
.B(n_12),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_167),
.Y(n_170)
);


endmodule