module real_jpeg_28134_n_18 (n_17, n_8, n_0, n_2, n_331, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_331;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_1),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_46),
.B(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_1),
.B(n_48),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_1),
.A2(n_62),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_1),
.B(n_62),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_103),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_1),
.A2(n_26),
.B1(n_34),
.B2(n_237),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_1),
.A2(n_49),
.B(n_253),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_36),
.B1(n_62),
.B2(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_2),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_131)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_4),
.A2(n_54),
.B1(n_62),
.B2(n_63),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_5),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_49),
.B1(n_50),
.B2(n_106),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_106),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_106),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_8),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_49),
.B1(n_50),
.B2(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_65),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_9),
.A2(n_62),
.B1(n_63),
.B2(n_87),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_87),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_87),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_10),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_156),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_10),
.A2(n_62),
.B1(n_63),
.B2(n_156),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_156),
.Y(n_237)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_11),
.A2(n_29),
.A3(n_62),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_12),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_145),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_145),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_145),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_13),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_13),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_226)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_16),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_16),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_16),
.A2(n_28),
.B1(n_29),
.B2(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_16),
.A2(n_49),
.B1(n_50),
.B2(n_74),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_16),
.A2(n_42),
.B1(n_43),
.B2(n_74),
.Y(n_322)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_17),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_310),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_121),
.A3(n_135),
.B1(n_308),
.B2(n_309),
.C(n_330),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_107),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_21),
.B(n_107),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_77),
.C(n_92),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_22),
.B(n_77),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_56),
.B1(n_57),
.B2(n_76),
.Y(n_22)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_37),
.B2(n_38),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_24),
.A2(n_38),
.B(n_56),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_25),
.B(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_35),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_26),
.A2(n_35),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_26),
.A2(n_96),
.B1(n_97),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_26),
.A2(n_32),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_26),
.A2(n_32),
.B1(n_231),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_26),
.A2(n_97),
.B1(n_226),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_27),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_33),
.B1(n_161),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_27),
.A2(n_33),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_28),
.A2(n_29),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_28),
.B(n_70),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_28),
.B(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_53),
.B2(n_55),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_40),
.A2(n_45),
.B1(n_48),
.B2(n_105),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_42),
.A2(n_52),
.B(n_154),
.C(n_159),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_46),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_44),
.A2(n_53),
.B1(n_55),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_44),
.A2(n_55),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_44),
.A2(n_55),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_45),
.A2(n_48),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_45),
.A2(n_48),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_45),
.A2(n_48),
.B1(n_105),
.B2(n_185),
.Y(n_199)
);

AO22x1_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_48)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_80),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g261 ( 
.A1(n_49),
.A2(n_63),
.A3(n_80),
.B1(n_254),
.B2(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_50),
.B(n_154),
.Y(n_254)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_66),
.B1(n_72),
.B2(n_75),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_67),
.B1(n_68),
.B2(n_99),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_62),
.B(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_66),
.A2(n_75),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_66),
.A2(n_75),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_67),
.A2(n_68),
.B1(n_73),
.B2(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_67),
.A2(n_68),
.B(n_90),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_67),
.A2(n_68),
.B1(n_99),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_67),
.A2(n_68),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_67),
.A2(n_68),
.B1(n_212),
.B2(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_67),
.A2(n_68),
.B1(n_150),
.B2(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_68),
.B(n_154),
.Y(n_238)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_91),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_85),
.B2(n_88),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_79),
.A2(n_83),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_79),
.A2(n_83),
.B1(n_146),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_79),
.A2(n_83),
.B1(n_168),
.B2(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_79),
.A2(n_83),
.B(n_318),
.Y(n_317)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_80),
.Y(n_263)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_88),
.Y(n_114)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_108),
.CI(n_120),
.CON(n_107),
.SN(n_107)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_108),
.C(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_92),
.A2(n_93),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.C(n_104),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_94),
.B(n_100),
.CI(n_104),
.CON(n_291),
.SN(n_291)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_95),
.B(n_98),
.Y(n_195)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_188),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_103),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_103),
.B1(n_115),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_102),
.A2(n_103),
.B1(n_144),
.B2(n_167),
.Y(n_166)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_107),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_119),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_109),
.A2(n_110),
.B1(n_125),
.B2(n_133),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_113),
.C(n_118),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_110),
.B(n_133),
.C(n_134),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_116),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_118),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_116),
.B(n_126),
.C(n_130),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_122),
.B(n_123),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_134),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_128),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_131),
.Y(n_318)
);

AOI321xp33_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_289),
.A3(n_297),
.B1(n_302),
.B2(n_307),
.C(n_331),
.Y(n_135)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_190),
.C(n_202),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_172),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_138),
.B(n_172),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_157),
.C(n_164),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_139),
.B(n_286),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_147),
.B2(n_148),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_148),
.C(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_154),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_157),
.A2(n_164),
.B1(n_165),
.B2(n_287),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_157),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_160),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_163),
.Y(n_178)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_166),
.B(n_274),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_169),
.B(n_171),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_170),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_180),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_179),
.C(n_180),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_177),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_186),
.C(n_189),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_191),
.A2(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_192),
.B(n_193),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_195),
.B(n_196),
.C(n_201),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_197),
.B(n_199),
.C(n_200),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_283),
.B(n_288),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_269),
.B(n_282),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_247),
.B(n_268),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_227),
.B(n_246),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_207),
.B(n_217),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_224),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_222),
.C(n_224),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_223),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_225),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_234),
.B(n_245),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_239),
.B(n_244),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_236),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_248),
.B(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_260),
.B1(n_266),
.B2(n_267),
.Y(n_249)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_255),
.B1(n_258),
.B2(n_259),
.Y(n_250)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_255),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_259),
.C(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_257),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_260),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_271),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_278),
.C(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_294),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_294),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_291),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_303),
.B(n_306),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_299),
.B(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_325),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_313),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_323),
.B2(n_324),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);


endmodule