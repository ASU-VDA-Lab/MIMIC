module fake_jpeg_15000_n_142 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_142);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_142;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_5),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_36),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_30),
.Y(n_63)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_SL g34 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_22),
.B(n_18),
.C(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_27),
.B1(n_15),
.B2(n_26),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_33),
.A2(n_25),
.B1(n_21),
.B2(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_15),
.B1(n_27),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_13),
.B1(n_21),
.B2(n_25),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_64),
.B1(n_44),
.B2(n_46),
.Y(n_83)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_2),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_4),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_12),
.B(n_53),
.C(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_20),
.B1(n_16),
.B2(n_22),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_38),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_67),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_49),
.B(n_2),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_80),
.B(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_8),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_8),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_7),
.Y(n_78)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_7),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_52),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_63),
.B1(n_46),
.B2(n_54),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

CKINVDCx10_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_57),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_55),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_63),
.C(n_52),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_99),
.C(n_77),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_84),
.B1(n_68),
.B2(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_48),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_81),
.B(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_99),
.C(n_93),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_73),
.B1(n_83),
.B2(n_79),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_105),
.B1(n_111),
.B2(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_108),
.B(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_92),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_114),
.A2(n_101),
.B1(n_102),
.B2(n_63),
.Y(n_124)
);

A2O1A1O1Ixp25_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_91),
.B(n_87),
.C(n_98),
.D(n_88),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_80),
.C(n_69),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_97),
.C(n_86),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_111),
.A2(n_97),
.B1(n_80),
.B2(n_69),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_120),
.B(n_96),
.C(n_117),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_106),
.A3(n_107),
.B1(n_82),
.B2(n_96),
.C(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_124),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_125),
.B(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_127),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_131),
.C(n_132),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_113),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_116),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_125),
.B(n_121),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_131),
.B(n_48),
.Y(n_138)
);

OAI321xp33_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_100),
.A3(n_62),
.B1(n_48),
.B2(n_68),
.C(n_57),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_136),
.B(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_89),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_137),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_134),
.B(n_45),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_45),
.B1(n_57),
.B2(n_139),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_45),
.Y(n_142)
);


endmodule