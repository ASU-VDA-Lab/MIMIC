module fake_jpeg_14851_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_6),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_17),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_21),
.A2(n_19),
.B1(n_17),
.B2(n_14),
.Y(n_39)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_27),
.Y(n_35)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_20),
.A2(n_16),
.B1(n_13),
.B2(n_19),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_41),
.B1(n_11),
.B2(n_10),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_10),
.C(n_11),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_26),
.B(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_23),
.A2(n_13),
.B1(n_16),
.B2(n_22),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_7),
.B1(n_8),
.B2(n_49),
.Y(n_55)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx12f_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_3),
.B(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_43),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.C(n_36),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_31),
.A2(n_35),
.B(n_37),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_55),
.B1(n_56),
.B2(n_50),
.Y(n_58)
);

XOR2x2_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_34),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.C(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_43),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_42),
.B(n_45),
.Y(n_61)
);

AOI31xp33_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_57),
.A3(n_54),
.B(n_51),
.Y(n_64)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_65),
.B(n_60),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_68),
.B(n_65),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_59),
.B(n_55),
.Y(n_68)
);


endmodule