module fake_jpeg_8580_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_44),
.Y(n_59)
);

INVx5_ASAP7_75t_SL g72 ( 
.A(n_59),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_62),
.Y(n_70)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_65),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_0),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx6f_ASAP7_75t_SL g67 ( 
.A(n_50),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_78),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_41),
.B1(n_54),
.B2(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_56),
.B1(n_57),
.B2(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_56),
.B1(n_55),
.B2(n_53),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_47),
.B1(n_51),
.B2(n_50),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_22),
.B1(n_38),
.B2(n_35),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_80),
.B1(n_83),
.B2(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_5),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_86),
.B(n_6),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_87)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_89),
.B(n_92),
.Y(n_99)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_8),
.Y(n_94)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_99),
.A2(n_90),
.B1(n_95),
.B2(n_71),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_98),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_94),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_107),
.A2(n_95),
.B1(n_91),
.B2(n_76),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_109),
.B(n_70),
.CI(n_11),
.CON(n_110),
.SN(n_110)
);

AOI322xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_10),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C1(n_16),
.C2(n_20),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_110),
.B(n_25),
.C(n_26),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_32),
.Y(n_114)
);


endmodule