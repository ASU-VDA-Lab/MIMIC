module fake_jpeg_22471_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_36),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

CKINVDCx9p33_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_1),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_31),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_21),
.Y(n_50)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_46),
.B1(n_21),
.B2(n_16),
.Y(n_51)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_22),
.B1(n_30),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_47),
.A2(n_57),
.B1(n_58),
.B2(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_48),
.B(n_66),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_52),
.Y(n_80)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_55),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_60),
.Y(n_87)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_20),
.B1(n_22),
.B2(n_30),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_20),
.B1(n_16),
.B2(n_46),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp67_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_15),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_24),
.Y(n_67)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OR2x2_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_40),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_26),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_45),
.A2(n_23),
.B1(n_25),
.B2(n_17),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_25),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_52),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_97),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_23),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_100),
.Y(n_117)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_26),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_56),
.B1(n_64),
.B2(n_74),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_27),
.B(n_86),
.C(n_79),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_106),
.Y(n_131)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_18),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_58),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_112),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_99),
.A2(n_78),
.B1(n_83),
.B2(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_121),
.B1(n_92),
.B2(n_96),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_72),
.C(n_51),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_9),
.Y(n_119)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_27),
.B1(n_3),
.B2(n_2),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_27),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_121),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_125),
.B(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_87),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_128),
.A2(n_140),
.B1(n_112),
.B2(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_95),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_80),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_27),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_3),
.Y(n_141)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_146),
.B(n_148),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_147),
.Y(n_161)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_110),
.B1(n_114),
.B2(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_131),
.B(n_129),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_143),
.B(n_111),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_157),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_3),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_135),
.Y(n_165)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_170),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_139),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_171),
.B(n_174),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_139),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_176),
.C(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_147),
.B1(n_145),
.B2(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_178),
.B(n_180),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_173),
.B(n_160),
.Y(n_180)
);

NAND2x1_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_175),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_179),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_167),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_177),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_185),
.B(n_186),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_142),
.C(n_128),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_128),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_8),
.Y(n_190)
);


endmodule