module fake_jpeg_18309_n_299 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_299);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx6_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_19),
.B1(n_16),
.B2(n_13),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_42),
.B1(n_45),
.B2(n_51),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_19),
.B1(n_13),
.B2(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_19),
.B1(n_13),
.B2(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_26),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_19),
.B1(n_16),
.B2(n_26),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_33),
.B1(n_35),
.B2(n_17),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_58),
.B1(n_72),
.B2(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_62),
.Y(n_82)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_39),
.B1(n_46),
.B2(n_35),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_28),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_70),
.C(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_32),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_63),
.B(n_64),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_66),
.Y(n_98)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_15),
.B1(n_28),
.B2(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_22),
.B1(n_18),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_20),
.B1(n_18),
.B2(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_30),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_17),
.B1(n_20),
.B2(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_78),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_14),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_52),
.C(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_21),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_15),
.B1(n_14),
.B2(n_27),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_90),
.B(n_95),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_63),
.B1(n_60),
.B2(n_68),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_29),
.B(n_15),
.C(n_25),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_27),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_89),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_56),
.B(n_59),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_62),
.A2(n_23),
.B1(n_25),
.B2(n_24),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_63),
.B1(n_64),
.B2(n_70),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_60),
.B1(n_68),
.B2(n_59),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_99),
.A2(n_101),
.B1(n_110),
.B2(n_115),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_102),
.B(n_106),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_108),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_61),
.C(n_70),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_83),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_94),
.C(n_91),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_118),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_58),
.B1(n_73),
.B2(n_55),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_57),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_87),
.B1(n_90),
.B2(n_98),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_54),
.B(n_57),
.Y(n_138)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_81),
.B1(n_93),
.B2(n_84),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_98),
.B1(n_55),
.B2(n_74),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_97),
.B1(n_78),
.B2(n_96),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_125),
.A2(n_132),
.B1(n_137),
.B2(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_140),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_104),
.B(n_107),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_130),
.B(n_0),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_74),
.B1(n_77),
.B2(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_6),
.B1(n_11),
.B2(n_2),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_77),
.B1(n_88),
.B2(n_54),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_147),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_67),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_134),
.B(n_142),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_120),
.B1(n_117),
.B2(n_116),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_143),
.B(n_153),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_27),
.B1(n_14),
.B2(n_23),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_103),
.C(n_106),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_25),
.B(n_24),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_57),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_103),
.B(n_25),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_1),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_154),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_67),
.B1(n_23),
.B2(n_24),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_117),
.A2(n_111),
.B(n_123),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_24),
.C(n_23),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_118),
.C(n_114),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_156),
.B(n_160),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_122),
.Y(n_158)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_135),
.B(n_100),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_179),
.C(n_186),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_100),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_126),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_166),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_167),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_172),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_178),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_6),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_128),
.A2(n_147),
.B1(n_153),
.B2(n_140),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_0),
.C(n_1),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_7),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_185),
.B1(n_150),
.B2(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_138),
.B(n_148),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_182),
.A2(n_183),
.B1(n_131),
.B2(n_153),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_125),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_7),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_143),
.Y(n_195)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_127),
.B(n_0),
.C(n_1),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_189),
.A2(n_175),
.B1(n_163),
.B2(n_170),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_203),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_168),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_168),
.B1(n_150),
.B2(n_171),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_137),
.Y(n_201)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_130),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_129),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_206),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_132),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_128),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_205),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_155),
.C(n_141),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_179),
.C(n_186),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_212),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_178),
.B1(n_163),
.B2(n_181),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_228),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_170),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_219),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_201),
.A2(n_169),
.B1(n_161),
.B2(n_174),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_204),
.B1(n_199),
.B2(n_182),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_193),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_161),
.B(n_173),
.C(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_195),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_173),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_174),
.B1(n_171),
.B2(n_183),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

INVx13_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_209),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_235),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_226),
.B(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_224),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_207),
.B(n_197),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_243),
.A2(n_236),
.B1(n_197),
.B2(n_233),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_228),
.B1(n_196),
.B2(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_247),
.C(n_225),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_250),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_241),
.C(n_238),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_252),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_258),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_213),
.C(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_190),
.C(n_221),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_237),
.A2(n_196),
.B1(n_200),
.B2(n_214),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_190),
.C(n_194),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_2),
.C(n_3),
.Y(n_268)
);

OAI321xp33_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_210),
.A3(n_240),
.B1(n_234),
.B2(n_194),
.C(n_232),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_267),
.B(n_5),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_256),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_246),
.B(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_4),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_3),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_271),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_257),
.Y(n_272)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_279),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_268),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_278),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_270),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_265),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_9),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_275),
.B(n_8),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_281),
.A2(n_284),
.B(n_9),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_9),
.B(n_10),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_10),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_287),
.B(n_276),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_291),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_285),
.A2(n_9),
.B(n_10),
.Y(n_290)
);

NAND3xp33_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_292),
.C(n_283),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_281),
.B(n_286),
.Y(n_295)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_293),
.C(n_282),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_296),
.A2(n_10),
.B(n_11),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_11),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_12),
.Y(n_299)
);


endmodule