module fake_jpeg_20342_n_407 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_407);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_407;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_2),
.B(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_44),
.B(n_47),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_46),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_48),
.B(n_71),
.Y(n_103)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_52),
.Y(n_128)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_54),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_62),
.B(n_63),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_65),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_68),
.B(n_69),
.Y(n_125)
);

INVx6_ASAP7_75t_SL g69 ( 
.A(n_16),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_70),
.B(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_17),
.B(n_12),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_32),
.B(n_13),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_75),
.B(n_85),
.Y(n_130)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_82),
.Y(n_123)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_27),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_30),
.B1(n_15),
.B2(n_40),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_88),
.A2(n_95),
.B1(n_99),
.B2(n_102),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_49),
.A2(n_31),
.B1(n_30),
.B2(n_15),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_90),
.A2(n_93),
.B1(n_105),
.B2(n_109),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_50),
.A2(n_30),
.B1(n_15),
.B2(n_31),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_40),
.B1(n_32),
.B2(n_42),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_27),
.C(n_37),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_104),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_20),
.B1(n_41),
.B2(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_100),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_42),
.B1(n_41),
.B2(n_36),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_38),
.B1(n_26),
.B2(n_28),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_86),
.A2(n_33),
.B1(n_28),
.B2(n_22),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_67),
.A2(n_33),
.B1(n_22),
.B2(n_20),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_119),
.B1(n_132),
.B2(n_137),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_68),
.A2(n_18),
.B1(n_26),
.B2(n_12),
.Y(n_119)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_18),
.B1(n_27),
.B2(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_0),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_135),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_69),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_58),
.A2(n_2),
.B1(n_3),
.B2(n_6),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_74),
.A2(n_2),
.B1(n_3),
.B2(n_7),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_138),
.A2(n_121),
.B1(n_108),
.B2(n_111),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_140),
.Y(n_187)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_147),
.B(n_151),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_54),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_59),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_149),
.B(n_158),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_110),
.B(n_60),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_157),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_103),
.B(n_8),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_8),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_152),
.B(n_166),
.Y(n_207)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_104),
.B(n_51),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_155),
.B(n_163),
.C(n_97),
.Y(n_201)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_72),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_96),
.B(n_66),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_164),
.Y(n_216)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_183),
.B1(n_92),
.B2(n_134),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_51),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_87),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_107),
.B(n_8),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_45),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_171),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_109),
.B(n_79),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_180),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_170),
.A2(n_89),
.B1(n_94),
.B2(n_101),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_8),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_172),
.Y(n_206)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_111),
.A2(n_78),
.B1(n_52),
.B2(n_11),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_126),
.A2(n_9),
.B(n_10),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_125),
.B(n_10),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_122),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_91),
.Y(n_179)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_10),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_108),
.A2(n_11),
.B1(n_121),
.B2(n_128),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_112),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_128),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_112),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_185),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_97),
.B(n_11),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_188),
.B(n_195),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_89),
.B1(n_101),
.B2(n_94),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_194),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_134),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_196),
.A2(n_201),
.B1(n_156),
.B2(n_157),
.Y(n_255)
);

AO21x2_ASAP7_75t_L g202 ( 
.A1(n_146),
.A2(n_140),
.B(n_158),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_202),
.A2(n_224),
.B1(n_173),
.B2(n_161),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_182),
.B1(n_169),
.B2(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_127),
.B1(n_122),
.B2(n_131),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_115),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_153),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_143),
.B(n_139),
.C(n_106),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_155),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_182),
.A2(n_180),
.B1(n_144),
.B2(n_168),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_163),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_106),
.B(n_127),
.C(n_124),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_144),
.A2(n_139),
.B1(n_145),
.B2(n_143),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_155),
.A2(n_163),
.B1(n_141),
.B2(n_142),
.Y(n_224)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_220),
.Y(n_229)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_222),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_231),
.B(n_233),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_147),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_160),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_171),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_243),
.Y(n_265)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_240),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_212),
.C(n_201),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_184),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_200),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_242),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_151),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_200),
.B(n_189),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_246),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_219),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_245),
.B(n_249),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_193),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_248),
.A2(n_226),
.B1(n_202),
.B2(n_209),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_190),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_250),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_197),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_251),
.A2(n_254),
.B(n_257),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_204),
.B1(n_192),
.B2(n_221),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_166),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_197),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_199),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_256),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_258),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_225),
.B(n_152),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_259),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_205),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_198),
.B(n_202),
.Y(n_290)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_261),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_267),
.A2(n_276),
.B1(n_285),
.B2(n_248),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_275),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_288),
.C(n_289),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_229),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_226),
.B1(n_202),
.B2(n_209),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_279),
.B1(n_231),
.B2(n_233),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_228),
.A2(n_202),
.B1(n_211),
.B2(n_198),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_281),
.A2(n_188),
.B(n_234),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_228),
.A2(n_202),
.B1(n_218),
.B2(n_196),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_238),
.B(n_196),
.C(n_195),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_244),
.B(n_195),
.C(n_225),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_290),
.A2(n_227),
.B(n_257),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_267),
.A2(n_236),
.B1(n_230),
.B2(n_258),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_303),
.B1(n_312),
.B2(n_314),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_293),
.B(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_269),
.B(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_296),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_269),
.B(n_243),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_300),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_255),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_299),
.B(n_315),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_280),
.Y(n_301)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_301),
.Y(n_338)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_304),
.Y(n_334)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_305),
.A2(n_311),
.B1(n_316),
.B2(n_317),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_251),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_306),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_278),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_254),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_246),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_262),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_279),
.A2(n_227),
.B1(n_239),
.B2(n_256),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_262),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_239),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_276),
.A2(n_250),
.B1(n_188),
.B2(n_219),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_321),
.B(n_308),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_303),
.A2(n_282),
.B1(n_284),
.B2(n_290),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_323),
.A2(n_326),
.B1(n_339),
.B2(n_297),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_299),
.C(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_328),
.C(n_336),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_293),
.A2(n_284),
.B1(n_285),
.B2(n_268),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_289),
.C(n_281),
.Y(n_328)
);

XOR2x2_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_281),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_329),
.A2(n_310),
.B1(n_302),
.B2(n_296),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_305),
.B(n_265),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_333),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_268),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_265),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_337),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_301),
.B(n_264),
.C(n_286),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_271),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_300),
.A2(n_275),
.B1(n_286),
.B2(n_283),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_340),
.B(n_333),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_320),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_341),
.B(n_344),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_321),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_322),
.B(n_291),
.Y(n_344)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_294),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_347),
.B(n_355),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_295),
.Y(n_348)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_348),
.Y(n_366)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_334),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_349),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_350),
.B(n_351),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_335),
.B(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_338),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_352),
.A2(n_357),
.B1(n_339),
.B2(n_318),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_328),
.B(n_206),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_353),
.A2(n_331),
.B1(n_330),
.B2(n_323),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_306),
.C(n_304),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_332),
.C(n_327),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_283),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_329),
.A2(n_277),
.B(n_264),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_371),
.C(n_346),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_360),
.B(n_368),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_363),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_319),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_367),
.B(n_370),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_324),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_346),
.B(n_207),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_354),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_372),
.A2(n_374),
.B(n_207),
.Y(n_389)
);

OA21x2_ASAP7_75t_SL g374 ( 
.A1(n_364),
.A2(n_340),
.B(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_369),
.B(n_370),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_376),
.B(n_378),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_365),
.A2(n_342),
.B1(n_352),
.B2(n_357),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_380),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_367),
.B(n_356),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_261),
.C(n_215),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_242),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_382),
.B(n_362),
.Y(n_386)
);

NOR2x1_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_363),
.Y(n_383)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_373),
.A2(n_359),
.B1(n_361),
.B2(n_371),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_386),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_241),
.C(n_240),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_387),
.B(n_375),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_389),
.A2(n_390),
.B(n_381),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_241),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_391),
.A2(n_375),
.B(n_377),
.Y(n_394)
);

AOI322xp5_ASAP7_75t_L g398 ( 
.A1(n_394),
.A2(n_395),
.A3(n_385),
.B1(n_383),
.B2(n_387),
.C1(n_384),
.C2(n_388),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_397),
.C(n_179),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_390),
.A2(n_261),
.B(n_263),
.Y(n_397)
);

AO221x1_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_400),
.B1(n_274),
.B2(n_210),
.C(n_181),
.Y(n_403)
);

FAx1_ASAP7_75t_SL g399 ( 
.A(n_393),
.B(n_312),
.CI(n_263),
.CON(n_399),
.SN(n_399)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_399),
.B(n_401),
.Y(n_402)
);

AOI322xp5_ASAP7_75t_L g400 ( 
.A1(n_392),
.A2(n_274),
.A3(n_177),
.B1(n_247),
.B2(n_237),
.C1(n_210),
.C2(n_162),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_403),
.A2(n_179),
.B(n_154),
.Y(n_405)
);

AOI321xp33_ASAP7_75t_L g404 ( 
.A1(n_402),
.A2(n_399),
.A3(n_274),
.B1(n_154),
.B2(n_181),
.C(n_165),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_405),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_179),
.Y(n_407)
);


endmodule