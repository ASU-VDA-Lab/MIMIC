module real_jpeg_31850_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_572;
wire n_405;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g102 ( 
.A(n_0),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_0),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_0),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_0),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_1),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_1),
.B(n_65),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g203 ( 
.A(n_1),
.B(n_144),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_1),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g344 ( 
.A(n_1),
.B(n_258),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_1),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_1),
.B(n_389),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_2),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_3),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_3),
.B(n_319),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_3),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_3),
.B(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_3),
.B(n_339),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_3),
.B(n_477),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_3),
.B(n_389),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_4),
.A2(n_21),
.B(n_24),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_5),
.B(n_229),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_5),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_5),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_5),
.B(n_400),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_5),
.B(n_75),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_5),
.B(n_480),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_6),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_6),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_6),
.B(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_6),
.B(n_331),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_7),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_9),
.Y(n_529)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_10),
.Y(n_259)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_10),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_L g245 ( 
.A(n_11),
.B(n_246),
.Y(n_245)
);

NAND2x1_ASAP7_75t_L g323 ( 
.A(n_11),
.B(n_99),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_11),
.B(n_351),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_11),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_11),
.B(n_492),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g527 ( 
.A(n_11),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_11),
.B(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_12),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_12),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_12),
.B(n_65),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_12),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_12),
.B(n_208),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_12),
.B(n_541),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_12),
.B(n_549),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_25),
.Y(n_24)
);

NAND2x1_ASAP7_75t_SL g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_14),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_14),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_14),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_14),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_14),
.B(n_101),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_14),
.B(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_15),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g74 ( 
.A(n_16),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_16),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_16),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_16),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_16),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_16),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_17),
.Y(n_135)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_18),
.B(n_192),
.Y(n_191)
);

NAND2x1_ASAP7_75t_L g231 ( 
.A(n_18),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_18),
.B(n_261),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_18),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_18),
.B(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_18),
.B(n_497),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_18),
.B(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_18),
.B(n_524),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_19),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_19),
.B(n_187),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_19),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_19),
.B(n_389),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

O2A1O1Ixp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_301),
.B(n_576),
.C(n_590),
.Y(n_25)
);

OAI211xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_177),
.B(n_285),
.C(n_286),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g573 ( 
.A(n_27),
.B(n_574),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_148),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_28),
.B(n_148),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_110),
.C(n_125),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_29),
.B(n_283),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_78),
.B(n_109),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_30),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_49),
.C(n_62),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_31),
.B(n_49),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_32),
.B(n_38),
.C(n_42),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_36),
.Y(n_173)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_36),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_36),
.Y(n_233)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_36),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_46),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_47),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.C(n_56),
.Y(n_49)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_50),
.B(n_53),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_52),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_55),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_56),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_58),
.B(n_326),
.Y(n_473)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g535 ( 
.A(n_60),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_61),
.Y(n_348)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_62),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_63),
.B(n_69),
.C(n_77),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_67),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_77),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_69),
.A2(n_70),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_69),
.B(n_113),
.C(n_117),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_98),
.C(n_100),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_74),
.A2(n_77),
.B1(n_100),
.B2(n_190),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_76),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_76),
.Y(n_477)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_76),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_96),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_96),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_79),
.A2(n_80),
.B1(n_96),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2x1_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_92),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_86),
.B1(n_87),
.B2(n_91),
.Y(n_81)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_85),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_91),
.C(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_89),
.Y(n_458)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_90),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_94),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_95),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_96),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.C(n_108),
.Y(n_96)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_97),
.Y(n_199)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_99),
.Y(n_299)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_100),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_100),
.A2(n_186),
.B1(n_190),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_103),
.B(n_108),
.Y(n_200)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_105),
.Y(n_294)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_105),
.Y(n_343)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_108),
.B(n_202),
.C(n_210),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_108),
.B(n_211),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_110),
.B(n_125),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_123),
.C(n_124),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_111),
.B(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_113),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_116),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_159),
.C(n_160),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_115),
.Y(n_209)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_115),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_123),
.B(n_124),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_147),
.C(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_132),
.C(n_136),
.Y(n_150)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_146),
.B2(n_147),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_175),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_150),
.B(n_151),
.C(n_175),
.Y(n_287)
);

XNOR2x1_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_161),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_153),
.B(n_158),
.C(n_161),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_159),
.B(n_164),
.C(n_170),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_170),
.B1(n_171),
.B2(n_174),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_163),
.A2(n_164),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_163),
.B(n_292),
.C(n_297),
.Y(n_586)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_279),
.B(n_284),
.Y(n_177)
);

NOR2xp67_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_268),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_179),
.B(n_268),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_R g179 ( 
.A(n_180),
.B(n_216),
.C(n_219),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_180),
.A2(n_181),
.B1(n_216),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_197),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.C(n_194),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_183),
.B(n_185),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.C(n_191),
.Y(n_185)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_189),
.Y(n_386)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_194),
.B(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_198),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_SL g269 ( 
.A(n_201),
.B(n_270),
.C(n_272),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_202),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.C(n_207),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_204),
.Y(n_242)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_215),
.Y(n_584)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_216),
.Y(n_363)
);

XNOR2x2_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_220),
.B(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_243),
.C(n_265),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.C(n_241),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_222),
.B(n_226),
.C(n_241),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_226),
.Y(n_374)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_239),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_231),
.B(n_240),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_234),
.Y(n_404)
);

INVx3_ASAP7_75t_SL g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_241),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_243),
.B(n_266),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_254),
.B(n_264),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.C(n_252),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_245),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_SL g356 ( 
.A(n_245),
.B(n_249),
.C(n_252),
.Y(n_356)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_249),
.A2(n_252),
.B1(n_253),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_260),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_255),
.B(n_260),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_255),
.B(n_260),
.Y(n_357)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_259),
.Y(n_402)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_259),
.Y(n_498)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_274),
.C(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_279),
.B(n_575),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_282),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_287),
.B(n_288),
.Y(n_589)
);

BUFx24_ASAP7_75t_SL g593 ( 
.A(n_288),
.Y(n_593)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.CI(n_291),
.CON(n_288),
.SN(n_288)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_296),
.A2(n_297),
.B1(n_580),
.B2(n_581),
.Y(n_579)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_300),
.B(n_582),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_573),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_412),
.B(n_570),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_364),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g570 ( 
.A1(n_304),
.A2(n_571),
.B(n_572),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_361),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_L g572 ( 
.A(n_305),
.B(n_361),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_310),
.C(n_359),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_307),
.B(n_359),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_310),
.B(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_334),
.C(n_352),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_368),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.C(n_328),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_313),
.B(n_315),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_316),
.A2(n_317),
.B1(n_328),
.B2(n_329),
.Y(n_439)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_321),
.B(n_324),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_379),
.Y(n_378)
);

AOI21xp33_ASAP7_75t_SL g324 ( 
.A1(n_319),
.A2(n_325),
.B(n_327),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_322),
.B1(n_327),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_327),
.Y(n_380)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

OA21x2_ASAP7_75t_SL g423 ( 
.A1(n_329),
.A2(n_330),
.B(n_333),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_333),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_353),
.B1(n_354),
.B2(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_345),
.C(n_349),
.Y(n_335)
);

XOR2x1_ASAP7_75t_L g408 ( 
.A(n_336),
.B(n_409),
.Y(n_408)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_342),
.C(n_344),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_337),
.A2(n_338),
.B1(n_344),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_340),
.Y(n_494)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_345),
.A2(n_346),
.B1(n_349),
.B2(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_358),
.Y(n_354)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_356),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_410),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_365),
.B(n_410),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.C(n_375),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_367),
.B(n_371),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_375),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_403),
.C(n_406),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_376),
.A2(n_377),
.B1(n_416),
.B2(n_417),
.Y(n_415)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.C(n_392),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_378),
.B(n_462),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_381),
.A2(n_392),
.B1(n_393),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_381),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_387),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_382),
.A2(n_383),
.B1(n_387),
.B2(n_388),
.Y(n_459)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_391),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_391),
.Y(n_551)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_398),
.C(n_399),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_394),
.A2(n_395),
.B1(n_399),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_398),
.B(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_402),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_403),
.A2(n_407),
.B1(n_408),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_403),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_466),
.B(n_568),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_440),
.B(n_443),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_414),
.B(n_440),
.C(n_569),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_419),
.C(n_436),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_419),
.B(n_437),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_423),
.C(n_424),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_423),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_424),
.B(n_446),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_430),
.C(n_432),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_425),
.B(n_482),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_426),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.Y(n_472)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_430),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_482)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_464),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_444),
.B(n_464),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.C(n_460),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_484),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_451),
.C(n_459),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_459),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.C(n_456),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_452),
.B(n_456),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_453),
.B(n_517),
.Y(n_516)
);

INVx3_ASAP7_75t_SL g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_458),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_485),
.B(n_567),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_483),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_SL g567 ( 
.A(n_468),
.B(n_483),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.C(n_481),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g564 ( 
.A(n_469),
.B(n_565),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_471),
.B(n_481),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.C(n_474),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_472),
.B(n_473),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_511),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

AO22x1_ASAP7_75t_L g507 ( 
.A1(n_475),
.A2(n_476),
.B1(n_478),
.B2(n_479),
.Y(n_507)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_562),
.B(n_566),
.Y(n_485)
);

OAI21x1_ASAP7_75t_SL g486 ( 
.A1(n_487),
.A2(n_519),
.B(n_561),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_508),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_488),
.B(n_508),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_501),
.C(n_507),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_489),
.A2(n_490),
.B1(n_557),
.B2(n_559),
.Y(n_556)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_495),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_514),
.C(n_515),
.Y(n_513)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_499),
.Y(n_495)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_496),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_501),
.A2(n_502),
.B1(n_507),
.B2(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_506),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_506),
.Y(n_537)
);

INVx4_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_507),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_510),
.B1(n_512),
.B2(n_518),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_509),
.B(n_513),
.C(n_516),
.Y(n_563)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_554),
.B(n_560),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_521),
.A2(n_538),
.B(n_553),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_530),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_522),
.B(n_530),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_523),
.B(n_527),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_523),
.B(n_527),
.Y(n_546)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx8_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_527),
.B(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_537),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_532),
.A2(n_533),
.B1(n_534),
.B2(n_536),
.Y(n_531)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_532),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_536),
.C(n_537),
.Y(n_555)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_539),
.A2(n_547),
.B(n_552),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_546),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_546),
.Y(n_552)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx3_ASAP7_75t_SL g549 ( 
.A(n_550),
.Y(n_549)
);

INVx8_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_556),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_555),
.B(n_556),
.Y(n_560)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_557),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_564),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_577),
.B(n_588),
.Y(n_576)
);

AOI221xp5_ASAP7_75t_L g577 ( 
.A1(n_578),
.A2(n_579),
.B1(n_585),
.B2(n_586),
.C(n_587),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_578),
.A2(n_579),
.B1(n_585),
.B2(n_586),
.Y(n_592)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_579),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_581),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_581),
.B(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_586),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_587),
.B(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);


endmodule