module fake_jpeg_2522_n_65 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_65);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_65;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_4),
.B(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_24),
.B(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_45),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_26),
.B1(n_22),
.B2(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_41),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.C(n_52),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_37),
.B(n_36),
.Y(n_49)
);

OAI31xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_51),
.A3(n_26),
.B(n_3),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_8),
.C(n_17),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_7),
.C(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_2),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_2),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_11),
.C(n_13),
.Y(n_60)
);

AOI31xp67_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.A3(n_5),
.B(n_6),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_59),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_64),
.Y(n_65)
);


endmodule