module real_jpeg_5715_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_2),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_2),
.B(n_51),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_3),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_3),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_3),
.B(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

NAND2x1p5_ASAP7_75t_L g39 ( 
.A(n_5),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_5),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_83),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_5),
.B(n_98),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_5),
.B(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_7),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_7),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_7),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_7),
.B(n_177),
.Y(n_176)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_8),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_8),
.Y(n_211)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_8),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_8),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_9),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_9),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_9),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_9),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_9),
.B(n_108),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_9),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_10),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_10),
.B(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_11),
.Y(n_183)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_13),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_13),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_13),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_14),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_14),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_14),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_14),
.B(n_37),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_14),
.B(n_245),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_14),
.B(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_15),
.Y(n_157)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_17),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_17),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_17),
.B(n_238),
.Y(n_237)
);

XNOR2x2_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_193),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_192),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_165),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_22),
.B(n_165),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_99),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_69),
.C(n_80),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_24),
.B(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_43),
.C(n_54),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_25),
.A2(n_26),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

MAJx2_ASAP7_75t_L g150 ( 
.A(n_27),
.B(n_35),
.C(n_42),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_28),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_32),
.Y(n_271)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_44),
.B(n_55),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_45),
.B(n_50),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_48),
.Y(n_142)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_48),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.C(n_65),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_56),
.B(n_65),
.Y(n_283)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_60),
.B(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_62),
.Y(n_266)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_63),
.Y(n_229)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_67),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_69),
.B(n_80),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_74),
.C(n_76),
.Y(n_115)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_89),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_82),
.B(n_84),
.C(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_89),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.C(n_96),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_90),
.B(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_93),
.A2(n_96),
.B1(n_97),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_93),
.Y(n_188)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_131),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_113),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_130),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_151),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_143),
.C(n_150),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_134),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_139),
.C(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_142),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_144),
.B(n_147),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_150),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx6_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_154),
.B1(n_163),
.B2(n_164),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_160),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_189),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_167),
.B(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_169),
.B(n_189),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.C(n_185),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_170),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.C(n_181),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_171),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_259)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_179),
.B(n_182),
.Y(n_279)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_190),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_304),
.B(n_308),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_291),
.B(n_303),
.Y(n_194)
);

AOI21x1_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_275),
.B(n_290),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_249),
.B(n_274),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_231),
.B(n_248),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_213),
.B(n_230),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_209),
.B(n_212),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_207),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_204),
.Y(n_214)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_215),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_222),
.B2(n_223),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_225),
.C(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_219),
.Y(n_239)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_247),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_239),
.C(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_237),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_240),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_262),
.C(n_263),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_244),
.Y(n_263)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_246),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_252),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_261),
.C(n_264),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_256),
.C(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_270),
.C(n_272),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_270),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_289),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_289),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_280),
.C(n_302),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_286),
.C(n_287),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_301),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_295),
.C(n_298),
.Y(n_307)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);


endmodule