module fake_jpeg_24343_n_344 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.C(n_1),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_19),
.B(n_20),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_58),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_19),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_30),
.B(n_20),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_34),
.B(n_35),
.C(n_31),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_69),
.Y(n_72)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_43),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_21),
.B1(n_22),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_21),
.B1(n_22),
.B2(n_34),
.Y(n_78)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_22),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_26),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_87),
.Y(n_110)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_77),
.A2(n_81),
.B1(n_89),
.B2(n_93),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_53),
.B(n_26),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_84),
.Y(n_106)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_91),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_39),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_85),
.A2(n_97),
.B(n_32),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_48),
.B1(n_21),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_43),
.B1(n_64),
.B2(n_63),
.Y(n_102)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_95),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_17),
.B1(n_18),
.B2(n_32),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_0),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_99),
.Y(n_123)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_98),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g97 ( 
.A(n_52),
.B(n_43),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_100),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_113),
.B1(n_119),
.B2(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_103),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_105),
.A2(n_107),
.B(n_128),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_41),
.B(n_40),
.C(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_112),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_63),
.B1(n_59),
.B2(n_17),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_62),
.C(n_70),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_127),
.C(n_90),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_25),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_76),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_80),
.A2(n_17),
.B1(n_18),
.B2(n_49),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_122),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_85),
.A2(n_49),
.B1(n_46),
.B2(n_44),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_100),
.B1(n_95),
.B2(n_91),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_37),
.C(n_41),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_86),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_129),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_92),
.B(n_37),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_133),
.B(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_144),
.B(n_117),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_74),
.C(n_84),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_160),
.C(n_111),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_84),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_146),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_85),
.B1(n_75),
.B2(n_101),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_145),
.Y(n_182)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_149),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_75),
.B1(n_77),
.B2(n_97),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_115),
.B1(n_126),
.B2(n_104),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_97),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_77),
.B1(n_81),
.B2(n_89),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_79),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_117),
.B1(n_111),
.B2(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_154),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g151 ( 
.A(n_108),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_159),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_99),
.B1(n_82),
.B2(n_96),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_123),
.B1(n_119),
.B2(n_113),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_87),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_46),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_110),
.B(n_37),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_161),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_40),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_SL g212 ( 
.A(n_164),
.B(n_178),
.C(n_180),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_176),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_109),
.B(n_131),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_184),
.B(n_185),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_172),
.B1(n_174),
.B2(n_192),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

CKINVDCx10_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_142),
.A2(n_105),
.B1(n_102),
.B2(n_107),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_181),
.C(n_161),
.Y(n_207)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_105),
.B1(n_107),
.B2(n_117),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_157),
.B1(n_139),
.B2(n_136),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_138),
.B(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_8),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_37),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

NOR2x1_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_37),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_141),
.A2(n_114),
.B(n_28),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_193),
.B(n_156),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_140),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_149),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_112),
.Y(n_190)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_190),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_191),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_142),
.A2(n_40),
.B1(n_28),
.B2(n_32),
.Y(n_192)
);

AOI21x1_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_35),
.B(n_1),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_181),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_202),
.C(n_204),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_182),
.A2(n_137),
.B1(n_152),
.B2(n_160),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_203),
.B1(n_210),
.B2(n_168),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_135),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_143),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_169),
.Y(n_228)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_211),
.C(n_220),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_148),
.B1(n_140),
.B2(n_154),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_134),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_145),
.B(n_158),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

OA21x2_ASAP7_75t_SL g214 ( 
.A1(n_164),
.A2(n_185),
.B(n_178),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_179),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_163),
.A2(n_133),
.B(n_112),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_165),
.B(n_180),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_174),
.B1(n_163),
.B2(n_162),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_217),
.A2(n_219),
.B1(n_170),
.B2(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_162),
.A2(n_112),
.B1(n_108),
.B2(n_33),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_108),
.C(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_188),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_35),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_176),
.C(n_191),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_223),
.B(n_192),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_224),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_231),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_228),
.A2(n_234),
.B(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_240),
.B(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_169),
.Y(n_233)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_249),
.C(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_171),
.Y(n_239)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_171),
.Y(n_243)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_194),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_195),
.B1(n_196),
.B2(n_213),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_248),
.B1(n_226),
.B2(n_240),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_204),
.C(n_198),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_195),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_258),
.C(n_265),
.Y(n_274)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_202),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_263),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_200),
.C(n_196),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_268),
.B1(n_224),
.B2(n_229),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_211),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_205),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_151),
.C(n_36),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_270),
.C(n_228),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_36),
.C(n_29),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_248),
.B1(n_33),
.B2(n_31),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_262),
.B(n_247),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_SL g294 ( 
.A(n_273),
.B(n_286),
.C(n_263),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_264),
.A2(n_229),
.B(n_241),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_285),
.B(n_267),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_279),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_278),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_257),
.B(n_225),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_284),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_230),
.C(n_244),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_288),
.C(n_290),
.Y(n_296)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_9),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_268),
.A2(n_233),
.B(n_245),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_227),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_255),
.B(n_227),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g305 ( 
.A1(n_287),
.A2(n_10),
.B(n_14),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_36),
.C(n_29),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_271),
.A2(n_27),
.B1(n_25),
.B2(n_9),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_289),
.A2(n_272),
.B1(n_256),
.B2(n_261),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_27),
.C(n_25),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_10),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_294),
.B(n_303),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_295),
.B(n_304),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_275),
.A2(n_285),
.B1(n_259),
.B2(n_277),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_301),
.B1(n_290),
.B2(n_288),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_266),
.C(n_269),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_300),
.C(n_274),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_270),
.C(n_253),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_273),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_305),
.A2(n_293),
.B(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_318),
.B1(n_12),
.B2(n_14),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_314),
.C(n_15),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_286),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_282),
.Y(n_310)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_282),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_313),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_10),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_7),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_2),
.Y(n_315)
);

NAND5xp2_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_2),
.C(n_3),
.D(n_4),
.E(n_5),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_7),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_11),
.A3(n_13),
.B1(n_15),
.B2(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_322),
.Y(n_330)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_296),
.B(n_295),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_321),
.B(n_311),
.Y(n_329)
);

INVx11_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_328),
.C(n_316),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_15),
.B1(n_3),
.B2(n_6),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_331),
.B(n_334),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_317),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_333),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_325),
.B(n_6),
.C(n_326),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_6),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_320),
.Y(n_339)
);

O2A1O1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_330),
.A2(n_327),
.B(n_326),
.C(n_322),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_339),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g341 ( 
.A1(n_337),
.A2(n_330),
.B(n_338),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_341),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_342),
.B(n_340),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_328),
.Y(n_344)
);


endmodule