module fake_jpeg_20072_n_274 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_241;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_23),
.B1(n_15),
.B2(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_25),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_16),
.B1(n_14),
.B2(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_49),
.Y(n_61)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_53),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_29),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_27),
.B1(n_25),
.B2(n_23),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_39),
.B1(n_27),
.B2(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_56),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_27),
.B1(n_26),
.B2(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_58),
.B1(n_36),
.B2(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_21),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_58),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_62),
.A2(n_65),
.B1(n_47),
.B2(n_50),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_71),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_21),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_78),
.C(n_54),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_39),
.B1(n_34),
.B2(n_26),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_47),
.B1(n_53),
.B2(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_59),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_34),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_24),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_49),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_57),
.C(n_56),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_64),
.B(n_60),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_85),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_90),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_88),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_72),
.B1(n_47),
.B2(n_83),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_49),
.C(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_92),
.Y(n_102)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_68),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_63),
.B1(n_73),
.B2(n_76),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_75),
.B(n_63),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_77),
.B(n_63),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_110),
.B1(n_79),
.B2(n_90),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_82),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_105),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_107),
.Y(n_147)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_89),
.A3(n_81),
.B1(n_96),
.B2(n_73),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_24),
.C(n_28),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_68),
.B1(n_71),
.B2(n_62),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_80),
.A2(n_67),
.B(n_72),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_118),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

XOR2x1_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_24),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_48),
.B1(n_90),
.B2(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_10),
.Y(n_168)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_83),
.B(n_14),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_141),
.B1(n_144),
.B2(n_70),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_72),
.B1(n_45),
.B2(n_74),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_128),
.Y(n_170)
);

AO22x1_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_45),
.B1(n_74),
.B2(n_39),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_137),
.Y(n_149)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_55),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_138),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_28),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_33),
.B(n_28),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_100),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_146),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_33),
.B(n_22),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_98),
.B(n_32),
.C(n_30),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_98),
.C(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_101),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_33),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_162),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_102),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_133),
.C(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_159),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_99),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_119),
.Y(n_160)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_108),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_10),
.B(n_9),
.Y(n_184)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_169),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_165),
.Y(n_188)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_132),
.B1(n_144),
.B2(n_122),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_126),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_124),
.B(n_147),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_127),
.B1(n_138),
.B2(n_141),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_191),
.B1(n_170),
.B2(n_165),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_186),
.C(n_193),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_161),
.A2(n_157),
.B1(n_156),
.B2(n_162),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_184),
.B(n_151),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_182),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_187),
.B(n_151),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_31),
.C(n_30),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_35),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_189),
.B(n_149),
.Y(n_200)
);

XNOR2x1_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_35),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_169),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_70),
.B1(n_51),
.B2(n_40),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_31),
.C(n_30),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_31),
.C(n_51),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_153),
.C(n_164),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_148),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_208),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_205),
.B(n_70),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_200),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_148),
.B1(n_166),
.B2(n_153),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_202),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_203),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_155),
.B(n_154),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_158),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

XOR2x1_ASAP7_75t_SL g209 ( 
.A(n_184),
.B(n_149),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_SL g217 ( 
.A(n_209),
.B(n_194),
.C(n_175),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_174),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_40),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_192),
.B1(n_191),
.B2(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_214),
.A2(n_223),
.B1(n_215),
.B2(n_216),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_193),
.CI(n_186),
.CON(n_218),
.SN(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_222),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_187),
.B1(n_182),
.B2(n_188),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_224),
.A2(n_202),
.B(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_200),
.B1(n_207),
.B2(n_8),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_198),
.C(n_201),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_228),
.C(n_22),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_198),
.C(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_231),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_220),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_227),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_35),
.B(n_40),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_235),
.Y(n_249)
);

OAI22x1_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_35),
.B1(n_7),
.B2(n_8),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_236),
.B1(n_214),
.B2(n_7),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_6),
.B1(n_8),
.B2(n_7),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_237),
.A2(n_221),
.B1(n_226),
.B2(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_240),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_6),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_243),
.Y(n_257)
);

NOR2xp67_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_17),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_245),
.A2(n_247),
.B(n_248),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_246),
.B(n_17),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_6),
.B(n_8),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_5),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_232),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_251),
.C(n_257),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_231),
.B(n_17),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_253),
.B(n_0),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_22),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_256),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_22),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_247),
.A2(n_4),
.B1(n_6),
.B2(n_5),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_258),
.A2(n_248),
.B1(n_5),
.B2(n_3),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_259),
.B(n_260),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_255),
.A2(n_19),
.A3(n_20),
.B1(n_3),
.B2(n_2),
.C1(n_0),
.C2(n_1),
.Y(n_262)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_262),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_19),
.B1(n_20),
.B2(n_2),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_265),
.B(n_260),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_269),
.B(n_267),
.Y(n_270)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_266),
.A2(n_261),
.A3(n_258),
.B1(n_19),
.B2(n_20),
.C1(n_2),
.C2(n_1),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_20),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_0),
.B1(n_1),
.B2(n_146),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_0),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_0),
.B(n_1),
.Y(n_274)
);


endmodule