module fake_jpeg_7141_n_199 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_199);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_46),
.Y(n_77)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_54),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_24),
.B1(n_30),
.B2(n_23),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_24),
.B1(n_29),
.B2(n_22),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_33),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_53),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_32),
.B1(n_29),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_19),
.B1(n_17),
.B2(n_31),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_25),
.Y(n_73)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_19),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_16),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_83),
.B1(n_50),
.B2(n_4),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_76),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_16),
.Y(n_74)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_31),
.B1(n_4),
.B2(n_5),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_27),
.B1(n_75),
.B2(n_78),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_50),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_44),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_97),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_60),
.C(n_49),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_41),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_100),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_51),
.B1(n_49),
.B2(n_56),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_5),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_6),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_109),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_114),
.C(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_66),
.C(n_74),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_82),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_103),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_84),
.B1(n_88),
.B2(n_75),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_69),
.Y(n_123)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_130),
.C(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_122),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_96),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_104),
.C(n_84),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_135),
.B1(n_110),
.B2(n_75),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_101),
.C(n_97),
.Y(n_133)
);

AO21x2_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_82),
.B(n_78),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_92),
.B(n_82),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_140),
.B(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_111),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_80),
.B(n_38),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_116),
.B(n_115),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_152),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_115),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_153),
.Y(n_156)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_117),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_149),
.C(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_119),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_151),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_117),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_51),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_78),
.B1(n_76),
.B2(n_51),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_49),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_125),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_161),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_135),
.A3(n_132),
.B1(n_131),
.B2(n_138),
.C1(n_136),
.C2(n_126),
.Y(n_158)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_151),
.A3(n_152),
.B1(n_153),
.B2(n_145),
.C1(n_149),
.C2(n_35),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_156),
.C(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_172),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_150),
.Y(n_170)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_156),
.B(n_31),
.Y(n_179)
);

NAND4xp25_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_11),
.C(n_13),
.D(n_8),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_56),
.B1(n_43),
.B2(n_41),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g181 ( 
.A1(n_175),
.A2(n_174),
.B(n_169),
.C(n_38),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_166),
.B1(n_162),
.B2(n_165),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_181),
.B1(n_173),
.B2(n_7),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_172),
.B(n_173),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_43),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_11),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_10),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_10),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_189),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_188),
.B(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_6),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_192),
.A2(n_193),
.B(n_6),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_178),
.C(n_181),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_188),
.B(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_14),
.C(n_7),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_7),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_198),
.Y(n_199)
);


endmodule