module fake_netlist_6_542_n_157 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_157);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_157;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_68;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_29),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_19),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_0),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_1),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_15),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_7),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_7),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_34),
.B(n_8),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_67),
.B(n_55),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_40),
.B(n_47),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_67),
.B(n_66),
.C(n_53),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_33),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_34),
.B(n_49),
.C(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_51),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_44),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_35),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_37),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_50),
.B(n_11),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_9),
.Y(n_84)
);

NAND2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_11),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_12),
.Y(n_86)
);

CKINVDCx8_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_53),
.B(n_55),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_55),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_61),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_78),
.B1(n_74),
.B2(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_93),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_97),
.Y(n_102)
);

CKINVDCx11_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_58),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_90),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_94),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_91),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_101),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_107),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_85),
.B1(n_103),
.B2(n_70),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_109),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_110),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_103),
.B1(n_61),
.B2(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_73),
.Y(n_128)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_83),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_125),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_57),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_64),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_122),
.C(n_68),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_130),
.C(n_131),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_121),
.B1(n_123),
.B2(n_59),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_62),
.B1(n_126),
.B2(n_61),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_137),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_142),
.B(n_136),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_62),
.Y(n_148)
);

NAND2x1p5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_59),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_12),
.Y(n_150)
);

OAI211xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_143),
.B(n_72),
.C(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_148),
.C(n_149),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_146),
.B(n_84),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_153),
.B(n_152),
.Y(n_156)
);

OAI221xp5_ASAP7_75t_R g157 ( 
.A1(n_156),
.A2(n_155),
.B1(n_13),
.B2(n_61),
.C(n_92),
.Y(n_157)
);


endmodule