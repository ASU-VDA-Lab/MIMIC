module fake_jpeg_7201_n_105 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_55),
.Y(n_84)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_73),
.B1(n_47),
.B2(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_4),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_74),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_74),
.A2(n_62),
.B1(n_53),
.B2(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_79),
.B1(n_5),
.B2(n_8),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_56),
.B1(n_54),
.B2(n_58),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_57),
.C(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_84),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_89),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_90),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_87),
.B1(n_83),
.B2(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_22),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_23),
.B(n_24),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_99),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_25),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_31),
.B(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_37),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_39),
.Y(n_105)
);


endmodule