module fake_jpeg_25694_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_149;
wire n_48;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_25),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_49),
.B1(n_67),
.B2(n_18),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_16),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_1),
.C(n_2),
.Y(n_50)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_1),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_54),
.A2(n_61),
.B1(n_38),
.B2(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_32),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_32),
.C(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_40),
.A2(n_24),
.B1(n_31),
.B2(n_30),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_29),
.B1(n_27),
.B2(n_26),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_28),
.C(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_34),
.B(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_27),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_33),
.A2(n_28),
.B1(n_18),
.B2(n_26),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_53),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_42),
.B1(n_33),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_63),
.B1(n_60),
.B2(n_52),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_50),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_42),
.B1(n_35),
.B2(n_43),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_55),
.B1(n_54),
.B2(n_44),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_86),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_89),
.B1(n_68),
.B2(n_65),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_2),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_43),
.A3(n_18),
.B1(n_38),
.B2(n_6),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_2),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_65),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_64),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_95),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_81),
.C(n_78),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_83),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_99),
.B(n_102),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_105),
.B(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_57),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_45),
.B(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_108),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_71),
.Y(n_123)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_112),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_44),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_127),
.C(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_103),
.B1(n_94),
.B2(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_134),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_73),
.B1(n_111),
.B2(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_120),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_111),
.B1(n_133),
.B2(n_125),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_93),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_151),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_117),
.B1(n_126),
.B2(n_95),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_117),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_98),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_117),
.A2(n_101),
.B1(n_100),
.B2(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_98),
.B(n_82),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_154),
.A2(n_124),
.B(n_75),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_158),
.C(n_161),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_115),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_110),
.B1(n_72),
.B2(n_85),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_72),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_75),
.A3(n_51),
.B1(n_76),
.B2(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_119),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_163),
.Y(n_186)
);

AO32x1_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_125),
.A3(n_120),
.B1(n_129),
.B2(n_119),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_131),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_169),
.B(n_176),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_142),
.Y(n_177)
);

AOI221xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_154),
.B1(n_162),
.B2(n_153),
.C(n_146),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_181),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_135),
.B(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_107),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_104),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_155),
.Y(n_188)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_158),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_148),
.C(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_197),
.C(n_202),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_151),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_195),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_206),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_44),
.C(n_76),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_172),
.A2(n_122),
.B1(n_68),
.B2(n_48),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_186),
.B1(n_185),
.B2(n_184),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_172),
.C(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_204),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

OAI322xp33_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_15),
.A3(n_5),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_10),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_216),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_164),
.B1(n_174),
.B2(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_220),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_164),
.C(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_205),
.C(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_185),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_221),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_165),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_222),
.A2(n_192),
.B(n_203),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_193),
.A2(n_180),
.B1(n_184),
.B2(n_171),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_204),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_191),
.C(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_226),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_192),
.C(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

XNOR2x1_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_212),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_195),
.C(n_200),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_208),
.B(n_171),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_236),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_200),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_3),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_237),
.A2(n_218),
.B(n_213),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_215),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_240),
.A2(n_227),
.B(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_214),
.B1(n_211),
.B2(n_220),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_243),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g244 ( 
.A(n_229),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_5),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_223),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_247),
.B1(n_237),
.B2(n_219),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_219),
.B1(n_48),
.B2(n_8),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_253),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_255),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_254),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_240),
.B(n_238),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_48),
.B1(n_11),
.B2(n_12),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_10),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_248),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_11),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_255),
.Y(n_263)
);

NOR4xp25_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.D(n_266),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_12),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

AOI321xp33_ASAP7_75t_L g271 ( 
.A1(n_268),
.A2(n_269),
.A3(n_257),
.B1(n_14),
.B2(n_13),
.C(n_38),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_267),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_271),
.A2(n_270),
.B(n_13),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_14),
.Y(n_273)
);


endmodule