module fake_jpeg_2890_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_55),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_52),
.B1(n_53),
.B2(n_50),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_59),
.B1(n_58),
.B2(n_56),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_77),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_71),
.B1(n_61),
.B2(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_71),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_87),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_3),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_67),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_92),
.B(n_105),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_72),
.B1(n_42),
.B2(n_54),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_95),
.B1(n_92),
.B2(n_105),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_51),
.B1(n_55),
.B2(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_46),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_94),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_51),
.B1(n_43),
.B2(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_97),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_76),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_0),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_104),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_17),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_110),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_113),
.B1(n_118),
.B2(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_93),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_38),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_115),
.B(n_117),
.Y(n_128)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_123),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_97),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_130),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_11),
.B(n_12),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_137),
.B(n_106),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_22),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_135),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_12),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_134),
.B(n_13),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_36),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_24),
.B(n_33),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_109),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_139),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_129),
.B1(n_136),
.B2(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_143),
.C(n_128),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_125),
.C(n_147),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_135),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_150),
.A2(n_151),
.B(n_130),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_142),
.B(n_137),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_153),
.C(n_146),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_133),
.B(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_14),
.Y(n_156)
);

AOI321xp33_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_18),
.C(n_20),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_25),
.B(n_28),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_29),
.B(n_34),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_122),
.Y(n_160)
);


endmodule