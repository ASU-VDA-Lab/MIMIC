module real_aes_2982_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_834, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_833, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_834;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_833;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g232 ( .A(n_0), .B(n_154), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_1), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g147 ( .A(n_2), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_3), .B(n_160), .Y(n_173) );
NAND2xp33_ASAP7_75t_SL g224 ( .A(n_4), .B(n_158), .Y(n_224) );
INVx1_ASAP7_75t_L g205 ( .A(n_5), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_6), .B(n_178), .Y(n_551) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_7), .A2(n_122), .B1(n_123), .B2(n_125), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g531 ( .A(n_8), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_9), .Y(n_115) );
AND2x2_ASAP7_75t_L g171 ( .A(n_10), .B(n_164), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_11), .Y(n_498) );
INVx2_ASAP7_75t_L g165 ( .A(n_12), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_13), .Y(n_124) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_14), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_14), .B(n_27), .Y(n_727) );
INVx1_ASAP7_75t_L g559 ( .A(n_15), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g817 ( .A1(n_16), .A2(n_27), .B1(n_781), .B2(n_818), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_16), .Y(n_818) );
AOI221x1_ASAP7_75t_L g218 ( .A1(n_17), .A2(n_142), .B1(n_219), .B2(n_221), .C(n_223), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_18), .B(n_160), .Y(n_193) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
INVx1_ASAP7_75t_L g557 ( .A(n_20), .Y(n_557) );
INVx1_ASAP7_75t_SL g480 ( .A(n_21), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_22), .B(n_161), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_23), .A2(n_142), .B(n_175), .Y(n_174) );
AOI221xp5_ASAP7_75t_SL g185 ( .A1(n_24), .A2(n_40), .B1(n_142), .B2(n_160), .C(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_25), .B(n_154), .Y(n_176) );
AOI33xp33_ASAP7_75t_L g517 ( .A1(n_26), .A2(n_53), .A3(n_208), .B1(n_214), .B2(n_518), .B3(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g781 ( .A(n_27), .Y(n_781) );
INVx1_ASAP7_75t_L g491 ( .A(n_28), .Y(n_491) );
OR2x2_ASAP7_75t_L g166 ( .A(n_29), .B(n_94), .Y(n_166) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_29), .A2(n_94), .B(n_165), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_30), .B(n_150), .Y(n_197) );
INVxp67_ASAP7_75t_L g217 ( .A(n_31), .Y(n_217) );
AND2x2_ASAP7_75t_L g248 ( .A(n_32), .B(n_163), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_33), .B(n_206), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_34), .A2(n_142), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_35), .B(n_150), .Y(n_187) );
AND2x2_ASAP7_75t_L g143 ( .A(n_36), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g158 ( .A(n_36), .B(n_147), .Y(n_158) );
INVx1_ASAP7_75t_L g213 ( .A(n_36), .Y(n_213) );
NOR3xp33_ASAP7_75t_L g113 ( .A(n_37), .B(n_114), .C(n_116), .Y(n_113) );
OR2x6_ASAP7_75t_L g791 ( .A(n_37), .B(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_38), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_39), .B(n_206), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_41), .A2(n_178), .B1(n_222), .B2(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_42), .B(n_549), .Y(n_548) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_43), .A2(n_84), .B1(n_142), .B2(n_211), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_44), .B(n_161), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_45), .B(n_154), .Y(n_246) );
INVx1_ASAP7_75t_L g789 ( .A(n_46), .Y(n_789) );
XNOR2xp5_ASAP7_75t_L g820 ( .A(n_47), .B(n_88), .Y(n_820) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_48), .B(n_198), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_49), .B(n_161), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_50), .Y(n_544) );
AND2x2_ASAP7_75t_L g235 ( .A(n_51), .B(n_163), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_52), .B(n_163), .Y(n_189) );
XOR2xp5_ASAP7_75t_L g812 ( .A(n_52), .B(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_54), .B(n_161), .Y(n_509) );
INVx1_ASAP7_75t_L g146 ( .A(n_55), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_55), .Y(n_156) );
AND2x2_ASAP7_75t_L g510 ( .A(n_56), .B(n_163), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g529 ( .A1(n_57), .A2(n_77), .B1(n_206), .B2(n_211), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_58), .B(n_206), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_59), .B(n_160), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_60), .A2(n_121), .B1(n_126), .B2(n_127), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_60), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_61), .B(n_222), .Y(n_500) );
AOI21xp5_ASAP7_75t_SL g469 ( .A1(n_62), .A2(n_211), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g167 ( .A(n_63), .B(n_163), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_64), .B(n_150), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_65), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_SL g200 ( .A(n_66), .B(n_164), .Y(n_200) );
INVx1_ASAP7_75t_L g554 ( .A(n_67), .Y(n_554) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_68), .B(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_69), .A2(n_142), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g508 ( .A(n_70), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_71), .B(n_150), .Y(n_177) );
AND2x2_ASAP7_75t_SL g285 ( .A(n_72), .B(n_198), .Y(n_285) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_73), .A2(n_211), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g144 ( .A(n_74), .Y(n_144) );
INVx1_ASAP7_75t_L g152 ( .A(n_74), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_75), .B(n_206), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_76), .Y(n_830) );
AND2x2_ASAP7_75t_L g482 ( .A(n_78), .B(n_221), .Y(n_482) );
INVx1_ASAP7_75t_L g555 ( .A(n_79), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_80), .A2(n_211), .B(n_479), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_81), .A2(n_211), .B(n_281), .C(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_82), .B(n_160), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_83), .A2(n_87), .B1(n_160), .B2(n_206), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_85), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g793 ( .A(n_85), .Y(n_793) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_86), .B(n_221), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_89), .A2(n_211), .B1(n_515), .B2(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_90), .B(n_154), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_91), .B(n_154), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_92), .B(n_795), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_93), .A2(n_142), .B(n_148), .Y(n_141) );
INVx1_ASAP7_75t_L g471 ( .A(n_95), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_96), .B(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g521 ( .A(n_97), .B(n_221), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_98), .A2(n_489), .B(n_490), .C(n_492), .Y(n_488) );
INVxp67_ASAP7_75t_L g220 ( .A(n_99), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_100), .B(n_160), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_101), .B(n_150), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_102), .A2(n_142), .B(n_195), .Y(n_194) );
BUFx2_ASAP7_75t_SL g787 ( .A(n_103), .Y(n_787) );
BUFx2_ASAP7_75t_L g804 ( .A(n_103), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_104), .B(n_161), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_117), .B(n_829), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_109), .Y(n_831) );
INVx3_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_SL g110 ( .A(n_111), .B(n_113), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_112), .B(n_793), .Y(n_792) );
HB1xp67_ASAP7_75t_L g130 ( .A(n_116), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g782 ( .A(n_116), .Y(n_782) );
OR2x2_ASAP7_75t_L g790 ( .A(n_116), .B(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_116), .B(n_798), .Y(n_797) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_805), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_783), .B(n_799), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_128), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g828 ( .A(n_120), .Y(n_828) );
INVxp33_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
INVx1_ASAP7_75t_L g125 ( .A(n_123), .Y(n_125) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
HB1xp67_ASAP7_75t_L g827 ( .A(n_129), .Y(n_827) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_457), .Y(n_129) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_396), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_289), .C(n_340), .Y(n_132) );
OAI211xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_179), .B(n_236), .C(n_267), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_168), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_138), .B(n_241), .Y(n_404) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g249 ( .A(n_139), .B(n_170), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_139), .B(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g266 ( .A(n_139), .B(n_256), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_139), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_139), .B(n_279), .Y(n_303) );
INVx2_ASAP7_75t_L g329 ( .A(n_139), .Y(n_329) );
AND2x4_ASAP7_75t_L g338 ( .A(n_139), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g443 ( .A(n_139), .B(n_310), .Y(n_443) );
AO21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_162), .B(n_167), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_159), .Y(n_140) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
BUFx3_ASAP7_75t_L g210 ( .A(n_143), .Y(n_210) );
AND2x6_ASAP7_75t_L g154 ( .A(n_144), .B(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g215 ( .A(n_144), .Y(n_215) );
AND2x4_ASAP7_75t_L g211 ( .A(n_145), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x4_ASAP7_75t_L g150 ( .A(n_146), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_147), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B(n_157), .Y(n_148) );
INVxp67_ASAP7_75t_L g560 ( .A(n_150), .Y(n_560) );
AND2x4_ASAP7_75t_L g161 ( .A(n_151), .B(n_155), .Y(n_161) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVxp67_ASAP7_75t_L g558 ( .A(n_154), .Y(n_558) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_157), .A2(n_176), .B(n_177), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_157), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_157), .A2(n_196), .B(n_197), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_157), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_157), .A2(n_245), .B(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_157), .A2(n_471), .B(n_472), .C(n_473), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_157), .A2(n_472), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_157), .A2(n_472), .B(n_508), .C(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g515 ( .A(n_157), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_157), .A2(n_472), .B(n_531), .C(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_157), .A2(n_547), .B(n_548), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_157), .B(n_178), .Y(n_561) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g160 ( .A(n_158), .B(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_158), .Y(n_492) );
INVx1_ASAP7_75t_L g225 ( .A(n_161), .Y(n_225) );
AO21x2_ASAP7_75t_L g241 ( .A1(n_162), .A2(n_242), .B(n_248), .Y(n_241) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_162), .A2(n_242), .B(n_248), .Y(n_256) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_162), .A2(n_476), .B(n_482), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_163), .Y(n_162) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_163), .A2(n_185), .B(n_189), .Y(n_184) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_165), .B(n_166), .Y(n_164) );
AND2x4_ASAP7_75t_L g178 ( .A(n_165), .B(n_166), .Y(n_178) );
AND2x2_ASAP7_75t_L g327 ( .A(n_168), .B(n_328), .Y(n_327) );
OAI32xp33_ASAP7_75t_L g410 ( .A1(n_168), .A2(n_332), .A3(n_336), .B1(n_343), .B2(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_168), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g264 ( .A(n_169), .B(n_265), .Y(n_264) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_169), .B(n_259), .C(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g363 ( .A(n_169), .B(n_266), .Y(n_363) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_170), .Y(n_253) );
INVx5_ASAP7_75t_L g288 ( .A(n_170), .Y(n_288) );
AND2x4_ASAP7_75t_L g344 ( .A(n_170), .B(n_256), .Y(n_344) );
OR2x2_ASAP7_75t_L g359 ( .A(n_170), .B(n_279), .Y(n_359) );
OR2x2_ASAP7_75t_L g385 ( .A(n_170), .B(n_241), .Y(n_385) );
AND2x2_ASAP7_75t_L g393 ( .A(n_170), .B(n_339), .Y(n_393) );
AND2x4_ASAP7_75t_SL g418 ( .A(n_170), .B(n_338), .Y(n_418) );
OR2x6_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_178), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_178), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_178), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_178), .B(n_220), .Y(n_219) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_178), .B(n_224), .C(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_178), .A2(n_469), .B(n_474), .Y(n_468) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_180), .B(n_338), .Y(n_414) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_190), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_181), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
OR2x6_ASAP7_75t_SL g238 ( .A(n_182), .B(n_239), .Y(n_238) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g263 ( .A(n_183), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_183), .B(n_298), .Y(n_316) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_183), .Y(n_454) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g271 ( .A(n_184), .Y(n_271) );
AND2x2_ASAP7_75t_L g296 ( .A(n_184), .B(n_227), .Y(n_296) );
INVx2_ASAP7_75t_L g324 ( .A(n_184), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_184), .B(n_191), .Y(n_365) );
BUFx3_ASAP7_75t_L g389 ( .A(n_184), .Y(n_389) );
OR2x2_ASAP7_75t_L g401 ( .A(n_184), .B(n_191), .Y(n_401) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_184), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_190), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_431) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_201), .Y(n_190) );
INVx1_ASAP7_75t_L g259 ( .A(n_191), .Y(n_259) );
OR2x2_ASAP7_75t_L g270 ( .A(n_191), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g277 ( .A(n_191), .Y(n_277) );
AND2x4_ASAP7_75t_SL g294 ( .A(n_191), .B(n_202), .Y(n_294) );
AND2x4_ASAP7_75t_L g299 ( .A(n_191), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g308 ( .A(n_191), .Y(n_308) );
OR2x2_ASAP7_75t_L g314 ( .A(n_191), .B(n_202), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_191), .B(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_191), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_191), .B(n_296), .Y(n_430) );
OR2x2_ASAP7_75t_L g446 ( .A(n_191), .B(n_349), .Y(n_446) );
OR2x6_ASAP7_75t_L g191 ( .A(n_192), .B(n_200), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_198), .Y(n_192) );
INVx2_ASAP7_75t_SL g281 ( .A(n_198), .Y(n_281) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_198), .A2(n_529), .B(n_533), .Y(n_528) );
BUFx4f_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx3_ASAP7_75t_L g222 ( .A(n_199), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_201), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g272 ( .A(n_201), .Y(n_272) );
AND2x2_ASAP7_75t_SL g379 ( .A(n_201), .B(n_263), .Y(n_379) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_226), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_202), .B(n_227), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_202), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_202), .B(n_271), .Y(n_275) );
INVx3_ASAP7_75t_L g300 ( .A(n_202), .Y(n_300) );
INVx1_ASAP7_75t_L g333 ( .A(n_202), .Y(n_333) );
AND2x2_ASAP7_75t_L g413 ( .A(n_202), .B(n_277), .Y(n_413) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_218), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_206), .B1(n_211), .B2(n_216), .Y(n_203) );
INVx1_ASAP7_75t_L g501 ( .A(n_206), .Y(n_501) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_210), .Y(n_206) );
INVx1_ASAP7_75t_L g542 ( .A(n_207), .Y(n_542) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
OR2x6_ASAP7_75t_L g472 ( .A(n_208), .B(n_215), .Y(n_472) );
INVxp33_ASAP7_75t_L g518 ( .A(n_208), .Y(n_518) );
INVx1_ASAP7_75t_L g543 ( .A(n_210), .Y(n_543) );
INVxp67_ASAP7_75t_L g499 ( .A(n_211), .Y(n_499) );
NOR2x1p5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
INVx1_ASAP7_75t_L g519 ( .A(n_214), .Y(n_519) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_221), .A2(n_488), .B1(n_493), .B2(n_494), .Y(n_487) );
INVx3_ASAP7_75t_L g494 ( .A(n_221), .Y(n_494) );
INVx4_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AOI21x1_ASAP7_75t_L g228 ( .A1(n_222), .A2(n_229), .B(n_235), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_222), .B(n_497), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_225), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_225), .A2(n_472), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_227), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g298 ( .A(n_227), .Y(n_298) );
AND2x2_ASAP7_75t_L g323 ( .A(n_227), .B(n_324), .Y(n_323) );
OR2x2_ASAP7_75t_L g349 ( .A(n_227), .B(n_271), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_227), .B(n_300), .Y(n_366) );
INVx1_ASAP7_75t_L g372 ( .A(n_227), .Y(n_372) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
AOI222xp33_ASAP7_75t_SL g236 ( .A1(n_237), .A2(n_240), .B1(n_250), .B2(n_257), .C1(n_260), .C2(n_264), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_249), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_241), .B(n_310), .Y(n_361) );
AND2x4_ASAP7_75t_L g377 ( .A(n_241), .B(n_288), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_247), .Y(n_242) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_252), .B(n_254), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g302 ( .A(n_253), .B(n_303), .Y(n_302) );
AOI222xp33_ASAP7_75t_L g267 ( .A1(n_254), .A2(n_268), .B1(n_273), .B2(n_278), .C1(n_286), .C2(n_833), .Y(n_267) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g406 ( .A(n_255), .B(n_310), .Y(n_406) );
OR2x2_ASAP7_75t_L g449 ( .A(n_255), .B(n_355), .Y(n_449) );
AND2x2_ASAP7_75t_L g278 ( .A(n_256), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g339 ( .A(n_256), .Y(n_339) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_256), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g367 ( .A1(n_257), .A2(n_368), .B(n_373), .C(n_374), .Y(n_367) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g395 ( .A(n_259), .Y(n_395) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g325 ( .A(n_264), .Y(n_325) );
AND2x2_ASAP7_75t_L g309 ( .A(n_265), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g318 ( .A(n_265), .B(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OAI31xp33_ASAP7_75t_L g360 ( .A1(n_268), .A2(n_286), .A3(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g362 ( .A1(n_269), .A2(n_319), .B(n_363), .C(n_364), .Y(n_362) );
OR2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
OR2x2_ASAP7_75t_L g351 ( .A(n_270), .B(n_300), .Y(n_351) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
BUFx2_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
AND2x2_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx6f_ASAP7_75t_L g310 ( .A(n_280), .Y(n_310) );
AOI21x1_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_285), .Y(n_280) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_281), .A2(n_513), .B(n_521), .Y(n_512) );
AO21x2_ASAP7_75t_L g572 ( .A1(n_281), .A2(n_513), .B(n_521), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_288), .B(n_345), .Y(n_437) );
OAI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_301), .B(n_304), .C(n_326), .Y(n_289) );
INVxp33_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_292), .B(n_297), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g330 ( .A(n_294), .B(n_323), .Y(n_330) );
OR2x2_ASAP7_75t_L g306 ( .A(n_295), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_310), .Y(n_336) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g412 ( .A(n_296), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g435 ( .A(n_297), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_299), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_299), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g447 ( .A(n_299), .B(n_323), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_299), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g390 ( .A(n_300), .B(n_372), .Y(n_390) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
AOI322xp5_ASAP7_75t_L g444 ( .A1(n_303), .A2(n_323), .A3(n_377), .B1(n_402), .B2(n_445), .C1(n_447), .C2(n_448), .Y(n_444) );
AOI211xp5_ASAP7_75t_SL g304 ( .A1(n_305), .A2(n_309), .B(n_311), .C(n_320), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_307), .B(n_335), .Y(n_357) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g322 ( .A(n_308), .B(n_323), .Y(n_322) );
NOR2x1p5_ASAP7_75t_L g388 ( .A(n_308), .B(n_389), .Y(n_388) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_308), .Y(n_421) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_309), .A2(n_327), .B(n_330), .C(n_331), .Y(n_326) );
AND2x4_ASAP7_75t_L g345 ( .A(n_310), .B(n_329), .Y(n_345) );
INVx2_ASAP7_75t_L g355 ( .A(n_310), .Y(n_355) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_310), .B(n_344), .Y(n_375) );
AND2x2_ASAP7_75t_L g417 ( .A(n_310), .B(n_418), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_310), .B(n_434), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_310), .B(n_338), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_315), .B(n_317), .Y(n_311) );
AND2x2_ASAP7_75t_L g407 ( .A(n_313), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g335 ( .A(n_316), .Y(n_335) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_325), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_328), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g422 ( .A(n_328), .Y(n_422) );
O2A1O1Ixp33_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_334), .B(n_336), .C(n_337), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_335), .Y(n_419) );
INVx3_ASAP7_75t_SL g434 ( .A(n_338), .Y(n_434) );
NAND5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_360), .C(n_367), .D(n_380), .E(n_391), .Y(n_340) );
AOI222xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_346), .B1(n_350), .B2(n_352), .C1(n_356), .C2(n_358), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_343), .A2(n_424), .B1(n_428), .B2(n_429), .Y(n_423) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g373 ( .A(n_344), .B(n_345), .Y(n_373) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_354), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_355), .B(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g392 ( .A(n_355), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g403 ( .A(n_355), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g433 ( .A(n_359), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g381 ( .A(n_366), .Y(n_381) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B(n_378), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_377), .A2(n_381), .B1(n_382), .B2(n_386), .Y(n_380) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g394 ( .A(n_379), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g399 ( .A(n_381), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_SL g427 ( .A(n_390), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_415), .C(n_438), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_414), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_405), .B2(n_407), .C(n_410), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g439 ( .A(n_401), .B(n_427), .Y(n_439) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
OAI321xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .A3(n_420), .B1(n_422), .B2(n_423), .C(n_431), .Y(n_415) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_429), .A2(n_451), .B1(n_455), .B2(n_456), .Y(n_450) );
INVx1_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B(n_444), .C(n_450), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_778), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_728), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_668), .B(n_727), .Y(n_459) );
NOR3xp33_ASAP7_75t_L g778 ( .A(n_460), .B(n_729), .C(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g823 ( .A(n_460), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_632), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_573), .C(n_602), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_463), .B(n_562), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_483), .B1(n_522), .B2(n_534), .Y(n_463) );
NAND2x1_ASAP7_75t_L g764 ( .A(n_464), .B(n_563), .Y(n_764) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
INVx2_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
INVx4_ASAP7_75t_L g578 ( .A(n_466), .Y(n_578) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_466), .Y(n_598) );
AND2x4_ASAP7_75t_L g609 ( .A(n_466), .B(n_577), .Y(n_609) );
AND2x2_ASAP7_75t_L g615 ( .A(n_466), .B(n_539), .Y(n_615) );
NOR2x1_ASAP7_75t_SL g688 ( .A(n_466), .B(n_550), .Y(n_688) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVxp67_ASAP7_75t_L g489 ( .A(n_472), .Y(n_489) );
INVx2_ASAP7_75t_L g549 ( .A(n_472), .Y(n_549) );
INVx2_ASAP7_75t_L g581 ( .A(n_475), .Y(n_581) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_475), .Y(n_595) );
INVx1_ASAP7_75t_L g606 ( .A(n_475), .Y(n_606) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_475), .Y(n_618) );
AND2x2_ASAP7_75t_L g650 ( .A(n_475), .B(n_550), .Y(n_650) );
INVx1_ASAP7_75t_L g676 ( .A(n_475), .Y(n_676) );
AND2x2_ASAP7_75t_L g738 ( .A(n_475), .B(n_566), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_502), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g631 ( .A(n_485), .B(n_570), .Y(n_631) );
INVx2_ASAP7_75t_L g673 ( .A(n_485), .Y(n_673) );
AND2x2_ASAP7_75t_L g775 ( .A(n_485), .B(n_502), .Y(n_775) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_486), .B(n_525), .Y(n_569) );
INVx2_ASAP7_75t_L g590 ( .A(n_486), .Y(n_590) );
AND2x4_ASAP7_75t_L g612 ( .A(n_486), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g647 ( .A(n_486), .Y(n_647) );
AND2x2_ASAP7_75t_L g771 ( .A(n_486), .B(n_528), .Y(n_771) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .Y(n_486) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_494), .A2(n_504), .B(n_510), .Y(n_503) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_494), .A2(n_504), .B(n_510), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_499), .B1(n_500), .B2(n_501), .Y(n_495) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g745 ( .A(n_502), .Y(n_745) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_511), .Y(n_502) );
NOR2xp67_ASAP7_75t_L g620 ( .A(n_503), .B(n_590), .Y(n_620) );
AND2x2_ASAP7_75t_L g625 ( .A(n_503), .B(n_590), .Y(n_625) );
INVx2_ASAP7_75t_L g638 ( .A(n_503), .Y(n_638) );
NOR2x1_ASAP7_75t_L g703 ( .A(n_503), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x4_ASAP7_75t_L g611 ( .A(n_511), .B(n_524), .Y(n_611) );
AND2x2_ASAP7_75t_L g626 ( .A(n_511), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g681 ( .A(n_511), .Y(n_681) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_512), .B(n_528), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_512), .B(n_525), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_514), .B(n_520), .Y(n_513) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVxp33_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
INVx3_ASAP7_75t_L g587 ( .A(n_524), .Y(n_587) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_525), .Y(n_585) );
AND2x2_ASAP7_75t_L g699 ( .A(n_525), .B(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g642 ( .A(n_526), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_526), .B(n_681), .Y(n_722) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g589 ( .A(n_527), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g570 ( .A(n_528), .B(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g613 ( .A(n_528), .Y(n_613) );
INVxp67_ASAP7_75t_L g627 ( .A(n_528), .Y(n_627) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_528), .Y(n_700) );
INVx1_ASAP7_75t_L g704 ( .A(n_528), .Y(n_704) );
INVx1_ASAP7_75t_L g682 ( .A(n_534), .Y(n_682) );
NOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_537), .Y(n_534) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_535), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g724 ( .A(n_536), .B(n_565), .Y(n_724) );
OR2x2_ASAP7_75t_L g776 ( .A(n_537), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g675 ( .A(n_538), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g711 ( .A(n_538), .B(n_598), .Y(n_711) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_550), .Y(n_538) );
AND2x4_ASAP7_75t_L g565 ( .A(n_539), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g577 ( .A(n_539), .Y(n_577) );
INVx2_ASAP7_75t_L g594 ( .A(n_539), .Y(n_594) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_539), .Y(n_720) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_545), .Y(n_539) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .C(n_544), .Y(n_541) );
INVx3_ASAP7_75t_L g566 ( .A(n_550), .Y(n_566) );
INVx2_ASAP7_75t_L g660 ( .A(n_550), .Y(n_660) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B(n_561), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_558), .B1(n_559), .B2(n_560), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_564), .B(n_640), .Y(n_657) );
NOR2x1_ASAP7_75t_L g749 ( .A(n_564), .B(n_578), .Y(n_749) );
INVx4_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_565), .B(n_640), .Y(n_726) );
AND2x2_ASAP7_75t_L g593 ( .A(n_566), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g607 ( .A(n_566), .Y(n_607) );
AOI22xp5_ASAP7_75t_SL g655 ( .A1(n_567), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g652 ( .A(n_568), .B(n_626), .Y(n_652) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g760 ( .A(n_569), .B(n_601), .Y(n_760) );
AND2x2_ASAP7_75t_L g583 ( .A(n_570), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g619 ( .A(n_570), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g762 ( .A(n_570), .B(n_673), .Y(n_762) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g637 ( .A(n_572), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g663 ( .A(n_572), .Y(n_663) );
AND2x2_ASAP7_75t_L g698 ( .A(n_572), .B(n_590), .Y(n_698) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_582), .B1(n_586), .B2(n_591), .C(n_596), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g654 ( .A(n_576), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_576), .B(n_650), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_576), .B(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NOR2xp67_ASAP7_75t_SL g622 ( .A(n_578), .B(n_623), .Y(n_622) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_578), .Y(n_635) );
AND2x4_ASAP7_75t_SL g719 ( .A(n_578), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g766 ( .A(n_578), .B(n_767), .Y(n_766) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx3_ASAP7_75t_L g640 ( .A(n_580), .Y(n_640) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_581), .Y(n_777) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI221x1_ASAP7_75t_L g730 ( .A1(n_583), .A2(n_731), .B1(n_733), .B2(n_734), .C(n_736), .Y(n_730) );
AND2x2_ASAP7_75t_L g656 ( .A(n_584), .B(n_612), .Y(n_656) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AND2x2_ASAP7_75t_L g599 ( .A(n_587), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_587), .B(n_589), .Y(n_773) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_593), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_593), .B(n_606), .Y(n_623) );
INVx2_ASAP7_75t_L g630 ( .A(n_593), .Y(n_630) );
INVx1_ASAP7_75t_L g692 ( .A(n_594), .Y(n_692) );
BUFx2_ASAP7_75t_L g712 ( .A(n_595), .Y(n_712) );
NAND2xp33_ASAP7_75t_SL g596 ( .A(n_597), .B(n_599), .Y(n_596) );
OR2x6_ASAP7_75t_L g629 ( .A(n_598), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g758 ( .A(n_598), .B(n_650), .Y(n_758) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_621), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_610), .B1(n_614), .B2(n_619), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_605), .B(n_609), .Y(n_667) );
AND2x4_ASAP7_75t_L g733 ( .A(n_605), .B(n_691), .Y(n_733) );
AND2x4_ASAP7_75t_SL g605 ( .A(n_606), .B(n_607), .Y(n_605) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_606), .Y(n_748) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_609), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_609), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_609), .B(n_640), .Y(n_732) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x2_ASAP7_75t_L g753 ( .A(n_611), .B(n_672), .Y(n_753) );
INVx3_ASAP7_75t_L g664 ( .A(n_612), .Y(n_664) );
AND2x2_ASAP7_75t_L g685 ( .A(n_612), .B(n_637), .Y(n_685) );
NAND2x1_ASAP7_75t_SL g756 ( .A(n_612), .B(n_663), .Y(n_756) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .B1(n_628), .B2(n_631), .Y(n_621) );
BUFx2_ASAP7_75t_L g677 ( .A(n_623), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_624), .A2(n_715), .B1(n_724), .B2(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_625), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g645 ( .A(n_626), .B(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_630), .B(n_710), .C(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
AOI211x1_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_641), .B(n_643), .C(n_661), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_636), .B(n_724), .Y(n_743) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_637), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g715 ( .A(n_637), .B(n_673), .Y(n_715) );
AND2x2_ASAP7_75t_L g770 ( .A(n_637), .B(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g693 ( .A(n_640), .Y(n_693) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g735 ( .A(n_642), .B(n_680), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_655), .Y(n_643) );
AOI22xp5_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_648), .B1(n_651), .B2(n_653), .Y(n_644) );
BUFx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g708 ( .A(n_647), .B(n_703), .Y(n_708) );
INVx1_ASAP7_75t_SL g750 ( .A(n_647), .Y(n_750) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_SL g718 ( .A(n_650), .B(n_719), .Y(n_718) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g754 ( .A(n_659), .B(n_676), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_666), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_663), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g678 ( .A(n_664), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_668), .Y(n_825) );
NAND3x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_705), .C(n_713), .Y(n_668) );
NAND4xp25_ASAP7_75t_L g779 ( .A(n_669), .B(n_705), .C(n_713), .D(n_780), .Y(n_779) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_670), .B(n_683), .Y(n_669) );
OAI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B1(n_677), .B2(n_678), .C1(n_680), .C2(n_682), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI21xp5_ASAP7_75t_SL g757 ( .A1(n_675), .A2(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_676), .B(n_691), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_679), .A2(n_737), .B1(n_739), .B2(n_740), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_694), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_687), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_693), .Y(n_689) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_691), .B(n_693), .Y(n_696) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B1(n_701), .B2(n_702), .Y(n_694) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
AND2x2_ASAP7_75t_L g702 ( .A(n_698), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_706), .B(n_709), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g739 ( .A(n_708), .Y(n_739) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_723), .Y(n_713) );
AOI22xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B1(n_718), .B2(n_721), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp33_ASAP7_75t_L g728 ( .A(n_727), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g824 ( .A(n_729), .Y(n_824) );
NAND3x1_ASAP7_75t_L g729 ( .A(n_730), .B(n_741), .C(n_761), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_733), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g767 ( .A(n_738), .Y(n_767) );
NOR2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_751), .Y(n_741) );
AOI21xp5_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_744), .B(n_750), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_757), .Y(n_751) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_756), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_765), .B2(n_768), .C(n_772), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVxp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B(n_776), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
INVxp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NOR3xp33_ASAP7_75t_L g826 ( .A(n_784), .B(n_827), .C(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_785), .B(n_794), .Y(n_784) );
INVxp33_ASAP7_75t_L g801 ( .A(n_785), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
CKINVDCx8_ASAP7_75t_R g786 ( .A(n_787), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_791), .Y(n_798) );
OAI32xp33_ASAP7_75t_L g799 ( .A1(n_791), .A2(n_800), .A3(n_801), .B1(n_802), .B2(n_834), .Y(n_799) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_794), .Y(n_800) );
INVx1_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NOR2x1_ASAP7_75t_R g803 ( .A(n_797), .B(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_800), .B(n_807), .Y(n_806) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g811 ( .A(n_804), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_812), .B(n_826), .Y(n_805) );
HB1xp67_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_809), .Y(n_808) );
BUFx3_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_814), .A2(n_815), .B1(n_821), .B2(n_822), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_819), .B2(n_820), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
AND3x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_824), .C(n_825), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
endmodule