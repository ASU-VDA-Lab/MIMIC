module real_aes_2932_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_0), .B(n_500), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_1), .A2(n_502), .B(n_503), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_2), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_3), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_4), .B(n_267), .Y(n_535) );
INVx1_ASAP7_75t_L g153 ( .A(n_5), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_6), .B(n_172), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_7), .B(n_267), .Y(n_562) );
INVx1_ASAP7_75t_L g236 ( .A(n_8), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_9), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_10), .Y(n_201) );
NAND2xp33_ASAP7_75t_L g524 ( .A(n_11), .B(n_264), .Y(n_524) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
AOI221x1_ASAP7_75t_L g568 ( .A1(n_13), .A2(n_26), .B1(n_500), .B2(n_502), .C(n_569), .Y(n_568) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_14), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_15), .B(n_500), .Y(n_520) );
INVx1_ASAP7_75t_L g265 ( .A(n_16), .Y(n_265) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_17), .A2(n_217), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_18), .B(n_176), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_19), .B(n_267), .Y(n_512) );
AO21x1_ASAP7_75t_L g530 ( .A1(n_20), .A2(n_500), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
INVx1_ASAP7_75t_L g262 ( .A(n_22), .Y(n_262) );
INVx1_ASAP7_75t_SL g182 ( .A(n_23), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_24), .B(n_159), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_25), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_27), .Y(n_787) );
AOI33xp33_ASAP7_75t_L g222 ( .A1(n_28), .A2(n_54), .A3(n_148), .B1(n_157), .B2(n_223), .B3(n_224), .Y(n_222) );
NAND2x1_ASAP7_75t_L g543 ( .A(n_29), .B(n_267), .Y(n_543) );
NAND2x1_ASAP7_75t_L g561 ( .A(n_30), .B(n_264), .Y(n_561) );
INVx1_ASAP7_75t_L g193 ( .A(n_31), .Y(n_193) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_32), .A2(n_86), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g173 ( .A(n_32), .B(n_86), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_33), .B(n_167), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_34), .B(n_264), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_35), .B(n_267), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_36), .B(n_264), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_37), .A2(n_502), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g147 ( .A(n_38), .Y(n_147) );
AND2x2_ASAP7_75t_L g165 ( .A(n_38), .B(n_153), .Y(n_165) );
AND2x2_ASAP7_75t_L g171 ( .A(n_38), .B(n_150), .Y(n_171) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_39), .B(n_107), .C(n_109), .Y(n_106) );
OR2x6_ASAP7_75t_L g122 ( .A(n_39), .B(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_40), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_41), .B(n_500), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_42), .B(n_167), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_43), .A2(n_140), .B1(n_172), .B2(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_44), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_45), .B(n_159), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_46), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_47), .B(n_264), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_48), .B(n_217), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_49), .B(n_159), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_50), .A2(n_502), .B(n_560), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_51), .Y(n_249) );
OAI222xp33_ASAP7_75t_L g125 ( .A1(n_52), .A2(n_126), .B1(n_783), .B2(n_784), .C1(n_787), .C2(n_788), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_52), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_53), .B(n_264), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_55), .B(n_159), .Y(n_212) );
INVx1_ASAP7_75t_L g152 ( .A(n_56), .Y(n_152) );
INVx1_ASAP7_75t_L g161 ( .A(n_56), .Y(n_161) );
AND2x2_ASAP7_75t_L g213 ( .A(n_57), .B(n_176), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g234 ( .A1(n_58), .A2(n_74), .B1(n_145), .B2(n_167), .C(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_59), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_60), .B(n_267), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_61), .B(n_140), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g144 ( .A1(n_62), .A2(n_145), .B(n_154), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_63), .A2(n_502), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g259 ( .A(n_64), .Y(n_259) );
AO21x1_ASAP7_75t_L g532 ( .A1(n_65), .A2(n_502), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_66), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g211 ( .A(n_67), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_68), .B(n_500), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_69), .A2(n_145), .B(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g554 ( .A(n_70), .B(n_177), .Y(n_554) );
INVx1_ASAP7_75t_L g150 ( .A(n_71), .Y(n_150) );
INVx1_ASAP7_75t_L g163 ( .A(n_71), .Y(n_163) );
AND2x2_ASAP7_75t_L g564 ( .A(n_72), .B(n_139), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_73), .B(n_167), .Y(n_225) );
AND2x2_ASAP7_75t_L g184 ( .A(n_75), .B(n_139), .Y(n_184) );
INVx1_ASAP7_75t_L g260 ( .A(n_76), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_77), .A2(n_145), .B(n_181), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_78), .A2(n_145), .B(n_216), .C(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g104 ( .A(n_79), .Y(n_104) );
AND2x2_ASAP7_75t_L g497 ( .A(n_80), .B(n_139), .Y(n_497) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_81), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_82), .B(n_500), .Y(n_514) );
OAI22xp5_ASAP7_75t_SL g798 ( .A1(n_83), .A2(n_488), .B1(n_799), .B2(n_800), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_83), .Y(n_799) );
AOI22xp5_ASAP7_75t_L g219 ( .A1(n_84), .A2(n_145), .B1(n_220), .B2(n_221), .Y(n_219) );
AND2x2_ASAP7_75t_L g531 ( .A(n_85), .B(n_172), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_87), .B(n_264), .Y(n_513) );
AND2x2_ASAP7_75t_L g546 ( .A(n_88), .B(n_139), .Y(n_546) );
INVx1_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_90), .B(n_267), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_91), .A2(n_502), .B(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_92), .B(n_264), .Y(n_570) );
AND2x2_ASAP7_75t_L g226 ( .A(n_93), .B(n_139), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_94), .B(n_267), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g190 ( .A1(n_95), .A2(n_191), .B(n_192), .C(n_195), .Y(n_190) );
INVx1_ASAP7_75t_SL g113 ( .A(n_96), .Y(n_113) );
BUFx2_ASAP7_75t_SL g796 ( .A(n_96), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_97), .A2(n_502), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_98), .B(n_159), .Y(n_158) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_110), .B(n_802), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_101), .Y(n_805) );
INVx3_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_106), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_104), .B(n_105), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_109), .B(n_121), .Y(n_120) );
OR2x6_ASAP7_75t_SL g487 ( .A(n_109), .B(n_121), .Y(n_487) );
AND2x6_ASAP7_75t_SL g782 ( .A(n_109), .B(n_122), .Y(n_782) );
OR2x2_ASAP7_75t_L g786 ( .A(n_109), .B(n_122), .Y(n_786) );
OA21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_125), .B(n_792), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_115), .A2(n_798), .B(n_801), .Y(n_797) );
NOR2xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_124), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_119), .Y(n_801) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_485), .B1(n_488), .B2(n_781), .Y(n_127) );
AOI22x1_ASAP7_75t_L g788 ( .A1(n_128), .A2(n_486), .B1(n_789), .B2(n_791), .Y(n_788) );
INVx1_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
AND3x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_375), .C(n_438), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_339), .Y(n_131) );
NOR3xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_280), .C(n_309), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g133 ( .A(n_134), .B(n_269), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_185), .B1(n_227), .B2(n_239), .Y(n_134) );
NAND2x1_ASAP7_75t_L g424 ( .A(n_135), .B(n_270), .Y(n_424) );
INVx2_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_174), .Y(n_136) );
INVx2_ASAP7_75t_L g241 ( .A(n_137), .Y(n_241) );
INVx4_ASAP7_75t_L g285 ( .A(n_137), .Y(n_285) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_137), .Y(n_305) );
AND2x4_ASAP7_75t_L g316 ( .A(n_137), .B(n_284), .Y(n_316) );
AND2x2_ASAP7_75t_L g322 ( .A(n_137), .B(n_244), .Y(n_322) );
NOR2x1_ASAP7_75t_SL g452 ( .A(n_137), .B(n_255), .Y(n_452) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_143), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_139), .A2(n_190), .B1(n_196), .B2(n_197), .Y(n_189) );
INVx3_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx4_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_140), .B(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx4f_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
AND2x4_ASAP7_75t_L g172 ( .A(n_142), .B(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_142), .B(n_173), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_166), .B(n_172), .Y(n_143) );
INVxp67_ASAP7_75t_L g202 ( .A(n_145), .Y(n_202) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_151), .Y(n_145) );
NOR2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx1_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OR2x6_ASAP7_75t_L g156 ( .A(n_149), .B(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g264 ( .A(n_150), .B(n_160), .Y(n_264) );
AND2x6_ASAP7_75t_L g502 ( .A(n_151), .B(n_171), .Y(n_502) );
AND2x2_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx2_ASAP7_75t_L g157 ( .A(n_152), .Y(n_157) );
AND2x4_ASAP7_75t_L g267 ( .A(n_152), .B(n_162), .Y(n_267) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_158), .C(n_164), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_SL g181 ( .A1(n_156), .A2(n_164), .B(n_182), .C(n_183), .Y(n_181) );
INVxp67_ASAP7_75t_L g191 ( .A(n_156), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_156), .A2(n_164), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_156), .A2(n_164), .B(n_236), .C(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g254 ( .A(n_156), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_156), .A2(n_194), .B1(n_259), .B2(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g168 ( .A(n_157), .B(n_169), .Y(n_168) );
INVxp33_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx1_ASAP7_75t_L g194 ( .A(n_159), .Y(n_194) );
AND2x4_ASAP7_75t_L g500 ( .A(n_159), .B(n_165), .Y(n_500) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_162), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g220 ( .A(n_164), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_164), .A2(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_164), .B(n_172), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_164), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_164), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_164), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_164), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_164), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_164), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_164), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_164), .A2(n_570), .B(n_571), .Y(n_569) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
INVx1_ASAP7_75t_L g204 ( .A(n_167), .Y(n_204) );
AND2x4_ASAP7_75t_L g167 ( .A(n_168), .B(n_170), .Y(n_167) );
INVx1_ASAP7_75t_L g247 ( .A(n_168), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_170), .Y(n_248) );
BUFx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_SL g508 ( .A(n_172), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_172), .A2(n_520), .B(n_521), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_172), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g288 ( .A(n_174), .Y(n_288) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_174), .Y(n_302) );
INVx1_ASAP7_75t_L g313 ( .A(n_174), .Y(n_313) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_174), .Y(n_325) );
AND2x2_ASAP7_75t_L g357 ( .A(n_174), .B(n_255), .Y(n_357) );
AND2x2_ASAP7_75t_L g389 ( .A(n_174), .B(n_273), .Y(n_389) );
INVx1_ASAP7_75t_L g396 ( .A(n_174), .Y(n_396) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_178), .B(n_184), .Y(n_174) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_175), .A2(n_558), .B(n_564), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_176), .A2(n_499), .B(n_501), .Y(n_498) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_176), .A2(n_568), .B(n_572), .Y(n_567) );
OA21x2_ASAP7_75t_L g607 ( .A1(n_176), .A2(n_568), .B(n_572), .Y(n_607) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_205), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g338 ( .A(n_187), .B(n_277), .Y(n_338) );
INVx2_ASAP7_75t_L g412 ( .A(n_187), .Y(n_412) );
AND2x2_ASAP7_75t_L g435 ( .A(n_187), .B(n_205), .Y(n_435) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_188), .B(n_230), .Y(n_276) );
INVx2_ASAP7_75t_L g297 ( .A(n_188), .Y(n_297) );
AND2x4_ASAP7_75t_L g319 ( .A(n_188), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g354 ( .A(n_188), .Y(n_354) );
AND2x2_ASAP7_75t_L g431 ( .A(n_188), .B(n_233), .Y(n_431) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_197), .A2(n_207), .B(n_213), .Y(n_206) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_197), .A2(n_207), .B(n_213), .Y(n_230) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_197), .A2(n_540), .B(n_546), .Y(n_539) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_197), .A2(n_548), .B(n_554), .Y(n_547) );
AO21x2_ASAP7_75t_L g575 ( .A1(n_197), .A2(n_540), .B(n_546), .Y(n_575) );
AO21x2_ASAP7_75t_L g593 ( .A1(n_197), .A2(n_548), .B(n_554), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g402 ( .A(n_205), .Y(n_402) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_214), .Y(n_205) );
NOR2xp67_ASAP7_75t_L g327 ( .A(n_206), .B(n_297), .Y(n_327) );
AND2x2_ASAP7_75t_L g332 ( .A(n_206), .B(n_297), .Y(n_332) );
INVx2_ASAP7_75t_L g345 ( .A(n_206), .Y(n_345) );
NOR2x1_ASAP7_75t_L g393 ( .A(n_206), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AND2x4_ASAP7_75t_L g318 ( .A(n_214), .B(n_229), .Y(n_318) );
AND2x2_ASAP7_75t_L g333 ( .A(n_214), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g386 ( .A(n_214), .Y(n_386) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_215), .B(n_233), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_215), .B(n_230), .Y(n_390) );
AO21x2_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_218), .B(n_226), .Y(n_215) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_216), .A2(n_218), .B(n_226), .Y(n_279) );
INVx2_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_217), .A2(n_234), .B(n_238), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_219), .B(n_225), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVxp33_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
INVx3_ASAP7_75t_L g294 ( .A(n_229), .Y(n_294) );
INVx3_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_230), .Y(n_292) );
AND2x2_ASAP7_75t_L g461 ( .A(n_230), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g349 ( .A(n_231), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_231), .B(n_386), .Y(n_481) );
BUFx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g296 ( .A(n_232), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x4_ASAP7_75t_L g277 ( .A(n_233), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g320 ( .A(n_233), .Y(n_320) );
INVxp67_ASAP7_75t_L g334 ( .A(n_233), .Y(n_334) );
INVx1_ASAP7_75t_L g394 ( .A(n_233), .Y(n_394) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_233), .Y(n_462) );
INVx1_ASAP7_75t_L g446 ( .A(n_239), .Y(n_446) );
NOR2x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NOR2x1_ASAP7_75t_L g366 ( .A(n_240), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g400 ( .A(n_241), .B(n_272), .Y(n_400) );
OR2x2_ASAP7_75t_L g436 ( .A(n_242), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g418 ( .A(n_243), .B(n_396), .Y(n_418) );
AND2x2_ASAP7_75t_L g470 ( .A(n_243), .B(n_305), .Y(n_470) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_255), .Y(n_243) );
AND2x4_ASAP7_75t_L g272 ( .A(n_244), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g284 ( .A(n_244), .Y(n_284) );
INVx2_ASAP7_75t_L g301 ( .A(n_244), .Y(n_301) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_244), .Y(n_479) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_250), .Y(n_244) );
NOR3xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .C(n_249), .Y(n_246) );
INVx3_ASAP7_75t_L g273 ( .A(n_255), .Y(n_273) );
INVx2_ASAP7_75t_L g367 ( .A(n_255), .Y(n_367) );
AND2x4_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_261), .B(n_268), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B1(n_265), .B2(n_266), .Y(n_261) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_274), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_271), .B(n_347), .Y(n_364) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_271), .B(n_285), .Y(n_406) );
INVx4_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_272), .B(n_347), .Y(n_484) );
AND2x2_ASAP7_75t_L g300 ( .A(n_273), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g314 ( .A(n_273), .Y(n_314) );
AOI22xp5_ASAP7_75t_SL g362 ( .A1(n_274), .A2(n_363), .B1(n_364), .B2(n_365), .Y(n_362) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_275), .B(n_333), .Y(n_359) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g420 ( .A(n_276), .B(n_308), .Y(n_420) );
AND2x2_ASAP7_75t_L g290 ( .A(n_277), .B(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g326 ( .A(n_277), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g422 ( .A(n_277), .B(n_412), .Y(n_422) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g344 ( .A(n_279), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g370 ( .A(n_279), .Y(n_370) );
AND2x2_ASAP7_75t_L g460 ( .A(n_279), .B(n_297), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_289), .B1(n_293), .B2(n_298), .C(n_303), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_L g361 ( .A(n_283), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_283), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_283), .B(n_357), .Y(n_476) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NOR2xp67_ASAP7_75t_SL g329 ( .A(n_285), .B(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_285), .Y(n_342) );
OR2x2_ASAP7_75t_L g426 ( .A(n_285), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_SL g478 ( .A(n_285), .B(n_479), .Y(n_478) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g347 ( .A(n_287), .Y(n_347) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_288), .Y(n_437) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI221x1_ASAP7_75t_L g377 ( .A1(n_290), .A2(n_378), .B1(n_380), .B2(n_383), .C(n_387), .Y(n_377) );
AND2x2_ASAP7_75t_L g363 ( .A(n_291), .B(n_319), .Y(n_363) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g306 ( .A(n_294), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_294), .B(n_296), .Y(n_433) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
AND2x2_ASAP7_75t_SL g304 ( .A(n_300), .B(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_300), .B(n_313), .Y(n_330) );
INVx2_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
INVx1_ASAP7_75t_L g382 ( .A(n_301), .Y(n_382) );
BUFx2_ASAP7_75t_L g471 ( .A(n_302), .Y(n_471) );
NAND2xp33_ASAP7_75t_SL g303 ( .A(n_304), .B(n_306), .Y(n_303) );
OR2x6_ASAP7_75t_L g336 ( .A(n_305), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g417 ( .A(n_305), .B(n_357), .Y(n_417) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_328), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_317), .B1(n_321), .B2(n_326), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_312), .B(n_316), .Y(n_374) );
AND2x4_ASAP7_75t_L g380 ( .A(n_312), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_SL g312 ( .A(n_313), .B(n_314), .Y(n_312) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_313), .Y(n_405) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_316), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_316), .B(n_347), .Y(n_379) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_316), .Y(n_463) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g410 ( .A(n_318), .B(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
NAND2x1_ASAP7_75t_SL g415 ( .A(n_319), .B(n_370), .Y(n_415) );
AND2x2_ASAP7_75t_L g449 ( .A(n_319), .B(n_344), .Y(n_449) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_331), .B1(n_335), .B2(n_338), .Y(n_328) );
BUFx2_ASAP7_75t_L g444 ( .A(n_330), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_331), .A2(n_400), .B1(n_474), .B2(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_332), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g352 ( .A(n_333), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_337), .B(n_469), .C(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
AOI211x1_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_348), .B(n_350), .C(n_368), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_343), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AND2x2_ASAP7_75t_L g430 ( .A(n_344), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_344), .B(n_411), .Y(n_442) );
AND2x2_ASAP7_75t_L g474 ( .A(n_344), .B(n_412), .Y(n_474) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g455 ( .A(n_347), .Y(n_455) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g384 ( .A(n_349), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_362), .Y(n_350) );
AOI22xp5_ASAP7_75t_SL g351 ( .A1(n_352), .A2(n_355), .B1(n_358), .B2(n_360), .Y(n_351) );
BUFx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g392 ( .A(n_354), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g407 ( .A(n_354), .Y(n_407) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_357), .B(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g413 ( .A(n_366), .B(n_396), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_372), .B(n_373), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_370), .B(n_392), .Y(n_467) );
OR2x2_ASAP7_75t_L g445 ( .A(n_371), .B(n_390), .Y(n_445) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND3x1_ASAP7_75t_L g376 ( .A(n_377), .B(n_397), .C(n_421), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_380), .A2(n_410), .B1(n_413), .B2(n_414), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_381), .B(n_396), .Y(n_395) );
INVx2_ASAP7_75t_SL g454 ( .A(n_381), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_381), .B(n_455), .Y(n_458) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI222xp33_ASAP7_75t_L g441 ( .A1(n_385), .A2(n_442), .B1(n_443), .B2(n_444), .C1(n_445), .C2(n_446), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .B1(n_391), .B2(n_395), .Y(n_387) );
INVx1_ASAP7_75t_SL g427 ( .A(n_389), .Y(n_427) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g464 ( .A(n_393), .B(n_460), .Y(n_464) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_408), .Y(n_397) );
AOI21xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_401), .B(n_407), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_416), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_415), .B(n_429), .Y(n_428) );
OAI21xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g443 ( .A(n_418), .Y(n_443) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_425), .B2(n_428), .C(n_432), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_434), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NAND3x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_465), .C(n_472), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_447), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_456), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_449), .B(n_450), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_451), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_459), .B1(n_463), .B2(n_464), .Y(n_456) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_466), .B(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
AOI22xp5_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_475), .B1(n_477), .B2(n_480), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
CKINVDCx11_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g800 ( .A(n_488), .Y(n_800) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g791 ( .A(n_489), .Y(n_791) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_690), .Y(n_489) );
NOR4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_608), .C(n_634), .D(n_674), .Y(n_490) );
OAI211xp5_ASAP7_75t_SL g491 ( .A1(n_492), .A2(n_525), .B(n_555), .C(n_594), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_506), .Y(n_493) );
AND2x2_ASAP7_75t_L g761 ( .A(n_494), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_495), .B(n_506), .Y(n_628) );
BUFx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_496), .B(n_581), .Y(n_580) );
INVx5_ASAP7_75t_L g614 ( .A(n_496), .Y(n_614) );
NOR2x1_ASAP7_75t_SL g656 ( .A(n_496), .B(n_507), .Y(n_656) );
AND2x2_ASAP7_75t_L g712 ( .A(n_496), .B(n_518), .Y(n_712) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_507), .B(n_518), .Y(n_584) );
AND2x2_ASAP7_75t_L g645 ( .A(n_507), .B(n_614), .Y(n_645) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_508), .B(n_516), .Y(n_515) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_508), .A2(n_509), .B(n_515), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
AND2x2_ASAP7_75t_L g657 ( .A(n_517), .B(n_581), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_517), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g701 ( .A(n_517), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g734 ( .A(n_517), .B(n_556), .Y(n_734) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g578 ( .A(n_518), .Y(n_578) );
AND2x2_ASAP7_75t_L g611 ( .A(n_518), .B(n_612), .Y(n_611) );
BUFx3_ASAP7_75t_L g646 ( .A(n_518), .Y(n_646) );
OR2x2_ASAP7_75t_L g722 ( .A(n_518), .B(n_581), .Y(n_722) );
INVx1_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
AOI211x1_ASAP7_75t_SL g651 ( .A1(n_527), .A2(n_643), .B(n_652), .C(n_654), .Y(n_651) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_527), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_527), .B(n_694), .Y(n_741) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g591 ( .A(n_528), .Y(n_591) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g566 ( .A(n_529), .Y(n_566) );
OAI21x1_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_532), .B(n_536), .Y(n_529) );
INVx1_ASAP7_75t_L g537 ( .A(n_531), .Y(n_537) );
AOI322xp5_ASAP7_75t_L g555 ( .A1(n_538), .A2(n_556), .A3(n_565), .B1(n_573), .B2(n_576), .C1(n_582), .C2(n_585), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_538), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_547), .Y(n_538) );
INVx2_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
INVxp67_ASAP7_75t_L g631 ( .A(n_539), .Y(n_631) );
BUFx3_ASAP7_75t_L g695 ( .A(n_539), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
INVx2_ASAP7_75t_L g604 ( .A(n_547), .Y(n_604) );
AND2x2_ASAP7_75t_L g653 ( .A(n_547), .B(n_567), .Y(n_653) );
AND2x2_ASAP7_75t_L g697 ( .A(n_547), .B(n_606), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_549), .B(n_553), .Y(n_548) );
AND2x2_ASAP7_75t_L g582 ( .A(n_556), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_556), .B(n_767), .Y(n_766) );
AND2x2_ASAP7_75t_SL g776 ( .A(n_556), .B(n_611), .Y(n_776) );
INVx4_ASAP7_75t_L g581 ( .A(n_557), .Y(n_581) );
AND2x2_ASAP7_75t_L g613 ( .A(n_557), .B(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_557), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_565), .B(n_650), .Y(n_675) );
INVx1_ASAP7_75t_SL g714 ( .A(n_565), .Y(n_714) );
AND2x4_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x4_ASAP7_75t_L g605 ( .A(n_566), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_566), .B(n_604), .Y(n_673) );
AND2x2_ASAP7_75t_L g725 ( .A(n_566), .B(n_575), .Y(n_725) );
OR2x2_ASAP7_75t_L g749 ( .A(n_566), .B(n_567), .Y(n_749) );
AND2x2_ASAP7_75t_L g573 ( .A(n_567), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g623 ( .A(n_567), .B(n_604), .Y(n_623) );
AND2x2_ASAP7_75t_SL g679 ( .A(n_567), .B(n_591), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_573), .B(n_686), .Y(n_703) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g638 ( .A(n_575), .Y(n_638) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_575), .B(n_592), .Y(n_678) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_579), .Y(n_576) );
OR2x2_ASAP7_75t_L g626 ( .A(n_577), .B(n_580), .Y(n_626) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g595 ( .A(n_578), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g743 ( .A(n_578), .B(n_656), .Y(n_743) );
AND2x2_ASAP7_75t_L g759 ( .A(n_578), .B(n_613), .Y(n_759) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI311xp33_ASAP7_75t_L g729 ( .A1(n_580), .A2(n_668), .A3(n_730), .B(n_732), .C(n_739), .Y(n_729) );
AND2x4_ASAP7_75t_L g596 ( .A(n_581), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g600 ( .A(n_581), .Y(n_600) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_581), .B(n_614), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_581), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g713 ( .A(n_581), .B(n_700), .Y(n_713) );
AND2x2_ASAP7_75t_L g599 ( .A(n_583), .B(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_584), .Y(n_617) );
OR2x2_ASAP7_75t_L g706 ( .A(n_584), .B(n_670), .Y(n_706) );
INVx1_ASAP7_75t_L g762 ( .A(n_584), .Y(n_762) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g671 ( .A(n_588), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g685 ( .A(n_588), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g760 ( .A(n_588), .B(n_633), .Y(n_760) );
BUFx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g603 ( .A(n_589), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g622 ( .A(n_589), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g684 ( .A(n_590), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_590), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x2_ASAP7_75t_L g633 ( .A(n_591), .B(n_604), .Y(n_633) );
AND2x4_ASAP7_75t_L g686 ( .A(n_591), .B(n_593), .Y(n_686) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI21xp33_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_599), .B(n_601), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_595), .A2(n_681), .B1(n_685), .B2(n_687), .Y(n_680) );
AND2x2_ASAP7_75t_SL g640 ( .A(n_596), .B(n_614), .Y(n_640) );
INVx2_ASAP7_75t_L g702 ( .A(n_596), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_596), .B(n_712), .Y(n_716) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g612 ( .A(n_598), .Y(n_612) );
INVx1_ASAP7_75t_L g665 ( .A(n_598), .Y(n_665) );
INVx1_ASAP7_75t_L g616 ( .A(n_600), .Y(n_616) );
AND3x2_ASAP7_75t_L g644 ( .A(n_600), .B(n_645), .C(n_646), .Y(n_644) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g708 ( .A(n_603), .Y(n_708) );
AND2x2_ASAP7_75t_L g636 ( .A(n_605), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g707 ( .A(n_605), .B(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_605), .A2(n_719), .B1(n_723), .B2(n_726), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_605), .B(n_753), .Y(n_757) );
BUFx2_ASAP7_75t_L g648 ( .A(n_606), .Y(n_648) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g619 ( .A(n_607), .Y(n_619) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_607), .Y(n_738) );
OAI221xp5_ASAP7_75t_SL g608 ( .A1(n_609), .A2(n_618), .B1(n_620), .B2(n_621), .C(n_624), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_615), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_L g700 ( .A(n_612), .Y(n_700) );
INVx2_ASAP7_75t_SL g689 ( .A(n_613), .Y(n_689) );
AND2x2_ASAP7_75t_L g771 ( .A(n_613), .B(n_638), .Y(n_771) );
INVx4_ASAP7_75t_L g662 ( .A(n_614), .Y(n_662) );
INVx1_ASAP7_75t_L g620 ( .A(n_615), .Y(n_620) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x4_ASAP7_75t_L g731 ( .A(n_619), .B(n_686), .Y(n_731) );
INVx1_ASAP7_75t_SL g770 ( .A(n_619), .Y(n_770) );
AND2x2_ASAP7_75t_L g775 ( .A(n_619), .B(n_678), .Y(n_775) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g717 ( .A(n_623), .Y(n_717) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_627), .B(n_629), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
INVx1_ASAP7_75t_L g650 ( .A(n_631), .Y(n_650) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g647 ( .A(n_633), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g737 ( .A(n_633), .B(n_738), .Y(n_737) );
OAI211xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_639), .B(n_641), .C(n_658), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g730 ( .A(n_637), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_638), .B(n_653), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_638), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g763 ( .A(n_638), .B(n_686), .Y(n_763) );
OAI221xp5_ASAP7_75t_SL g674 ( .A1(n_639), .A2(n_663), .B1(n_675), .B2(n_676), .C(n_680), .Y(n_674) );
INVx3_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g745 ( .A(n_640), .B(n_646), .Y(n_745) );
OAI32xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_647), .A3(n_649), .B1(n_651), .B2(n_655), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_645), .Y(n_735) );
INVx2_ASAP7_75t_L g668 ( .A(n_646), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_646), .A2(n_698), .B(n_778), .C(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g683 ( .A(n_648), .Y(n_683) );
OR2x2_ASAP7_75t_L g779 ( .A(n_648), .B(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_652), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g740 ( .A(n_655), .Y(n_740) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g721 ( .A(n_656), .Y(n_721) );
OAI21xp33_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_667), .B(n_671), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
OR2x2_ASAP7_75t_L g698 ( .A(n_661), .B(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_662), .B(n_665), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_664), .A2(n_696), .B1(n_765), .B2(n_768), .C(n_772), .Y(n_764) );
INVx2_ASAP7_75t_L g767 ( .A(n_664), .Y(n_767) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OR2x2_ASAP7_75t_L g688 ( .A(n_668), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g755 ( .A(n_668), .B(n_713), .Y(n_755) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVxp67_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
INVx1_ASAP7_75t_L g753 ( .A(n_678), .Y(n_753) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_686), .B(n_716), .Y(n_773) );
INVx2_ASAP7_75t_L g780 ( .A(n_686), .Y(n_780) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_688), .A2(n_751), .B1(n_754), .B2(n_756), .C(n_758), .Y(n_750) );
AND5x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_729), .C(n_744), .D(n_764), .E(n_774), .Y(n_690) );
NOR2xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_709), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_698), .B1(n_701), .B2(n_703), .C(n_704), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI221xp5_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_714), .B1(n_715), .B2(n_717), .C(n_718), .Y(n_709) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_714), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
OR2x2_ASAP7_75t_L g727 ( .A(n_722), .B(n_728), .Y(n_727) );
CKINVDCx16_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx2_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_735), .B(n_736), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B(n_750), .Y(n_744) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVxp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B1(n_761), .B2(n_763), .Y(n_758) );
O2A1O1Ixp33_ASAP7_75t_L g774 ( .A1(n_760), .A2(n_775), .B(n_776), .C(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_L g778 ( .A(n_771), .Y(n_778) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx11_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_782), .Y(n_790) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx3_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx3_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
CKINVDCx11_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
CKINVDCx8_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
endmodule