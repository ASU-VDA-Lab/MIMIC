module fake_jpeg_8794_n_295 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx13_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_45),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_0),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_28),
.C(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_25),
.B(n_17),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_48),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_48),
.A2(n_37),
.B1(n_19),
.B2(n_33),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_55),
.B(n_59),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_48),
.B1(n_47),
.B2(n_33),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_76),
.B1(n_21),
.B2(n_27),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_38),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_0),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_19),
.B1(n_37),
.B2(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_46),
.B1(n_27),
.B2(n_34),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_37),
.B1(n_29),
.B2(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_70),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_29),
.B1(n_18),
.B2(n_35),
.Y(n_59)
);

INVxp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_18),
.B1(n_35),
.B2(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_66),
.B1(n_75),
.B2(n_46),
.Y(n_91)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_20),
.B1(n_24),
.B2(n_32),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_24),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_44),
.Y(n_82)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_41),
.B(n_30),
.C(n_23),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_78),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_84),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_40),
.C(n_44),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_97),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_84),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_46),
.B1(n_36),
.B2(n_34),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_90),
.A2(n_77),
.B1(n_1),
.B2(n_4),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_106),
.B1(n_1),
.B2(n_40),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_67),
.B1(n_65),
.B2(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_70),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_13),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_51),
.B(n_44),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_109),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_40),
.B(n_44),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_54),
.A2(n_46),
.B1(n_36),
.B2(n_31),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_65),
.B1(n_75),
.B2(n_69),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_100),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_77),
.B1(n_71),
.B2(n_40),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_12),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_36),
.B1(n_31),
.B2(n_2),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_57),
.A2(n_36),
.B1(n_31),
.B2(n_3),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_11),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_11),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_39),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_0),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_1),
.Y(n_140)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_67),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_67),
.B1(n_69),
.B2(n_75),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_133),
.B1(n_136),
.B2(n_102),
.Y(n_149)
);

CKINVDCx6p67_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_140),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_1),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_95),
.B(n_96),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_134),
.B(n_145),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_135),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_12),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_88),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_93),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_80),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_147),
.B(n_151),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_148),
.B(n_152),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_159),
.B1(n_172),
.B2(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_79),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_79),
.Y(n_154)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_111),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_155),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_166),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_86),
.B1(n_85),
.B2(n_79),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_81),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_78),
.Y(n_180)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_168),
.B(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_97),
.B(n_112),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_130),
.B(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_99),
.B1(n_83),
.B2(n_92),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_173),
.A2(n_114),
.B1(n_87),
.B2(n_101),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_118),
.A2(n_114),
.B1(n_101),
.B2(n_94),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_115),
.A2(n_114),
.B1(n_101),
.B2(n_81),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_105),
.B1(n_87),
.B2(n_104),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_141),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_138),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_132),
.B1(n_115),
.B2(n_136),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_187),
.B1(n_195),
.B2(n_204),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_154),
.C(n_150),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_185),
.C(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_182),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_125),
.C(n_144),
.Y(n_181)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_158),
.C(n_156),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_130),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_175),
.C(n_160),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_121),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_193),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_159),
.A2(n_120),
.B(n_142),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_192),
.B(n_197),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_167),
.B(n_120),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_131),
.B1(n_146),
.B2(n_101),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_143),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_147),
.C(n_172),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_177),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_173),
.A2(n_113),
.B1(n_98),
.B2(n_129),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_176),
.B1(n_157),
.B2(n_149),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_224),
.B(n_195),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_169),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_211),
.C(n_205),
.Y(n_243)
);

OAI21xp33_ASAP7_75t_SL g244 ( 
.A1(n_212),
.A2(n_185),
.B(n_14),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_189),
.A2(n_161),
.B1(n_158),
.B2(n_148),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_213),
.A2(n_214),
.B1(n_227),
.B2(n_191),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_161),
.B1(n_152),
.B2(n_168),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_156),
.C(n_177),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_14),
.C(n_17),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_219),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_221),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_8),
.B(n_12),
.C(n_14),
.D(n_15),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_226),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_178),
.A2(n_162),
.B(n_98),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_162),
.B1(n_15),
.B2(n_16),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_207),
.B1(n_224),
.B2(n_215),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_228),
.A2(n_225),
.B1(n_217),
.B2(n_216),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_230),
.A2(n_234),
.B1(n_239),
.B2(n_218),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_196),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_205),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_192),
.B(n_184),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_17),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_184),
.B(n_183),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_236),
.B1(n_241),
.B2(n_223),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_183),
.B1(n_194),
.B2(n_198),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_194),
.B(n_198),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_181),
.B1(n_196),
.B2(n_201),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_245),
.C(n_219),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_240),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_259),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_233),
.B1(n_255),
.B2(n_261),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g250 ( 
.A(n_242),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_253),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_256),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_240),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_254),
.Y(n_272)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_231),
.C(n_243),
.Y(n_266)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_258),
.A2(n_261),
.B1(n_236),
.B2(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_228),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_266),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_230),
.B1(n_239),
.B2(n_232),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_265),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g267 ( 
.A(n_248),
.B(n_234),
.CI(n_241),
.CON(n_267),
.SN(n_267)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_269),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_273),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_245),
.C(n_246),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_269),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_267),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_253),
.B(n_258),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_278),
.A2(n_267),
.B(n_273),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_270),
.A2(n_252),
.B1(n_249),
.B2(n_259),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_272),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_281),
.B(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_280),
.B(n_264),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_283),
.A2(n_284),
.B(n_285),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_268),
.B1(n_266),
.B2(n_257),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_286),
.A2(n_276),
.B(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_277),
.C(n_268),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_287),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_291),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_277),
.Y(n_295)
);


endmodule