module fake_netlist_1_1060_n_698 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_698);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_698;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_55), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_53), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_63), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_44), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_26), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_21), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_3), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_62), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_69), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_50), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_11), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_29), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_14), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_12), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_7), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_4), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_51), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_12), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_38), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_37), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_65), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_11), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_60), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_4), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_52), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_47), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_64), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_58), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_18), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_49), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_0), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_9), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_40), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_2), .Y(n_116) );
OR2x2_ASAP7_75t_L g117 ( .A(n_71), .B(n_77), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_5), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_22), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_74), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_0), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_28), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_25), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_98), .A2(n_1), .B1(n_3), .B2(n_5), .Y(n_126) );
AND2x6_ASAP7_75t_L g127 ( .A(n_87), .B(n_35), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_80), .B(n_6), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
BUFx12f_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_124), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_112), .B(n_6), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_124), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_115), .B(n_7), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_78), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_112), .B(n_8), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_79), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_88), .B(n_8), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_93), .B(n_10), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_93), .B(n_10), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_95), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_97), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
CKINVDCx8_ASAP7_75t_R g149 ( .A(n_82), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_85), .B(n_13), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_89), .B(n_13), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_101), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_89), .B(n_14), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_86), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_125), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_96), .B(n_15), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_106), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_109), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_111), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_118), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_92), .B(n_15), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_103), .B(n_16), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_119), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_117), .B(n_42), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_121), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_122), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_127), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_153), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_130), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_153), .Y(n_172) );
OR2x2_ASAP7_75t_L g173 ( .A(n_136), .B(n_91), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_140), .B(n_92), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_127), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_130), .A2(n_123), .B1(n_120), .B2(n_102), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_159), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_131), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_140), .B(n_102), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_163), .B(n_105), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_146), .B(n_108), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_131), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_146), .B(n_108), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_147), .B(n_82), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_163), .B(n_117), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_136), .B(n_110), .Y(n_195) );
CKINVDCx11_ASAP7_75t_R g196 ( .A(n_149), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_163), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_159), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_147), .B(n_83), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_134), .B(n_113), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_135), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_134), .B(n_83), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_135), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
AND2x6_ASAP7_75t_L g211 ( .A(n_155), .B(n_116), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_154), .B(n_104), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_149), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_154), .B(n_114), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_127), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_161), .B(n_114), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_161), .B(n_99), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_165), .B(n_90), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_160), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_165), .B(n_84), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_127), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_138), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_159), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_135), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_150), .Y(n_229) );
AND2x6_ASAP7_75t_L g230 ( .A(n_155), .B(n_107), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_127), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_150), .Y(n_232) );
BUFx4f_ASAP7_75t_L g233 ( .A(n_211), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_176), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_210), .B(n_128), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g236 ( .A1(n_211), .A2(n_127), .B1(n_132), .B2(n_129), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_208), .Y(n_237) );
AO22x1_ASAP7_75t_L g238 ( .A1(n_230), .A2(n_126), .B1(n_127), .B2(n_84), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_225), .B(n_166), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_196), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_208), .B(n_166), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_217), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_217), .B(n_142), .Y(n_243) );
NOR2xp67_ASAP7_75t_L g244 ( .A(n_173), .B(n_144), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_214), .B(n_148), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_202), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_211), .A2(n_132), .B1(n_129), .B2(n_143), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_173), .B(n_166), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_214), .B(n_220), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_214), .B(n_148), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_203), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_220), .B(n_221), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_170), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_205), .Y(n_254) );
NAND3xp33_ASAP7_75t_SL g255 ( .A(n_171), .B(n_107), .C(n_120), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_194), .A2(n_126), .B1(n_151), .B2(n_164), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_220), .B(n_137), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_221), .B(n_143), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_177), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_221), .B(n_137), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_176), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_230), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_177), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_195), .B(n_158), .Y(n_266) );
INVx1_ASAP7_75t_SL g267 ( .A(n_196), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_218), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_180), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_169), .B(n_168), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_218), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_169), .B(n_168), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_172), .Y(n_274) );
AND3x2_ASAP7_75t_SL g275 ( .A(n_183), .B(n_123), .C(n_139), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_175), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_174), .B(n_139), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_180), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_185), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_207), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_194), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_204), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_185), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_231), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_219), .B(n_168), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_174), .B(n_168), .Y(n_287) );
INVx5_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_187), .B(n_168), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_211), .A2(n_162), .B1(n_160), .B2(n_167), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_187), .B(n_162), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_204), .B(n_167), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_189), .B(n_167), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_230), .A2(n_167), .B1(n_162), .B2(n_160), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_204), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_212), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_188), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_195), .B(n_162), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_188), .B(n_167), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_188), .Y(n_300) );
BUFx4f_ASAP7_75t_L g301 ( .A(n_281), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_295), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_268), .Y(n_303) );
INVx5_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_268), .Y(n_305) );
AO21x1_ASAP7_75t_L g306 ( .A1(n_293), .A2(n_212), .B(n_213), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_253), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_262), .B(n_182), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_281), .B(n_198), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_262), .B(n_197), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_283), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_249), .B(n_169), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_248), .A2(n_230), .B1(n_191), .B2(n_192), .Y(n_316) );
AO21x1_ASAP7_75t_L g317 ( .A1(n_293), .A2(n_213), .B(n_216), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_249), .B(n_215), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
INVx5_ASAP7_75t_L g320 ( .A(n_288), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_235), .B(n_201), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_259), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_288), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_288), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_233), .Y(n_325) );
AOI21xp33_ASAP7_75t_L g326 ( .A1(n_266), .A2(n_223), .B(n_199), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_253), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_243), .B(n_230), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_244), .B(n_230), .Y(n_329) );
INVx5_ASAP7_75t_L g330 ( .A(n_259), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_249), .A2(n_199), .B1(n_226), .B2(n_184), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_253), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_259), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_259), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_233), .B(n_231), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_233), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_274), .Y(n_338) );
AOI22xp5_ASAP7_75t_L g339 ( .A1(n_256), .A2(n_215), .B1(n_184), .B2(n_226), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_242), .B(n_162), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_298), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_265), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_265), .Y(n_343) );
OAI22x1_ASAP7_75t_L g344 ( .A1(n_275), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_274), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_239), .B(n_160), .Y(n_346) );
BUFx8_ASAP7_75t_SL g347 ( .A(n_240), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_274), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_247), .B(n_222), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_277), .B(n_222), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_277), .Y(n_351) );
NAND3xp33_ASAP7_75t_L g352 ( .A(n_236), .B(n_216), .C(n_222), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_265), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_304), .B(n_237), .Y(n_354) );
CKINVDCx6p67_ASAP7_75t_R g355 ( .A(n_311), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_304), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_321), .B(n_277), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_304), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_301), .A2(n_247), .B1(n_241), .B2(n_236), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_304), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_347), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_301), .A2(n_255), .B1(n_240), .B2(n_267), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_301), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g364 ( .A1(n_326), .A2(n_257), .B1(n_252), .B2(n_238), .C(n_245), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_304), .B(n_245), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_328), .A2(n_264), .B1(n_245), .B2(n_287), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_328), .A2(n_287), .B1(n_289), .B2(n_276), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_318), .A2(n_287), .B1(n_289), .B2(n_276), .Y(n_368) );
INVx4_ASAP7_75t_SL g369 ( .A(n_308), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_308), .B(n_276), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_318), .A2(n_289), .B1(n_257), .B2(n_299), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_327), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_352), .A2(n_272), .B(n_270), .Y(n_373) );
O2A1O1Ixp33_ASAP7_75t_SL g374 ( .A1(n_329), .A2(n_272), .B(n_270), .C(n_294), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_307), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_327), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_SL g377 ( .A1(n_346), .A2(n_246), .B(n_280), .C(n_251), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_311), .B(n_254), .Y(n_378) );
CKINVDCx5p33_ASAP7_75t_R g379 ( .A(n_347), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_318), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_302), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_339), .B(n_250), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g383 ( .A1(n_316), .A2(n_261), .B(n_258), .C(n_341), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g384 ( .A1(n_351), .A2(n_275), .B1(n_291), .B2(n_292), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_351), .A2(n_299), .B1(n_292), .B2(n_286), .Y(n_385) );
INVx8_ASAP7_75t_L g386 ( .A(n_320), .Y(n_386) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_382), .A2(n_344), .B1(n_337), .B2(n_319), .C(n_340), .Y(n_387) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_383), .A2(n_308), .B(n_286), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_364), .A2(n_349), .B(n_309), .Y(n_389) );
AOI33xp33_ASAP7_75t_L g390 ( .A1(n_384), .A2(n_292), .A3(n_344), .B1(n_299), .B2(n_290), .B3(n_331), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_380), .A2(n_310), .B1(n_309), .B2(n_312), .Y(n_391) );
CKINVDCx8_ASAP7_75t_R g392 ( .A(n_361), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_357), .B(n_309), .Y(n_393) );
OAI221xp5_ASAP7_75t_SL g394 ( .A1(n_362), .A2(n_290), .B1(n_350), .B2(n_308), .C(n_315), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_357), .B(n_306), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_317), .B1(n_306), .B2(n_310), .C(n_314), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_370), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_370), .A2(n_310), .B1(n_348), .B2(n_345), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_377), .A2(n_317), .B(n_348), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_307), .B(n_345), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_378), .A2(n_314), .B1(n_320), .B2(n_336), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_355), .A2(n_332), .B1(n_338), .B2(n_320), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_354), .A2(n_314), .B1(n_332), .B2(n_338), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_325), .B1(n_336), .B2(n_324), .C(n_323), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_330), .B1(n_305), .B2(n_303), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_378), .B(n_330), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g407 ( .A1(n_373), .A2(n_367), .B(n_385), .Y(n_407) );
AOI222xp33_ASAP7_75t_L g408 ( .A1(n_381), .A2(n_313), .B1(n_325), .B2(n_323), .C1(n_324), .C2(n_320), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_354), .A2(n_313), .B1(n_305), .B2(n_303), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_354), .A2(n_303), .B1(n_305), .B2(n_323), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_354), .A2(n_305), .B1(n_303), .B2(n_324), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_355), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_381), .A2(n_342), .B1(n_334), .B2(n_303), .C(n_305), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_413), .B(n_361), .Y(n_415) );
INVx4_ASAP7_75t_L g416 ( .A(n_397), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_411), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_411), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_395), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_397), .B(n_369), .Y(n_420) );
AOI33xp33_ASAP7_75t_L g421 ( .A1(n_387), .A2(n_366), .A3(n_376), .B1(n_372), .B2(n_365), .B3(n_374), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_395), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_407), .A2(n_365), .B1(n_370), .B2(n_369), .Y(n_423) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_413), .A2(n_370), .B1(n_363), .B2(n_379), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_365), .B1(n_369), .B2(n_363), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_406), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_393), .B(n_376), .Y(n_427) );
OAI21xp5_ASAP7_75t_L g428 ( .A1(n_389), .A2(n_365), .B(n_375), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_392), .A2(n_379), .B(n_386), .C(n_360), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_392), .A2(n_386), .B(n_360), .C(n_358), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_388), .A2(n_369), .B1(n_386), .B2(n_358), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_403), .B(n_375), .Y(n_433) );
OAI31xp33_ASAP7_75t_L g434 ( .A1(n_394), .A2(n_358), .A3(n_360), .B(n_335), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
NAND4xp25_ASAP7_75t_L g436 ( .A(n_390), .B(n_17), .C(n_229), .D(n_227), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_391), .A2(n_386), .B1(n_356), .B2(n_334), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_404), .A2(n_386), .B1(n_356), .B2(n_320), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_401), .A2(n_334), .B1(n_342), .B2(n_356), .C(n_330), .Y(n_440) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_399), .A2(n_342), .B1(n_356), .B2(n_330), .C(n_353), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_400), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_408), .A2(n_356), .B1(n_330), .B2(n_343), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_402), .A2(n_150), .B1(n_152), .B2(n_156), .C(n_234), .Y(n_444) );
OAI211xp5_ASAP7_75t_SL g445 ( .A1(n_410), .A2(n_193), .B(n_179), .C(n_229), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_412), .B(n_343), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_409), .A2(n_353), .B1(n_343), .B2(n_333), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_414), .Y(n_448) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_387), .A2(n_353), .B1(n_343), .B2(n_333), .C(n_322), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g450 ( .A(n_394), .B(n_353), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_436), .B(n_156), .C(n_152), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_419), .B(n_156), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_436), .A2(n_156), .B1(n_152), .B2(n_150), .C(n_279), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_422), .B(n_156), .Y(n_455) );
NAND4xp25_ASAP7_75t_SL g456 ( .A(n_429), .B(n_19), .C(n_20), .D(n_23), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_417), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_417), .Y(n_458) );
INVx5_ASAP7_75t_SL g459 ( .A(n_420), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
OR2x6_ASAP7_75t_L g461 ( .A(n_416), .B(n_353), .Y(n_461) );
OAI22xp33_ASAP7_75t_L g462 ( .A1(n_450), .A2(n_343), .B1(n_333), .B2(n_322), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_437), .A2(n_434), .B1(n_432), .B2(n_425), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_418), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_419), .B(n_152), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_422), .B(n_152), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_427), .B(n_333), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_418), .Y(n_468) );
INVx4_ASAP7_75t_L g469 ( .A(n_420), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_421), .B(n_200), .C(n_232), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_416), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g472 ( .A(n_434), .B(n_200), .C(n_232), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_422), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_420), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_427), .B(n_24), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_433), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_420), .B(n_27), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_433), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_415), .B(n_30), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_449), .A2(n_333), .B(n_322), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_442), .B(n_31), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
AND2x4_ASAP7_75t_L g485 ( .A(n_435), .B(n_32), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_435), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_423), .B(n_186), .C(n_232), .Y(n_487) );
NOR2xp33_ASAP7_75t_SL g488 ( .A(n_424), .B(n_322), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_439), .A2(n_322), .B1(n_179), .B2(n_227), .C(n_190), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_430), .B(n_34), .Y(n_490) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_441), .A2(n_190), .B(n_193), .Y(n_491) );
OAI33xp33_ASAP7_75t_L g492 ( .A1(n_448), .A2(n_206), .A3(n_209), .B1(n_279), .B2(n_278), .B3(n_296), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_448), .B(n_36), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_446), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_450), .B(n_39), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_440), .A2(n_431), .A3(n_438), .B(n_443), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_445), .A2(n_265), .B1(n_285), .B2(n_282), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
OAI322xp33_ASAP7_75t_L g501 ( .A1(n_437), .A2(n_206), .A3(n_209), .B1(n_228), .B2(n_232), .C1(n_181), .C2(n_200), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_451), .A2(n_296), .B(n_284), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_493), .B(n_41), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_457), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_493), .B(n_45), .Y(n_506) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_485), .A2(n_46), .A3(n_48), .B(n_56), .Y(n_507) );
AOI211x1_ASAP7_75t_L g508 ( .A1(n_477), .A2(n_57), .B(n_59), .C(n_61), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_481), .B(n_66), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_464), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_468), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_453), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_460), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_495), .B(n_67), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_471), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_474), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_495), .B(n_68), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_480), .B(n_70), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_486), .Y(n_521) );
NAND2x1p5_ASAP7_75t_L g522 ( .A(n_485), .B(n_285), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_486), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_454), .B(n_186), .C(n_232), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_476), .Y(n_526) );
BUFx4f_ASAP7_75t_SL g527 ( .A(n_469), .Y(n_527) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_485), .B(n_186), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_478), .B(n_73), .Y(n_529) );
AOI31xp33_ASAP7_75t_L g530 ( .A1(n_479), .A2(n_75), .A3(n_76), .B(n_263), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_473), .B(n_178), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_484), .B(n_178), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_469), .B(n_178), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_494), .A2(n_269), .B(n_284), .C(n_278), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_469), .B(n_178), .Y(n_535) );
INVx3_ASAP7_75t_L g536 ( .A(n_475), .Y(n_536) );
AND2x4_ASAP7_75t_SL g537 ( .A(n_479), .B(n_263), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_452), .B(n_178), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_467), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_452), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_465), .B(n_466), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_465), .B(n_181), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_466), .B(n_181), .Y(n_543) );
NOR3xp33_ASAP7_75t_SL g544 ( .A(n_456), .B(n_181), .C(n_186), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_475), .B(n_181), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_455), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_455), .Y(n_547) );
OAI31xp33_ASAP7_75t_L g548 ( .A1(n_472), .A2(n_269), .A3(n_234), .B(n_228), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_476), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_459), .B(n_186), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_497), .B(n_200), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_461), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_461), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_459), .B(n_200), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g555 ( .A(n_463), .B(n_228), .C(n_271), .D(n_273), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_461), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_459), .B(n_228), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_461), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_497), .B(n_228), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_488), .B(n_271), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_523), .B(n_459), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_513), .B(n_483), .Y(n_564) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_549), .B(n_498), .C(n_470), .D(n_490), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_511), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_512), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_514), .B(n_491), .Y(n_568) );
NAND4xp25_ASAP7_75t_L g569 ( .A(n_526), .B(n_496), .C(n_487), .D(n_483), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_539), .B(n_491), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_517), .B(n_500), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_516), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_523), .B(n_541), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_541), .B(n_496), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_521), .Y(n_576) );
CKINVDCx16_ASAP7_75t_R g577 ( .A(n_527), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_524), .Y(n_578) );
XOR2x2_ASAP7_75t_L g579 ( .A(n_528), .B(n_491), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_540), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_547), .B(n_482), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_540), .B(n_499), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_547), .B(n_462), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_537), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_546), .B(n_489), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_532), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g587 ( .A1(n_519), .A2(n_492), .B1(n_501), .B2(n_282), .C(n_285), .Y(n_587) );
OR2x6_ASAP7_75t_L g588 ( .A(n_528), .B(n_271), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_536), .B(n_556), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_552), .B(n_271), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_552), .B(n_273), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_551), .B(n_273), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_536), .B(n_273), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_551), .B(n_282), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_536), .B(n_282), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_532), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_529), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_530), .B(n_285), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_504), .A2(n_518), .B1(n_506), .B2(n_515), .C(n_559), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_529), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_537), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_520), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_551), .B(n_559), .Y(n_603) );
AOI21xp33_ASAP7_75t_SL g604 ( .A1(n_522), .A2(n_507), .B(n_510), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_559), .B(n_553), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_504), .B(n_506), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_520), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_515), .B(n_518), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_531), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_558), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_577), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_571), .B(n_522), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_572), .B(n_522), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_567), .B(n_555), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_569), .A2(n_525), .B1(n_535), .B2(n_557), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_579), .B(n_544), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_565), .A2(n_548), .B1(n_545), .B2(n_502), .C(n_535), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_573), .B(n_543), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_610), .B(n_533), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_574), .B(n_542), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_580), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_564), .A2(n_557), .B1(n_560), .B2(n_554), .C(n_550), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_604), .A2(n_534), .B(n_533), .C(n_538), .Y(n_623) );
INVx1_ASAP7_75t_SL g624 ( .A(n_584), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_574), .B(n_538), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
AND3x1_ASAP7_75t_L g627 ( .A(n_599), .B(n_550), .C(n_554), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_542), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_562), .B(n_508), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_566), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_563), .B(n_533), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_581), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_589), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_575), .Y(n_634) );
INVx1_ASAP7_75t_SL g635 ( .A(n_601), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_578), .B(n_597), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_568), .Y(n_638) );
INVx3_ASAP7_75t_L g639 ( .A(n_579), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_600), .B(n_602), .Y(n_640) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_586), .Y(n_641) );
OAI21xp33_ASAP7_75t_L g642 ( .A1(n_605), .A2(n_568), .B(n_581), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_603), .B(n_605), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_607), .A2(n_609), .B1(n_606), .B2(n_608), .C1(n_603), .C2(n_582), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_606), .A2(n_585), .B1(n_582), .B2(n_598), .C(n_570), .Y(n_645) );
INVx8_ASAP7_75t_L g646 ( .A(n_588), .Y(n_646) );
CKINVDCx6p67_ASAP7_75t_R g647 ( .A(n_588), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_570), .B(n_585), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_587), .B(n_598), .Y(n_649) );
AOI21xp5_ASAP7_75t_SL g650 ( .A1(n_588), .A2(n_583), .B(n_561), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_561), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_588), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_593), .A2(n_595), .B(n_592), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_590), .Y(n_655) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_594), .B(n_592), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_591), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_594), .A2(n_577), .B1(n_527), .B2(n_549), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_591), .Y(n_659) );
AOI21xp33_ASAP7_75t_SL g660 ( .A1(n_577), .A2(n_530), .B(n_598), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_571), .B(n_572), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_577), .A2(n_527), .B1(n_549), .B2(n_599), .Y(n_662) );
AOI221x1_ASAP7_75t_L g663 ( .A1(n_660), .A2(n_639), .B1(n_662), .B2(n_650), .C(n_658), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_616), .A2(n_649), .B(n_646), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_639), .A2(n_611), .B(n_645), .C(n_646), .Y(n_665) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_639), .A2(n_635), .B1(n_624), .B2(n_661), .Y(n_666) );
OAI211xp5_ASAP7_75t_L g667 ( .A1(n_645), .A2(n_649), .B(n_623), .C(n_644), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_648), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_646), .A2(n_627), .B(n_615), .Y(n_669) );
O2A1O1Ixp33_ASAP7_75t_L g670 ( .A1(n_629), .A2(n_614), .B(n_617), .C(n_633), .Y(n_670) );
NAND4xp75_ASAP7_75t_L g671 ( .A(n_619), .B(n_653), .C(n_612), .D(n_613), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_636), .Y(n_672) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_653), .A2(n_642), .B(n_622), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_640), .A2(n_656), .B1(n_638), .B2(n_632), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_647), .A2(n_655), .B1(n_643), .B2(n_651), .Y(n_675) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_652), .B(n_638), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_667), .A2(n_637), .B1(n_632), .B2(n_655), .C(n_636), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_672), .Y(n_678) );
O2A1O1Ixp5_ASAP7_75t_L g679 ( .A1(n_664), .A2(n_631), .B(n_634), .C(n_626), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_670), .B(n_625), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_665), .A2(n_659), .B1(n_654), .B2(n_657), .C(n_634), .Y(n_681) );
INVx2_ASAP7_75t_SL g682 ( .A(n_666), .Y(n_682) );
NOR3xp33_ASAP7_75t_SL g683 ( .A(n_669), .B(n_628), .C(n_630), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_673), .A2(n_625), .B(n_620), .C(n_618), .Y(n_684) );
NAND2xp33_ASAP7_75t_L g685 ( .A(n_683), .B(n_671), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_677), .A2(n_673), .B1(n_675), .B2(n_668), .C(n_674), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_678), .Y(n_687) );
NOR4xp75_ASAP7_75t_L g688 ( .A(n_682), .B(n_663), .C(n_620), .D(n_618), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_687), .Y(n_689) );
OR3x1_ASAP7_75t_L g690 ( .A(n_688), .B(n_684), .C(n_679), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_685), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_689), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_691), .A2(n_686), .B1(n_681), .B2(n_680), .C(n_676), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_692), .Y(n_694) );
NOR3x1_ASAP7_75t_L g695 ( .A(n_693), .B(n_691), .C(n_690), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_694), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_696), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_695), .B1(n_641), .B2(n_626), .C(n_621), .Y(n_698) );
endmodule