module fake_jpeg_2663_n_76 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_31;
wire n_17;
wire n_25;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx6p67_ASAP7_75t_R g25 ( 
.A(n_19),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_10),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_23),
.B1(n_11),
.B2(n_8),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_32),
.B1(n_19),
.B2(n_21),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_20),
.A2(n_12),
.B1(n_17),
.B2(n_11),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_25),
.B1(n_26),
.B2(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

OAI22x1_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_23),
.B1(n_11),
.B2(n_9),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_27),
.B1(n_34),
.B2(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_46),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_34),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_47),
.C(n_48),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_44),
.C(n_34),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_40),
.C(n_53),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_47),
.B(n_25),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_26),
.C(n_4),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_25),
.B(n_38),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_51),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_58),
.B(n_26),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_62),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_4),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_56),
.B(n_6),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_73),
.Y(n_76)
);


endmodule