module real_jpeg_25125_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_348, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_348;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_1),
.A2(n_27),
.B1(n_29),
.B2(n_59),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_125),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_2),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_57),
.B1(n_75),
.B2(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_125),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_125),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_5),
.B(n_68),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_5),
.B(n_47),
.C(n_50),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_130),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_30),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_106),
.B1(n_210),
.B2(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_6),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_7),
.A2(n_70),
.B1(n_71),
.B2(n_74),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_7),
.A2(n_50),
.B1(n_51),
.B2(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_70),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_34),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_8),
.A2(n_26),
.B1(n_58),
.B2(n_74),
.Y(n_296)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_10),
.A2(n_42),
.B1(n_75),
.B2(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_119)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_11),
.B(n_29),
.C(n_64),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_12),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_127),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_127),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_12),
.A2(n_58),
.B1(n_66),
.B2(n_127),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_13),
.A2(n_58),
.B1(n_66),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_13),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_27),
.B1(n_29),
.B2(n_133),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_133),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_133),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_15),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_97),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_76),
.C(n_80),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_20),
.A2(n_76),
.B1(n_331),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_20),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_22),
.B(n_44),
.C(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_24),
.A2(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_25),
.A2(n_30),
.B(n_38),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_25),
.A2(n_38),
.B(n_83),
.Y(n_276)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_29),
.B1(n_32),
.B2(n_36),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_27),
.A2(n_29),
.B1(n_62),
.B2(n_64),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_27),
.A2(n_62),
.B(n_129),
.C(n_154),
.Y(n_153)
);

HAxp5_ASAP7_75t_SL g227 ( 
.A(n_27),
.B(n_130),
.CON(n_227),
.SN(n_227)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_29),
.B(n_32),
.C(n_34),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_30),
.A2(n_38),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_30),
.A2(n_38),
.B1(n_170),
.B2(n_227),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_30),
.A2(n_38),
.B1(n_82),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_31),
.B(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_31),
.A2(n_143),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_31),
.A2(n_37),
.B(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_31)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_33),
.A2(n_36),
.B(n_226),
.C(n_228),
.Y(n_225)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_34),
.B(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_38),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_38),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_76),
.C(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_43),
.A2(n_44),
.B1(n_81),
.B2(n_334),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_45),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_45),
.A2(n_49),
.B1(n_185),
.B2(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_45),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_45),
.A2(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_49),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_49),
.B(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_49),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_49),
.B(n_130),
.Y(n_208)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_51),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_51),
.B(n_216),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_117),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_53),
.B(n_183),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_61),
.B(n_77),
.Y(n_76)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_69),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_60),
.A2(n_68),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_60),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_60),
.A2(n_68),
.B1(n_140),
.B2(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_132),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_68),
.B(n_296),
.Y(n_295)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_75),
.B(n_130),
.CON(n_129),
.SN(n_129)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_76),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_76),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_80),
.B(n_338),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_81),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_93),
.B2(n_94),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_90),
.A2(n_138),
.B(n_320),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_328),
.A3(n_340),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_305),
.B(n_327),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_279),
.B(n_304),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_172),
.B(n_260),
.C(n_278),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_156),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_102),
.B(n_156),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_134),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_120),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_104),
.B(n_120),
.C(n_134),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_105),
.B(n_114),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_110),
.B(n_112),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_106),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_106),
.A2(n_203),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_106),
.A2(n_112),
.B(n_192),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_106),
.A2(n_192),
.B(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_111),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_107),
.B(n_113),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_107),
.A2(n_164),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_108),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_108),
.Y(n_211)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_115),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_116),
.B(n_250),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_117),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_117),
.A2(n_183),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_117),
.A2(n_183),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.C(n_128),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_123),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_122),
.Y(n_288)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_130),
.B(n_217),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_144),
.B2(n_155),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_137),
.B(n_141),
.C(n_155),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_138),
.A2(n_294),
.B(n_295),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_146),
.B1(n_153),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_152),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_157),
.B(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_159),
.B(n_161),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_162),
.A2(n_166),
.B1(n_167),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_165),
.B(n_189),
.Y(n_266)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_259),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_254),
.B(n_258),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_238),
.B(n_253),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_221),
.B(n_237),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_199),
.B(n_220),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_186),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_181),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_194),
.C(n_197),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_198),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_219),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_205),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_218),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_236),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_231),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_232),
.C(n_233),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_229),
.B2(n_230),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_240),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_248),
.C(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_277),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_271),
.C(n_277),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_270),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_270),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_269),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_274),
.C(n_276),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_275),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_281),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_303),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_290),
.B1(n_301),
.B2(n_302),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_302),
.C(n_303),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_289),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_284),
.A2(n_285),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_284),
.A2(n_315),
.B(n_319),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_285),
.B(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_290),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_297),
.C(n_300),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_292)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_296),
.Y(n_320)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_299),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_306),
.B(n_307),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_308),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_307)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_314),
.B1(n_322),
.B2(n_323),
.Y(n_308)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_310),
.B(n_312),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_313),
.A2(n_330),
.B1(n_335),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_322),
.C(n_326),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_321),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_324),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_337),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_337),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.C(n_336),
.Y(n_329)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);


endmodule