module real_jpeg_154_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_0),
.A2(n_54),
.B1(n_62),
.B2(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_46),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_2),
.A2(n_46),
.B1(n_62),
.B2(n_66),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_3),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_86),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_86),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_62),
.B1(n_66),
.B2(n_86),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_5),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_148),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_148),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_5),
.A2(n_62),
.B1(n_66),
.B2(n_148),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_6),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_126),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_6),
.A2(n_62),
.B1(n_66),
.B2(n_126),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_8),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_180),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_180),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_8),
.A2(n_62),
.B1(n_66),
.B2(n_180),
.Y(n_290)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_12),
.A2(n_42),
.B1(n_43),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_12),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_78),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_12),
.A2(n_62),
.B1(n_66),
.B2(n_78),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_38),
.B1(n_62),
.B2(n_66),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_15),
.B(n_42),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_15),
.B(n_55),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_15),
.A2(n_25),
.B(n_26),
.C(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_15),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_15),
.B(n_31),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_15),
.A2(n_26),
.B1(n_27),
.B2(n_230),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_15),
.B(n_62),
.C(n_65),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_230),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_15),
.B(n_116),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_15),
.B(n_60),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_91),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_79),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_79),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_58),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_39),
.B1(n_56),
.B2(n_57),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_24),
.B(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_24),
.A2(n_31),
.B1(n_197),
.B2(n_214),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_30),
.C(n_31),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_26),
.Y(n_30)
);

AO22x2_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_27),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_26),
.A2(n_43),
.A3(n_49),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g202 ( 
.A(n_27),
.B(n_51),
.Y(n_202)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_31),
.B(n_177),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_32),
.A2(n_33),
.B1(n_64),
.B2(n_65),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_32),
.A2(n_35),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_33),
.B(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_37),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_48),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

O2A1O1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_43),
.A2(n_76),
.B(n_230),
.C(n_239),
.Y(n_238)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_47),
.B(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_47),
.A2(n_55),
.B1(n_147),
.B2(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_76),
.B1(n_77),
.B2(n_85),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_48),
.A2(n_85),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_48),
.B(n_125),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_48),
.A2(n_123),
.B(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_71),
.C(n_75),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_59),
.A2(n_71),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_59),
.B(n_84),
.C(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_59),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_67),
.B(n_69),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_60),
.A2(n_67),
.B1(n_121),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_60),
.A2(n_67),
.B1(n_142),
.B2(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_60),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_70),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_61),
.A2(n_102),
.B1(n_103),
.B2(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_61),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_61),
.A2(n_246),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_61),
.A2(n_102),
.B1(n_223),
.B2(n_257),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_61)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_62),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_62),
.B(n_286),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_67),
.A2(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_67),
.B(n_226),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_74),
.B1(n_90),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_72),
.A2(n_74),
.B1(n_100),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_72),
.A2(n_196),
.B(n_198),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_72),
.A2(n_198),
.B(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_74),
.A2(n_144),
.B(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_74),
.A2(n_176),
.B(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_76),
.A2(n_146),
.B(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_87),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_80),
.A2(n_84),
.B1(n_105),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_80),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_156),
.B(n_327),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_151),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_127),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_96),
.B(n_127),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_108),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_99),
.B(n_101),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_104),
.C(n_108),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_102),
.A2(n_225),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_122),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_110),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_111),
.A2(n_112),
.B1(n_122),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_111),
.A2(n_112),
.B1(n_119),
.B2(n_166),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_116),
.B(n_117),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_113),
.A2(n_116),
.B1(n_139),
.B2(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_113),
.A2(n_230),
.B(n_263),
.Y(n_287)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_114),
.A2(n_115),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_114),
.A2(n_115),
.B1(n_205),
.B2(n_220),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_114),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_114),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_114),
.A2(n_115),
.B1(n_261),
.B2(n_295),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_115),
.A2(n_220),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_115),
.B(n_234),
.Y(n_263)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_116),
.A2(n_233),
.B(n_290),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.C(n_134),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_129),
.B1(n_133),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_143),
.C(n_145),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_135),
.A2(n_136),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_137),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_145),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_150),
.B(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_151),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_152),
.B(n_155),
.Y(n_329)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_181),
.B(n_326),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_158),
.B(n_161),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.C(n_167),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_165),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.C(n_178),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_169),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_170),
.B(n_172),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_171),
.Y(n_245)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_207),
.B(n_325),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_183),
.B(n_185),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.C(n_192),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_186),
.B(n_190),
.Y(n_310)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_192),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_199),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_193),
.B(n_195),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_199),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_200),
.A2(n_203),
.B1(n_204),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AOI31xp33_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_307),
.A3(n_317),
.B(n_322),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_251),
.B(n_306),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_235),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_210),
.B(n_235),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_221),
.C(n_227),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_216),
.C(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_221),
.B(n_227),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_231),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_247),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_236),
.B(n_248),
.C(n_250),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_237),
.B(n_242),
.C(n_243),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_301),
.B(n_305),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_270),
.B(n_300),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_264),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_264),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_260),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_282),
.B(n_299),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_278),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_278),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_273),
.A2(n_274),
.B1(n_276),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_279),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_293),
.B(n_298),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_288),
.B(n_292),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_291),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_290),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_296),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_309),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.C(n_315),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_319),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_314),
.Y(n_320)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_321),
.Y(n_323)
);


endmodule