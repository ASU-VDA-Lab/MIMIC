module fake_jpeg_12283_n_237 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_0),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_58),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_63),
.Y(n_76)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_24),
.B(n_1),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_25),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_37),
.B(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_15),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_80),
.B1(n_87),
.B2(n_61),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_39),
.B1(n_33),
.B2(n_29),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_93),
.B1(n_94),
.B2(n_47),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_39),
.B1(n_62),
.B2(n_48),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_70),
.A2(n_18),
.A3(n_63),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_37),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_78),
.B(n_79),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_30),
.B1(n_17),
.B2(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_38),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_92),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_30),
.B1(n_33),
.B2(n_20),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_57),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_20),
.B1(n_25),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_42),
.A2(n_35),
.B1(n_19),
.B2(n_32),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_45),
.B(n_34),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_18),
.Y(n_117)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_102),
.Y(n_129)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_19),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_111),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_34),
.B1(n_23),
.B2(n_32),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_119),
.B1(n_123),
.B2(n_11),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_110),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_26),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_71),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_69),
.C(n_68),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g150 ( 
.A(n_115),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_26),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_84),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_67),
.A2(n_70),
.B1(n_80),
.B2(n_87),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_23),
.B1(n_54),
.B2(n_57),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_121),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_18),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_71),
.A2(n_89),
.B(n_18),
.C(n_16),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_124),
.B(n_1),
.C(n_6),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_13),
.B(n_2),
.C(n_6),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_73),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_8),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_86),
.B(n_84),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_140),
.C(n_126),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_107),
.B(n_105),
.C(n_103),
.D(n_115),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_72),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_145),
.Y(n_160)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_69),
.A3(n_68),
.B1(n_83),
.B2(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_132),
.Y(n_166)
);

AOI22x1_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_83),
.B1(n_84),
.B2(n_9),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_114),
.B1(n_108),
.B2(n_141),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_106),
.B1(n_99),
.B2(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_102),
.B(n_6),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_166),
.B1(n_139),
.B2(n_138),
.C(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_123),
.B1(n_112),
.B2(n_113),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_161),
.B1(n_168),
.B2(n_171),
.Y(n_188)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_143),
.A2(n_127),
.B1(n_112),
.B2(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_169),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_116),
.C(n_98),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_165),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_100),
.C(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_172),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_104),
.B1(n_103),
.B2(n_10),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_8),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_11),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_173),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_154),
.B(n_129),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_177),
.B(n_138),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_135),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_190),
.C(n_160),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_183),
.B(n_186),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_128),
.B(n_144),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_167),
.B(n_154),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_131),
.B(n_144),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_189),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_196),
.Y(n_206)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_198),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_176),
.A2(n_161),
.B1(n_142),
.B2(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_172),
.B1(n_137),
.B2(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_201),
.Y(n_211)
);

OAI322xp33_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_151),
.A3(n_170),
.B1(n_173),
.B2(n_157),
.C1(n_171),
.C2(n_168),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_159),
.B1(n_152),
.B2(n_136),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_148),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_147),
.C(n_148),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_147),
.C(n_150),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_182),
.C(n_179),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_190),
.C(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_187),
.C(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_178),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_211),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_197),
.B(n_203),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_217),
.B(n_219),
.C(n_220),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_204),
.B(n_202),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_188),
.C(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_211),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_224),
.B(n_226),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_213),
.C(n_195),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_215),
.A2(n_199),
.B1(n_175),
.B2(n_146),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_146),
.C(n_225),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_222),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_225),
.A2(n_223),
.B1(n_221),
.B2(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_232),
.Y(n_235)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_233),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g237 ( 
.A(n_236),
.B(n_234),
.CI(n_231),
.CON(n_237),
.SN(n_237)
);


endmodule