module real_jpeg_33598_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_0),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_0),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g387 ( 
.A(n_0),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_1),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_1),
.A2(n_86),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g183 ( 
.A1(n_1),
.A2(n_86),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_1),
.A2(n_39),
.B1(n_86),
.B2(n_260),
.Y(n_259)
);

CKINVDCx11_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_2),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_2),
.B(n_485),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_4),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_5),
.Y(n_199)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_6),
.A2(n_51),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_6),
.A2(n_51),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_6),
.A2(n_51),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_6),
.B(n_310),
.Y(n_309)
);

OAI32xp33_ASAP7_75t_L g325 ( 
.A1(n_6),
.A2(n_326),
.A3(n_328),
.B1(n_330),
.B2(n_336),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_6),
.B(n_97),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_6),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_6),
.B(n_163),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_7),
.Y(n_341)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

AOI221xp5_ASAP7_75t_L g14 ( 
.A1(n_10),
.A2(n_15),
.B1(n_16),
.B2(n_468),
.C(n_483),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_11),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_111),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_11),
.A2(n_111),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_11),
.A2(n_111),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_12),
.Y(n_142)
);

AOI22x1_ASAP7_75t_L g38 ( 
.A1(n_13),
.A2(n_39),
.B1(n_42),
.B2(n_46),
.Y(n_38)
);

INVx2_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_13),
.A2(n_46),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_13),
.A2(n_46),
.B1(n_291),
.B2(n_293),
.Y(n_290)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_262),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_239),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_206),
.Y(n_20)
);

OAI21x1_ASAP7_75t_SL g478 ( 
.A1(n_21),
.A2(n_479),
.B(n_480),
.Y(n_478)
);

NOR2x1_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_148),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_22),
.B(n_148),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_129),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_23),
.B(n_24),
.C(n_130),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.C(n_94),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_24),
.A2(n_25),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_25),
.B(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_26),
.Y(n_273)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_27),
.B(n_213),
.C(n_270),
.Y(n_432)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g424 ( 
.A1(n_28),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_28),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_38),
.B(n_47),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_29),
.A2(n_38),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_29),
.B(n_135),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_SL g246 ( 
.A1(n_29),
.A2(n_247),
.B(n_253),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_29),
.A2(n_135),
.B1(n_247),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_55),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_30),
.Y(n_310)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_35),
.Y(n_283)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_41),
.Y(n_252)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_46),
.A2(n_145),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_46),
.B(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_47),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.Y(n_47)
);

INVxp33_ASAP7_75t_SL g136 ( 
.A(n_48),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_48),
.B(n_205),
.Y(n_204)
);

OAI21x1_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_51),
.B(n_52),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_51),
.B(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_51),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_51),
.B(n_374),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g276 ( 
.A1(n_52),
.A2(n_248),
.A3(n_277),
.B1(n_281),
.B2(n_284),
.Y(n_276)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

AOI22x1_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_59),
.Y(n_286)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_62),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_63),
.A2(n_64),
.B1(n_94),
.B2(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_64),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_64),
.B(n_132),
.C(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_85),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_65),
.B(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_77),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_77),
.Y(n_66)
);

NAND2x1p5_ASAP7_75t_L g162 ( 
.A(n_67),
.B(n_77),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_75),
.Y(n_67)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_68),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_69),
.Y(n_157)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_69),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_69),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_69),
.Y(n_377)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_72),
.Y(n_372)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_76),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_77),
.B(n_229),
.Y(n_350)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_79),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_82),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_83),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_85),
.A2(n_155),
.B1(n_161),
.B2(n_163),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_88),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22x1_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_99),
.B1(n_102),
.B2(n_106),
.Y(n_98)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_92),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_93),
.Y(n_180)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_108),
.B(n_115),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_96),
.A2(n_108),
.B1(n_139),
.B2(n_147),
.Y(n_138)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_R g245 ( 
.A(n_96),
.B(n_147),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_96),
.A2(n_147),
.B(n_165),
.Y(n_426)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_97),
.B(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_116),
.B(n_120),
.Y(n_215)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_119),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_120),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_127),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_126),
.Y(n_335)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_128),
.Y(n_288)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_132),
.B(n_213),
.C(n_216),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_132),
.B(n_164),
.C(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g430 ( 
.A1(n_133),
.A2(n_134),
.B1(n_164),
.B2(n_307),
.Y(n_430)
);

AOI22x1_ASAP7_75t_L g449 ( 
.A1(n_133),
.A2(n_134),
.B1(n_213),
.B2(n_271),
.Y(n_449)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_138),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_139),
.Y(n_244)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g280 ( 
.A(n_142),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_142),
.Y(n_327)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_171),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OA21x2_ASAP7_75t_L g234 ( 
.A1(n_153),
.A2(n_154),
.B(n_164),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_164),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_163),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AO22x2_ASAP7_75t_L g226 ( 
.A1(n_161),
.A2(n_163),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_164),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_164),
.A2(n_307),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_208),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_182),
.B(n_203),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_172),
.B(n_237),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_181),
.B(n_182),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_173),
.B(n_181),
.Y(n_446)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_175),
.B(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_176),
.Y(n_227)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_182),
.A2(n_203),
.B1(n_204),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_182),
.A2(n_238),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_190),
.Y(n_292)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_190),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_191),
.B(n_299),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_200),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_218),
.B1(n_219),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_193),
.A2(n_290),
.B1(n_296),
.B2(n_299),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_193),
.B(n_299),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_197),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_199),
.Y(n_380)
);

INVx3_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g475 ( 
.A(n_205),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_207),
.B(n_210),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_234),
.C(n_235),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_212),
.B(n_234),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_213),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_269)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_213),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_213),
.A2(n_271),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_216),
.B(n_449),
.Y(n_448)
);

NAND2x1_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.Y(n_216)
);

OAI22x1_ASAP7_75t_L g417 ( 
.A1(n_217),
.A2(n_323),
.B1(n_402),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_217),
.Y(n_418)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_220),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_221),
.A2(n_316),
.B(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_226),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_226),
.B(n_354),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_226),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_236),
.B(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_256),
.Y(n_239)
);

A2O1A1O1Ixp25_ASAP7_75t_L g477 ( 
.A1(n_240),
.A2(n_256),
.B(n_478),
.C(n_481),
.D(n_482),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_241),
.B(n_242),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_242),
.Y(n_490)
);

FAx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.CI(n_254),
.CON(n_242),
.SN(n_242)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_246),
.C(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx11_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_257),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_R g482 ( 
.A(n_257),
.B(n_261),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_257),
.B(n_488),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2x1_ASAP7_75t_L g474 ( 
.A(n_259),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_460),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_409),
.B(n_459),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_343),
.B(n_408),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_317),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_267),
.B(n_317),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_268),
.B(n_275),
.C(n_306),
.Y(n_434)
);

XNOR2x1_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_270),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_271),
.B(n_396),
.C(n_406),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_273),
.B(n_441),
.C(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_273),
.B(n_441),
.C(n_442),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_306),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_289),
.B1(n_304),
.B2(n_305),
.Y(n_275)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_276),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_276),
.B(n_305),
.Y(n_415)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_289),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_289),
.B(n_389),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_289),
.B(n_389),
.Y(n_390)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx4f_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_305),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.C(n_311),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_309),
.B1(n_311),
.B2(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_311),
.B(n_358),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_SL g391 ( 
.A(n_311),
.B(n_358),
.Y(n_391)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_312),
.B(n_383),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_315),
.B(n_316),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_322),
.C(n_324),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_318),
.A2(n_319),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_353),
.C(n_354),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_323),
.A2(n_324),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_324),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_342),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_325),
.B(n_342),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx4f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_399),
.B(n_407),
.Y(n_343)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_355),
.B(n_398),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_352),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_346),
.B(n_352),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_347),
.Y(n_406)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_349),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_349),
.B(n_359),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_349),
.B(n_421),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_349),
.B(n_421),
.Y(n_431)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_356),
.A2(n_392),
.B(n_397),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_381),
.B(n_391),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_360),
.A2(n_365),
.B1(n_373),
.B2(n_378),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_369),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_378),
.B(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_388),
.B(n_390),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx4_ASAP7_75t_SL g386 ( 
.A(n_387),
.Y(n_386)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_393),
.B(n_395),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_405),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_405),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_401),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_437),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_433),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_411),
.B(n_464),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_428),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_412),
.B(n_428),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_416),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_413),
.B(n_457),
.C(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_417),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

XNOR2x1_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_424),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_426),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_431),
.C(n_432),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_429),
.B(n_436),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_432),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_435),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_452),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_450),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_450),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_443),
.C(n_447),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_448),
.Y(n_455)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_456),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_467),
.Y(n_460)
);

A2O1A1Ixp33_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_463),
.B(n_465),
.C(n_466),
.Y(n_461)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_477),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_474),
.Y(n_488)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_486),
.Y(n_485)
);


endmodule