module fake_jpeg_7061_n_12 (n_3, n_2, n_1, n_0, n_4, n_12);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_12;

wire n_11;
wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

AOI22xp33_ASAP7_75t_SL g5 ( 
.A1(n_2),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_5)
);

INVx1_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

OAI32xp33_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVxp33_ASAP7_75t_SL g9 ( 
.A(n_7),
.Y(n_9)
);

AOI322xp5_ASAP7_75t_L g11 ( 
.A1(n_10),
.A2(n_9),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_0),
.C2(n_3),
.Y(n_11)
);

OAI321xp33_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_10),
.A3(n_7),
.B1(n_4),
.B2(n_2),
.C(n_1),
.Y(n_12)
);


endmodule