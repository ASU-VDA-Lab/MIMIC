module fake_jpeg_13316_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx8_ASAP7_75t_SL g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_60),
.Y(n_109)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_52),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_53),
.B(n_59),
.Y(n_101)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_62),
.B(n_66),
.Y(n_118)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_0),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_72),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_83),
.Y(n_120)
);

INVx2_ASAP7_75t_R g70 ( 
.A(n_43),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_30),
.B(n_1),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_78),
.Y(n_148)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

CKINVDCx6p67_ASAP7_75t_R g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_82),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_22),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_87),
.Y(n_137)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_22),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_32),
.B(n_4),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_90),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_35),
.B(n_5),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_18),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_91),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_45),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_18),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_95),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_26),
.B1(n_44),
.B2(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_102),
.A2(n_104),
.B1(n_112),
.B2(n_121),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_48),
.A2(n_45),
.B1(n_40),
.B2(n_46),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_115),
.B(n_34),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g160 ( 
.A(n_119),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_50),
.A2(n_45),
.B1(n_40),
.B2(n_46),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_70),
.A2(n_20),
.B1(n_42),
.B2(n_28),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_93),
.B1(n_61),
.B2(n_19),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_84),
.A2(n_52),
.B1(n_80),
.B2(n_56),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_143),
.B1(n_147),
.B2(n_17),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_72),
.A2(n_39),
.B(n_38),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_33),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_54),
.A2(n_65),
.B1(n_67),
.B2(n_71),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_58),
.B1(n_47),
.B2(n_78),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_51),
.A2(n_44),
.B1(n_26),
.B2(n_20),
.Y(n_143)
);

HAxp5_ASAP7_75t_SL g144 ( 
.A(n_63),
.B(n_20),
.CON(n_144),
.SN(n_144)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_128),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_94),
.A2(n_44),
.B1(n_26),
.B2(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_135),
.B(n_137),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_149),
.B(n_127),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_77),
.B1(n_42),
.B2(n_28),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_150),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_108),
.B(n_68),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_179),
.Y(n_193)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_42),
.B1(n_28),
.B2(n_23),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_161),
.B1(n_177),
.B2(n_178),
.Y(n_208)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_23),
.B1(n_19),
.B2(n_17),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_166),
.B(n_173),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_57),
.B1(n_55),
.B2(n_82),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_167),
.B1(n_172),
.B2(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_89),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_168),
.B(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_171),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_101),
.A2(n_64),
.B1(n_39),
.B2(n_38),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_128),
.A2(n_17),
.B1(n_19),
.B2(n_15),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_117),
.A2(n_15),
.B1(n_34),
.B2(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_96),
.B(n_15),
.Y(n_179)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_98),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

INVx11_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_104),
.A2(n_121),
.B1(n_147),
.B2(n_143),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_182),
.A2(n_189),
.B1(n_111),
.B2(n_103),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_83),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_186),
.C(n_124),
.Y(n_211)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_185),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_83),
.Y(n_186)
);

NOR2xp67_ASAP7_75t_SL g205 ( 
.A(n_187),
.B(n_116),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_118),
.B(n_32),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_191),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_92),
.B1(n_81),
.B2(n_8),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_109),
.A2(n_81),
.B1(n_6),
.B2(n_8),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_100),
.B1(n_131),
.B2(n_106),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_126),
.B(n_5),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_120),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_212),
.C(n_222),
.Y(n_237)
);

FAx1_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_144),
.CI(n_116),
.CON(n_201),
.SN(n_201)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_201),
.B(n_205),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_162),
.A2(n_99),
.B(n_107),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_211),
.Y(n_247)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_162),
.B(n_132),
.C(n_142),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_165),
.A2(n_117),
.B1(n_129),
.B2(n_148),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_213),
.A2(n_170),
.B1(n_152),
.B2(n_171),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_224),
.B1(n_189),
.B2(n_167),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_188),
.B(n_127),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_201),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_187),
.A2(n_145),
.B(n_131),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_181),
.B(n_176),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_166),
.B(n_5),
.Y(n_222)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_224),
.A2(n_182),
.B1(n_160),
.B2(n_157),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_229),
.A2(n_234),
.B1(n_238),
.B2(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_230),
.Y(n_273)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_207),
.Y(n_231)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_231),
.Y(n_278)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_236),
.Y(n_255)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_235),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_169),
.B1(n_173),
.B2(n_160),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_193),
.B(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_199),
.A2(n_173),
.B1(n_160),
.B2(n_164),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_158),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_242),
.Y(n_268)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_249),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_159),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_197),
.A2(n_198),
.B1(n_206),
.B2(n_217),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_166),
.B1(n_186),
.B2(n_183),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_244),
.A2(n_246),
.B1(n_155),
.B2(n_217),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_197),
.A2(n_186),
.B1(n_183),
.B2(n_111),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_248),
.A2(n_184),
.B(n_153),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_175),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_211),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_214),
.B(n_151),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_221),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_203),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_261),
.C(n_262),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_258),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_225),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_275),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_222),
.C(n_220),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_216),
.C(n_196),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_201),
.B(n_208),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_264),
.A2(n_276),
.B(n_240),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_218),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_218),
.C(n_223),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_238),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g274 ( 
.A1(n_234),
.A2(n_223),
.B(n_204),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_246),
.B(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_180),
.C(n_204),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_253),
.A2(n_202),
.B(n_163),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_248),
.B(n_250),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_241),
.B1(n_239),
.B2(n_249),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_282),
.A2(n_297),
.B1(n_267),
.B2(n_260),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_283),
.A2(n_284),
.B(n_291),
.Y(n_308)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_292),
.Y(n_317)
);

AO21x1_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_274),
.B(n_267),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_251),
.B1(n_244),
.B2(n_228),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_296),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_5),
.C(n_6),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_278),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_271),
.A2(n_227),
.B1(n_240),
.B2(n_233),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_277),
.B(n_233),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_299),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_202),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_301),
.B(n_263),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_274),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_303),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_305),
.B(n_311),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_257),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_309),
.B(n_315),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_310),
.A2(n_274),
.B1(n_294),
.B2(n_297),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_265),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_258),
.C(n_262),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_312),
.B(n_319),
.C(n_276),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_313),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_285),
.B(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_256),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_293),
.B(n_261),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_268),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_255),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_268),
.C(n_255),
.Y(n_319)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_317),
.A2(n_288),
.B1(n_299),
.B2(n_303),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_337),
.Y(n_343)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_332),
.C(n_279),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_282),
.Y(n_332)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_283),
.CI(n_291),
.CON(n_334),
.SN(n_334)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_334),
.B(n_340),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_336),
.A2(n_320),
.B1(n_322),
.B2(n_321),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_317),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_340),
.C(n_308),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_316),
.B(n_284),
.C(n_269),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_342),
.A2(n_351),
.B1(n_341),
.B2(n_327),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_329),
.B(n_315),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_349),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_309),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_355),
.C(n_333),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_348),
.B(n_331),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_325),
.A2(n_308),
.B(n_324),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_326),
.B(n_307),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_350),
.B(n_346),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_336),
.A2(n_304),
.B1(n_320),
.B2(n_307),
.Y(n_351)
);

NOR3xp33_ASAP7_75t_SL g353 ( 
.A(n_335),
.B(n_304),
.C(n_323),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_353),
.A2(n_296),
.B1(n_290),
.B2(n_287),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_323),
.B(n_302),
.Y(n_354)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_354),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_356),
.A2(n_359),
.B(n_366),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_338),
.C(n_332),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_365),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_358),
.A2(n_343),
.B1(n_344),
.B2(n_354),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_348),
.A2(n_334),
.B(n_339),
.Y(n_359)
);

OAI21x1_ASAP7_75t_L g375 ( 
.A1(n_361),
.A2(n_364),
.B(n_334),
.Y(n_375)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_352),
.Y(n_362)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_362),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_352),
.A2(n_329),
.B(n_328),
.Y(n_364)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_363),
.B(n_343),
.Y(n_369)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_355),
.C(n_354),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_370),
.B(n_374),
.C(n_113),
.Y(n_378)
);

BUFx24_ASAP7_75t_SL g373 ( 
.A(n_359),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_373),
.A2(n_375),
.B1(n_358),
.B2(n_360),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_351),
.C(n_344),
.Y(n_374)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_372),
.A2(n_353),
.B1(n_286),
.B2(n_221),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_379),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_9),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_374),
.A2(n_103),
.B1(n_113),
.B2(n_146),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_146),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_380),
.A2(n_371),
.B(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_384),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_386),
.A2(n_387),
.B(n_380),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_377),
.B(n_9),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_388),
.A2(n_383),
.B(n_11),
.Y(n_392)
);

MAJx2_ASAP7_75t_L g389 ( 
.A(n_385),
.B(n_378),
.C(n_381),
.Y(n_389)
);

AOI21xp33_ASAP7_75t_L g391 ( 
.A1(n_389),
.A2(n_382),
.B(n_383),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_391),
.Y(n_393)
);

AOI321xp33_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_390),
.A3(n_392),
.B1(n_12),
.B2(n_13),
.C(n_9),
.Y(n_394)
);

AO221x1_ASAP7_75t_L g395 ( 
.A1(n_394),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_353),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_395),
.A2(n_11),
.B(n_12),
.Y(n_396)
);


endmodule