module fake_jpeg_1606_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_52),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_60),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_59),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_44),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_43),
.B1(n_46),
.B2(n_45),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_42),
.B1(n_1),
.B2(n_2),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_49),
.B(n_39),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_49),
.B(n_43),
.C(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_39),
.B1(n_50),
.B2(n_47),
.Y(n_68)
);

AOI22x1_ASAP7_75t_L g75 ( 
.A1(n_68),
.A2(n_41),
.B1(n_42),
.B2(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_70),
.B(n_38),
.Y(n_74)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_72),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_4),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_71),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_83),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_82),
.B(n_84),
.Y(n_85)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_67),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_5),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_75),
.B(n_5),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_69),
.C(n_61),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_61),
.C(n_20),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_108),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_104),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_18),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_111),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_107),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_23),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_6),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_110),
.B(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_7),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_91),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_27),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_92),
.C(n_25),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_119),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_24),
.C(n_35),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_115),
.Y(n_125)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_36),
.B1(n_16),
.B2(n_30),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_100),
.B1(n_13),
.B2(n_14),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_123),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_135),
.A2(n_138),
.B1(n_116),
.B2(n_122),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_121),
.C(n_132),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_120),
.B1(n_116),
.B2(n_124),
.Y(n_138)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_136),
.B(n_133),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_34),
.Y(n_146)
);


endmodule