module fake_jpeg_14424_n_54 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_54);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_17;
wire n_25;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_6),
.B(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_2),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_28),
.B1(n_23),
.B2(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_27),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_36),
.Y(n_40)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_44),
.C(n_41),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_37),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_47),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_17),
.B(n_42),
.Y(n_47)
);

OAI21xp33_ASAP7_75t_L g48 ( 
.A1(n_47),
.A2(n_21),
.B(n_28),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_29),
.B(n_25),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_20),
.B2(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_53),
.B(n_29),
.Y(n_54)
);


endmodule