module fake_jpeg_17532_n_209 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_46),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_17),
.B1(n_14),
.B2(n_21),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_42),
.B1(n_17),
.B2(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_25),
.A2(n_14),
.B1(n_17),
.B2(n_13),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_45),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_27),
.A2(n_20),
.B(n_23),
.C(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_56),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_17),
.B1(n_28),
.B2(n_32),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_36),
.A2(n_33),
.B1(n_31),
.B2(n_18),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_50),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_47),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_78),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_34),
.B(n_24),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_72),
.B(n_73),
.C(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_34),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_84),
.B(n_92),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_54),
.B1(n_51),
.B2(n_41),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_87),
.B1(n_95),
.B2(n_76),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_62),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_0),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_41),
.B1(n_49),
.B2(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_86),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_22),
.C(n_15),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_61),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_22),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_41),
.B1(n_59),
.B2(n_33),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_103),
.B1(n_67),
.B2(n_75),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_77),
.B(n_64),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_102),
.A2(n_111),
.B(n_91),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_63),
.B1(n_78),
.B2(n_67),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_80),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_85),
.B(n_22),
.C(n_15),
.D(n_71),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_68),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_109),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_85),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_69),
.B(n_67),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_97),
.B(n_15),
.Y(n_138)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_84),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_62),
.B1(n_24),
.B2(n_15),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_81),
.C(n_87),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_98),
.C(n_111),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_118),
.A2(n_126),
.B1(n_101),
.B2(n_106),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_12),
.C(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_121),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_33),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_31),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_98),
.B(n_105),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_131),
.B1(n_6),
.B2(n_10),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_133),
.C(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_96),
.C(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_135),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_104),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_122),
.B1(n_112),
.B2(n_116),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_138),
.A2(n_126),
.B1(n_18),
.B2(n_31),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_9),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_7),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_114),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_148),
.C(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_113),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_112),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_153),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_155),
.A2(n_139),
.B(n_136),
.C(n_145),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_149),
.B1(n_153),
.B2(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_150),
.B1(n_138),
.B2(n_154),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_140),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_143),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_6),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_129),
.C(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_167),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_136),
.C(n_138),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_158),
.B1(n_7),
.B2(n_10),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_168),
.B1(n_167),
.B2(n_166),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_164),
.B1(n_10),
.B2(n_11),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_177),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_3),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_5),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_39),
.C(n_4),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_169),
.B(n_5),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_164),
.B(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_184),
.Y(n_195)
);

AOI21x1_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_4),
.B(n_12),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_186),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_11),
.B(n_12),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_172),
.C(n_176),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_184),
.C(n_39),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_176),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_175),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_199),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_40),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_3),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_3),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_200),
.A2(n_196),
.B(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.C(n_201),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

AOI321xp33_ASAP7_75t_L g206 ( 
.A1(n_204),
.A2(n_198),
.A3(n_40),
.B1(n_2),
.B2(n_1),
.C(n_0),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_39),
.B(n_1),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_0),
.B1(n_2),
.B2(n_191),
.Y(n_209)
);


endmodule