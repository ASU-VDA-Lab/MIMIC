module real_aes_8642_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_729;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g116 ( .A(n_0), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_1), .A2(n_153), .B(n_158), .C(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_2), .A2(n_148), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g464 ( .A(n_3), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_4), .B(n_172), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_5), .A2(n_16), .B1(n_731), .B2(n_732), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_5), .Y(n_732) );
AOI21xp33_ASAP7_75t_L g481 ( .A1(n_6), .A2(n_148), .B(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_L g153 ( .A(n_7), .B(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_8), .A2(n_726), .B1(n_727), .B2(n_728), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_8), .Y(n_726) );
INVx1_ASAP7_75t_L g182 ( .A(n_9), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_10), .B(n_44), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_11), .A2(n_260), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_12), .B(n_163), .Y(n_199) );
INVx1_ASAP7_75t_L g486 ( .A(n_13), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_14), .B(n_162), .Y(n_534) );
INVx1_ASAP7_75t_L g146 ( .A(n_15), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_16), .Y(n_731) );
INVx1_ASAP7_75t_L g546 ( .A(n_17), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_18), .A2(n_183), .B(n_208), .C(n_210), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_19), .B(n_172), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_20), .B(n_475), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_21), .B(n_148), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_22), .B(n_268), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_23), .A2(n_162), .B(n_164), .C(n_168), .Y(n_161) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_24), .A2(n_48), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_24), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_24), .B(n_172), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_25), .B(n_163), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_26), .A2(n_166), .B(n_210), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_27), .B(n_163), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_28), .Y(n_228) );
INVx1_ASAP7_75t_L g242 ( .A(n_29), .Y(n_242) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_30), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_31), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_32), .B(n_163), .Y(n_465) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_33), .A2(n_449), .B1(n_724), .B2(n_725), .C1(n_734), .C2(n_735), .Y(n_448) );
INVx1_ASAP7_75t_L g265 ( .A(n_34), .Y(n_265) );
INVx1_ASAP7_75t_L g499 ( .A(n_35), .Y(n_499) );
INVx2_ASAP7_75t_L g151 ( .A(n_36), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_37), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_38), .A2(n_162), .B(n_221), .C(n_223), .Y(n_220) );
INVxp67_ASAP7_75t_L g266 ( .A(n_39), .Y(n_266) );
CKINVDCx14_ASAP7_75t_R g219 ( .A(n_40), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_41), .A2(n_158), .B(n_241), .C(n_247), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_42), .A2(n_153), .B(n_158), .C(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_43), .A2(n_93), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_43), .Y(n_132) );
INVx1_ASAP7_75t_L g498 ( .A(n_45), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_46), .A2(n_180), .B(n_181), .C(n_184), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_47), .B(n_163), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_48), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_49), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g262 ( .A(n_50), .Y(n_262) );
INVx1_ASAP7_75t_L g156 ( .A(n_51), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_52), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_53), .B(n_148), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_54), .A2(n_158), .B1(n_168), .B2(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_55), .B(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_56), .Y(n_518) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_57), .Y(n_461) );
CKINVDCx14_ASAP7_75t_R g178 ( .A(n_58), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_59), .A2(n_180), .B(n_223), .C(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_60), .Y(n_527) );
INVx1_ASAP7_75t_L g483 ( .A(n_61), .Y(n_483) );
INVx1_ASAP7_75t_L g154 ( .A(n_62), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_63), .A2(n_105), .B1(n_118), .B2(n_739), .Y(n_104) );
INVx1_ASAP7_75t_L g145 ( .A(n_64), .Y(n_145) );
INVx1_ASAP7_75t_SL g222 ( .A(n_65), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_66), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_67), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g231 ( .A(n_68), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_SL g474 ( .A1(n_69), .A2(n_223), .B(n_475), .C(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g477 ( .A(n_70), .Y(n_477) );
INVx1_ASAP7_75t_L g111 ( .A(n_71), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_72), .A2(n_148), .B(n_177), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_73), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_74), .A2(n_148), .B(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_75), .Y(n_502) );
INVx1_ASAP7_75t_L g521 ( .A(n_76), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_77), .A2(n_260), .B(n_261), .Y(n_259) );
INVx1_ASAP7_75t_L g206 ( .A(n_78), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_79), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_80), .A2(n_153), .B(n_158), .C(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_81), .A2(n_148), .B(n_155), .Y(n_147) );
INVx1_ASAP7_75t_L g209 ( .A(n_82), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_83), .B(n_243), .Y(n_515) );
INVx2_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
INVx1_ASAP7_75t_L g196 ( .A(n_85), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_86), .B(n_475), .Y(n_516) );
A2O1A1Ixp33_ASAP7_75t_L g462 ( .A1(n_87), .A2(n_153), .B(n_158), .C(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g113 ( .A(n_88), .B(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g451 ( .A(n_88), .Y(n_451) );
OR2x2_ASAP7_75t_L g723 ( .A(n_88), .B(n_115), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_89), .A2(n_158), .B(n_230), .C(n_233), .Y(n_229) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_90), .A2(n_729), .B1(n_730), .B2(n_733), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_90), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_91), .B(n_175), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_92), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_93), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_94), .A2(n_153), .B(n_158), .C(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_95), .Y(n_538) );
INVx1_ASAP7_75t_L g473 ( .A(n_96), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_97), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_98), .B(n_243), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_99), .B(n_141), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_100), .B(n_141), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g165 ( .A(n_102), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_103), .A2(n_148), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx6p67_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g740 ( .A(n_108), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_113), .Y(n_444) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_114), .B(n_451), .Y(n_737) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OR2x2_ASAP7_75t_L g450 ( .A(n_115), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
AO21x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_447), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_SL g738 ( .A(n_121), .Y(n_738) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_443), .B(n_445), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_129), .B1(n_441), .B2(n_442), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_126), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_129), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_133), .B1(n_439), .B2(n_440), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_130), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_133), .A2(n_450), .B1(n_452), .B2(n_721), .Y(n_449) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g440 ( .A(n_134), .Y(n_440) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_365), .Y(n_134) );
NOR4xp25_ASAP7_75t_L g135 ( .A(n_136), .B(n_307), .C(n_337), .D(n_347), .Y(n_135) );
OAI211xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_212), .B(n_270), .C(n_297), .Y(n_136) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_137), .A2(n_312), .B1(n_393), .B2(n_394), .C1(n_395), .C2(n_396), .Y(n_392) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_187), .Y(n_137) );
AOI33xp33_ASAP7_75t_L g318 ( .A1(n_138), .A2(n_305), .A3(n_306), .B1(n_319), .B2(n_324), .B3(n_326), .Y(n_318) );
OAI211xp5_ASAP7_75t_SL g375 ( .A1(n_138), .A2(n_376), .B(n_378), .C(n_380), .Y(n_375) );
OR2x2_ASAP7_75t_L g391 ( .A(n_138), .B(n_377), .Y(n_391) );
INVx1_ASAP7_75t_L g424 ( .A(n_138), .Y(n_424) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_174), .Y(n_138) );
INVx2_ASAP7_75t_L g301 ( .A(n_139), .Y(n_301) );
AND2x2_ASAP7_75t_L g317 ( .A(n_139), .B(n_203), .Y(n_317) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_139), .Y(n_352) );
AND2x2_ASAP7_75t_L g381 ( .A(n_139), .B(n_174), .Y(n_381) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_147), .B(n_171), .Y(n_139) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_140), .A2(n_204), .B(n_211), .Y(n_203) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_140), .A2(n_217), .B(n_225), .Y(n_216) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_141), .A2(n_471), .B(n_478), .Y(n_470) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g258 ( .A(n_142), .Y(n_258) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x2_ASAP7_75t_SL g175 ( .A(n_143), .B(n_144), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx2_ASAP7_75t_L g260 ( .A(n_148), .Y(n_260) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_149), .B(n_153), .Y(n_193) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g246 ( .A(n_150), .Y(n_246) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
INVx1_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
INVx1_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_152), .Y(n_163) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_152), .Y(n_167) );
INVx3_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
INVx1_ASAP7_75t_L g475 ( .A(n_152), .Y(n_475) );
INVx4_ASAP7_75t_SL g170 ( .A(n_153), .Y(n_170) );
BUFx3_ASAP7_75t_L g247 ( .A(n_153), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_SL g155 ( .A1(n_156), .A2(n_157), .B(n_161), .C(n_170), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g177 ( .A1(n_157), .A2(n_170), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g205 ( .A1(n_157), .A2(n_170), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_157), .A2(n_170), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_SL g261 ( .A1(n_157), .A2(n_170), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_157), .A2(n_170), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_157), .A2(n_170), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_157), .A2(n_170), .B(n_543), .C(n_544), .Y(n_542) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
BUFx3_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_159), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_162), .B(n_222), .Y(n_221) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g180 ( .A(n_163), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_166), .B(n_209), .Y(n_208) );
OAI22xp33_ASAP7_75t_L g264 ( .A1(n_166), .A2(n_243), .B1(n_265), .B2(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_166), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g198 ( .A(n_167), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_167), .A2(n_198), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g466 ( .A(n_168), .Y(n_466) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g233 ( .A(n_170), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_170), .A2(n_193), .B1(n_496), .B2(n_500), .Y(n_495) );
OA21x2_ASAP7_75t_L g480 ( .A1(n_172), .A2(n_481), .B(n_487), .Y(n_480) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_173), .B(n_202), .Y(n_201) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_173), .A2(n_227), .B(n_234), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_173), .B(n_249), .Y(n_248) );
NOR2xp33_ASAP7_75t_SL g517 ( .A(n_173), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g281 ( .A(n_174), .Y(n_281) );
BUFx3_ASAP7_75t_L g289 ( .A(n_174), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_174), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g300 ( .A(n_174), .B(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_174), .B(n_188), .Y(n_329) );
AND2x2_ASAP7_75t_L g398 ( .A(n_174), .B(n_332), .Y(n_398) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_186), .Y(n_174) );
INVx1_ASAP7_75t_L g190 ( .A(n_175), .Y(n_190) );
INVx2_ASAP7_75t_L g236 ( .A(n_175), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_175), .A2(n_193), .B(n_239), .C(n_240), .Y(n_238) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_175), .A2(n_541), .B(n_547), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
INVx5_ASAP7_75t_L g243 ( .A(n_183), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_183), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_183), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g200 ( .A(n_184), .Y(n_200) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g210 ( .A(n_185), .Y(n_210) );
INVx2_ASAP7_75t_SL g292 ( .A(n_187), .Y(n_292) );
OR2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_203), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_188), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g334 ( .A(n_188), .Y(n_334) );
AND2x2_ASAP7_75t_L g345 ( .A(n_188), .B(n_301), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_188), .B(n_330), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_188), .B(n_332), .Y(n_377) );
AND2x2_ASAP7_75t_L g436 ( .A(n_188), .B(n_381), .Y(n_436) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g306 ( .A(n_189), .B(n_203), .Y(n_306) );
AND2x2_ASAP7_75t_L g316 ( .A(n_189), .B(n_317), .Y(n_316) );
BUFx3_ASAP7_75t_L g338 ( .A(n_189), .Y(n_338) );
AND3x2_ASAP7_75t_L g397 ( .A(n_189), .B(n_398), .C(n_399), .Y(n_397) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_201), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_190), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_190), .B(n_527), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_190), .B(n_538), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_194), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_193), .A2(n_228), .B(n_229), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_193), .A2(n_461), .B(n_462), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_193), .A2(n_521), .B(n_522), .Y(n_520) );
O2A1O1Ixp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .C(n_200), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_197), .A2(n_200), .B(n_231), .C(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_200), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_200), .A2(n_524), .B(n_525), .Y(n_523) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
INVx1_ASAP7_75t_SL g332 ( .A(n_203), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g344 ( .A(n_203), .B(n_281), .C(n_345), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_250), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_213), .A2(n_316), .B(n_368), .C(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_215), .B(n_237), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_215), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g384 ( .A(n_215), .Y(n_384) );
AND2x2_ASAP7_75t_L g405 ( .A(n_215), .B(n_252), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_215), .B(n_314), .Y(n_433) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
AND2x2_ASAP7_75t_L g278 ( .A(n_216), .B(n_269), .Y(n_278) );
INVx2_ASAP7_75t_L g285 ( .A(n_216), .Y(n_285) );
AND2x2_ASAP7_75t_L g305 ( .A(n_216), .B(n_252), .Y(n_305) );
AND2x2_ASAP7_75t_L g355 ( .A(n_216), .B(n_237), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_216), .Y(n_359) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_224), .Y(n_535) );
INVx2_ASAP7_75t_SL g269 ( .A(n_226), .Y(n_269) );
BUFx2_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
AND2x2_ASAP7_75t_L g422 ( .A(n_226), .B(n_237), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
INVx1_ASAP7_75t_L g268 ( .A(n_236), .Y(n_268) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_236), .A2(n_530), .B(n_537), .Y(n_529) );
INVx3_ASAP7_75t_SL g252 ( .A(n_237), .Y(n_252) );
AND2x2_ASAP7_75t_L g277 ( .A(n_237), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g284 ( .A(n_237), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g314 ( .A(n_237), .B(n_274), .Y(n_314) );
OR2x2_ASAP7_75t_L g323 ( .A(n_237), .B(n_269), .Y(n_323) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_237), .Y(n_341) );
AND2x2_ASAP7_75t_L g346 ( .A(n_237), .B(n_299), .Y(n_346) );
AND2x2_ASAP7_75t_L g374 ( .A(n_237), .B(n_254), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_237), .B(n_410), .Y(n_409) );
OR2x2_ASAP7_75t_L g412 ( .A(n_237), .B(n_253), .Y(n_412) );
OR2x6_ASAP7_75t_L g237 ( .A(n_238), .B(n_248), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_244), .C(n_245), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_243), .A2(n_464), .B(n_465), .C(n_466), .Y(n_463) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_246), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
AND2x2_ASAP7_75t_L g336 ( .A(n_252), .B(n_285), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_252), .B(n_278), .Y(n_364) );
AND2x2_ASAP7_75t_L g382 ( .A(n_252), .B(n_299), .Y(n_382) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_269), .Y(n_253) );
AND2x2_ASAP7_75t_L g283 ( .A(n_254), .B(n_269), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_254), .B(n_312), .Y(n_311) );
BUFx3_ASAP7_75t_L g321 ( .A(n_254), .Y(n_321) );
OR2x2_ASAP7_75t_L g369 ( .A(n_254), .B(n_289), .Y(n_369) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_259), .B(n_267), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AO21x2_ASAP7_75t_L g274 ( .A1(n_256), .A2(n_275), .B(n_276), .Y(n_274) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_256), .A2(n_520), .B(n_526), .Y(n_519) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AOI21xp5_ASAP7_75t_SL g511 ( .A1(n_257), .A2(n_512), .B(n_513), .Y(n_511) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AO21x2_ASAP7_75t_L g459 ( .A1(n_258), .A2(n_460), .B(n_467), .Y(n_459) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_258), .A2(n_495), .B(n_501), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_258), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g275 ( .A(n_259), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_267), .Y(n_276) );
AND2x2_ASAP7_75t_L g304 ( .A(n_269), .B(n_274), .Y(n_304) );
INVx1_ASAP7_75t_L g312 ( .A(n_269), .Y(n_312) );
AND2x2_ASAP7_75t_L g407 ( .A(n_269), .B(n_285), .Y(n_407) );
AOI222xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_279), .B1(n_282), .B2(n_286), .C1(n_290), .C2(n_293), .Y(n_270) );
INVx1_ASAP7_75t_L g402 ( .A(n_271), .Y(n_402) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_277), .Y(n_271) );
AND2x2_ASAP7_75t_L g298 ( .A(n_272), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g309 ( .A(n_272), .B(n_278), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_272), .B(n_300), .Y(n_325) );
OAI222xp33_ASAP7_75t_L g347 ( .A1(n_272), .A2(n_348), .B1(n_353), .B2(n_354), .C1(n_362), .C2(n_364), .Y(n_347) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g335 ( .A(n_274), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_274), .B(n_355), .Y(n_395) );
AND2x2_ASAP7_75t_L g406 ( .A(n_274), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g414 ( .A(n_277), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_279), .B(n_330), .Y(n_393) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_281), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g351 ( .A(n_281), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx3_ASAP7_75t_L g296 ( .A(n_284), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g386 ( .A1(n_284), .A2(n_387), .B(n_390), .C(n_392), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_284), .B(n_321), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_284), .B(n_304), .Y(n_426) );
AND2x2_ASAP7_75t_L g299 ( .A(n_285), .B(n_295), .Y(n_299) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g326 ( .A(n_288), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_289), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g378 ( .A(n_289), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g417 ( .A(n_289), .B(n_317), .Y(n_417) );
INVx1_ASAP7_75t_L g429 ( .A(n_289), .Y(n_429) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_292), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx1_ASAP7_75t_L g410 ( .A(n_295), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_300), .B(n_302), .C(n_306), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_298), .A2(n_328), .B1(n_343), .B2(n_346), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_299), .B(n_313), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_299), .B(n_321), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_300), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g363 ( .A(n_300), .Y(n_363) );
AND2x2_ASAP7_75t_L g370 ( .A(n_300), .B(n_350), .Y(n_370) );
INVx2_ASAP7_75t_L g331 ( .A(n_301), .Y(n_331) );
INVxp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
NOR4xp25_ASAP7_75t_L g308 ( .A(n_305), .B(n_309), .C(n_310), .D(n_313), .Y(n_308) );
INVx1_ASAP7_75t_SL g379 ( .A(n_306), .Y(n_379) );
AND2x2_ASAP7_75t_L g423 ( .A(n_306), .B(n_424), .Y(n_423) );
OAI211xp5_ASAP7_75t_SL g307 ( .A1(n_308), .A2(n_315), .B(n_318), .C(n_327), .Y(n_307) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_314), .B(n_384), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_316), .A2(n_435), .B1(n_436), .B2(n_437), .Y(n_434) );
INVx1_ASAP7_75t_SL g389 ( .A(n_317), .Y(n_389) );
AND2x2_ASAP7_75t_L g428 ( .A(n_317), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_321), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_325), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_326), .B(n_351), .Y(n_411) );
OAI21xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_333), .B(n_335), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g403 ( .A(n_330), .Y(n_403) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx2_ASAP7_75t_L g431 ( .A(n_331), .Y(n_431) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_332), .Y(n_358) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_339), .B(n_342), .Y(n_337) );
CKINVDCx16_ASAP7_75t_R g350 ( .A(n_338), .Y(n_350) );
OR2x2_ASAP7_75t_L g388 ( .A(n_338), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI21xp33_ASAP7_75t_SL g383 ( .A1(n_341), .A2(n_384), .B(n_385), .Y(n_383) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_345), .A2(n_372), .B1(n_375), .B2(n_382), .C(n_383), .Y(n_371) );
INVx1_ASAP7_75t_SL g415 ( .A(n_346), .Y(n_415) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OR2x2_ASAP7_75t_L g362 ( .A(n_350), .B(n_363), .Y(n_362) );
INVxp67_ASAP7_75t_L g399 ( .A(n_352), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_359), .B2(n_360), .Y(n_354) );
INVx1_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_358), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR4xp25_ASAP7_75t_L g365 ( .A(n_366), .B(n_400), .C(n_413), .D(n_425), .Y(n_365) );
NAND3xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_371), .C(n_386), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_369), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_376), .B(n_381), .Y(n_385) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI221xp5_ASAP7_75t_SL g413 ( .A1(n_388), .A2(n_414), .B1(n_415), .B2(n_416), .C(n_418), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_L g404 ( .A1(n_390), .A2(n_405), .B(n_406), .C(n_408), .Y(n_404) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_391), .A2(n_409), .B1(n_411), .B2(n_412), .Y(n_408) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B(n_403), .C(n_404), .Y(n_400) );
INVx1_ASAP7_75t_L g419 ( .A(n_412), .Y(n_419) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_420), .B(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI221xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_427), .B1(n_430), .B2(n_432), .C(n_434), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_440), .A2(n_450), .B1(n_453), .B2(n_723), .Y(n_734) );
INVx1_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_444), .Y(n_446) );
AOI21xp33_ASAP7_75t_SL g447 ( .A1(n_445), .A2(n_448), .B(n_738), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_637), .Y(n_453) );
NOR5xp2_ASAP7_75t_L g454 ( .A(n_455), .B(n_560), .C(n_592), .D(n_607), .E(n_624), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_488), .B(n_507), .C(n_548), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_469), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_457), .B(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_457), .B(n_612), .Y(n_675) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_458), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_458), .B(n_504), .Y(n_561) );
AND2x2_ASAP7_75t_L g602 ( .A(n_458), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_458), .B(n_571), .Y(n_606) );
OR2x2_ASAP7_75t_L g643 ( .A(n_458), .B(n_494), .Y(n_643) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g493 ( .A(n_459), .B(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g551 ( .A(n_459), .Y(n_551) );
OR2x2_ASAP7_75t_L g714 ( .A(n_459), .B(n_554), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_469), .A2(n_617), .B1(n_618), .B2(n_621), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_469), .B(n_551), .Y(n_700) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_479), .Y(n_469) );
AND2x2_ASAP7_75t_L g506 ( .A(n_470), .B(n_494), .Y(n_506) );
AND2x2_ASAP7_75t_L g553 ( .A(n_470), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g558 ( .A(n_470), .Y(n_558) );
INVx3_ASAP7_75t_L g571 ( .A(n_470), .Y(n_571) );
OR2x2_ASAP7_75t_L g591 ( .A(n_470), .B(n_554), .Y(n_591) );
AND2x2_ASAP7_75t_L g610 ( .A(n_470), .B(n_480), .Y(n_610) );
BUFx2_ASAP7_75t_L g642 ( .A(n_470), .Y(n_642) );
AND2x4_ASAP7_75t_L g557 ( .A(n_479), .B(n_558), .Y(n_557) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g492 ( .A(n_480), .Y(n_492) );
INVx2_ASAP7_75t_L g505 ( .A(n_480), .Y(n_505) );
OR2x2_ASAP7_75t_L g573 ( .A(n_480), .B(n_554), .Y(n_573) );
AND2x2_ASAP7_75t_L g603 ( .A(n_480), .B(n_494), .Y(n_603) );
AND2x2_ASAP7_75t_L g620 ( .A(n_480), .B(n_551), .Y(n_620) );
AND2x2_ASAP7_75t_L g660 ( .A(n_480), .B(n_571), .Y(n_660) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_480), .B(n_506), .Y(n_696) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp33_ASAP7_75t_SL g489 ( .A(n_490), .B(n_503), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_491), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
OAI21xp33_ASAP7_75t_L g634 ( .A1(n_492), .A2(n_506), .B(n_635), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_492), .B(n_494), .Y(n_690) );
AND2x2_ASAP7_75t_L g626 ( .A(n_493), .B(n_627), .Y(n_626) );
INVx3_ASAP7_75t_L g554 ( .A(n_494), .Y(n_554) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_494), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_503), .B(n_551), .Y(n_719) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_504), .A2(n_662), .B1(n_663), .B2(n_668), .Y(n_661) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g552 ( .A(n_505), .B(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g590 ( .A(n_505), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g627 ( .A(n_505), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_506), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g681 ( .A(n_506), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_528), .Y(n_508) );
INVx4_ASAP7_75t_L g567 ( .A(n_509), .Y(n_567) );
AND2x2_ASAP7_75t_L g645 ( .A(n_509), .B(n_612), .Y(n_645) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
INVx3_ASAP7_75t_L g564 ( .A(n_510), .Y(n_564) );
AND2x2_ASAP7_75t_L g578 ( .A(n_510), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
INVx2_ASAP7_75t_L g596 ( .A(n_510), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_510), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g653 ( .A(n_510), .B(n_648), .Y(n_653) );
AND2x2_ASAP7_75t_L g718 ( .A(n_510), .B(n_688), .Y(n_718) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_517), .Y(n_510) );
AND2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_540), .Y(n_559) );
INVx2_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g630 ( .A(n_528), .B(n_578), .Y(n_630) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
INVx2_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
INVx1_ASAP7_75t_L g577 ( .A(n_529), .Y(n_577) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_529), .B(n_579), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_536), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B(n_535), .Y(n_532) );
AND2x2_ASAP7_75t_L g612 ( .A(n_539), .B(n_569), .Y(n_612) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g565 ( .A(n_540), .Y(n_565) );
AND2x2_ASAP7_75t_L g648 ( .A(n_540), .B(n_579), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_555), .B(n_559), .Y(n_548) );
INVx1_ASAP7_75t_SL g593 ( .A(n_549), .Y(n_593) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_550), .B(n_557), .Y(n_650) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g599 ( .A(n_551), .B(n_554), .Y(n_599) );
AND2x2_ASAP7_75t_L g628 ( .A(n_551), .B(n_572), .Y(n_628) );
OR2x2_ASAP7_75t_L g631 ( .A(n_551), .B(n_591), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_552), .A2(n_644), .B1(n_696), .B2(n_697), .C1(n_699), .C2(n_701), .Y(n_695) );
BUFx2_ASAP7_75t_L g609 ( .A(n_554), .Y(n_609) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g598 ( .A(n_557), .B(n_599), .Y(n_598) );
INVx3_ASAP7_75t_SL g615 ( .A(n_557), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_557), .B(n_609), .Y(n_669) );
AND2x2_ASAP7_75t_L g604 ( .A(n_559), .B(n_564), .Y(n_604) );
INVx1_ASAP7_75t_L g623 ( .A(n_559), .Y(n_623) );
OAI221xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_562), .B1(n_566), .B2(n_570), .C(n_574), .Y(n_560) );
OR2x2_ASAP7_75t_L g632 ( .A(n_562), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_587), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_564), .B(n_577), .Y(n_657) );
AND2x2_ASAP7_75t_L g662 ( .A(n_564), .B(n_612), .Y(n_662) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_564), .Y(n_672) );
NAND2x1_ASAP7_75t_SL g683 ( .A(n_564), .B(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g568 ( .A(n_565), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g588 ( .A(n_565), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_565), .B(n_583), .Y(n_614) );
INVx1_ASAP7_75t_L g680 ( .A(n_565), .Y(n_680) );
INVx1_ASAP7_75t_L g655 ( .A(n_566), .Y(n_655) );
OR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx1_ASAP7_75t_L g667 ( .A(n_567), .Y(n_667) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_567), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g684 ( .A(n_568), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_568), .B(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g587 ( .A(n_569), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_569), .B(n_579), .Y(n_600) );
INVx1_ASAP7_75t_L g666 ( .A(n_569), .Y(n_666) );
INVx1_ASAP7_75t_L g687 ( .A(n_570), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_580), .B(n_589), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
AND2x2_ASAP7_75t_L g720 ( .A(n_576), .B(n_653), .Y(n_720) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g688 ( .A(n_577), .B(n_648), .Y(n_688) );
AOI32xp33_ASAP7_75t_L g601 ( .A1(n_578), .A2(n_584), .A3(n_602), .B1(n_604), .B2(n_605), .Y(n_601) );
AOI322xp5_ASAP7_75t_L g703 ( .A1(n_578), .A2(n_610), .A3(n_693), .B1(n_704), .B2(n_705), .C1(n_706), .C2(n_708), .Y(n_703) );
INVx2_ASAP7_75t_L g583 ( .A(n_579), .Y(n_583) );
INVx1_ASAP7_75t_L g693 ( .A(n_579), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_584), .B1(n_585), .B2(n_586), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_581), .B(n_587), .Y(n_636) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_582), .B(n_648), .Y(n_698) );
INVx1_ASAP7_75t_L g585 ( .A(n_583), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_583), .B(n_612), .Y(n_702) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_591), .B(n_686), .Y(n_685) );
OAI221xp5_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B1(n_597), .B2(n_600), .C(n_601), .Y(n_592) );
OR2x2_ASAP7_75t_L g613 ( .A(n_594), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g622 ( .A(n_594), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g647 ( .A(n_595), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g651 ( .A(n_605), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B1(n_613), .B2(n_615), .C(n_616), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_609), .A2(n_640), .B1(n_644), .B2(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_610), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g715 ( .A(n_610), .Y(n_715) );
INVx1_ASAP7_75t_L g709 ( .A(n_612), .Y(n_709) );
INVx1_ASAP7_75t_SL g644 ( .A(n_613), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_615), .B(n_643), .Y(n_705) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_620), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g686 ( .A(n_620), .Y(n_686) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_629), .B1(n_631), .B2(n_632), .C(n_634), .Y(n_624) );
NOR2xp33_ASAP7_75t_SL g625 ( .A(n_626), .B(n_628), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_626), .A2(n_644), .B1(n_690), .B2(n_691), .Y(n_689) );
CKINVDCx14_ASAP7_75t_R g629 ( .A(n_630), .Y(n_629) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_631), .A2(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR3xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_670), .C(n_694), .Y(n_637) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_639), .B(n_646), .C(n_654), .D(n_661), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
INVx1_ASAP7_75t_L g717 ( .A(n_642), .Y(n_717) );
INVx3_ASAP7_75t_SL g711 ( .A(n_643), .Y(n_711) );
OR2x2_ASAP7_75t_L g716 ( .A(n_643), .B(n_717), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_649), .B1(n_651), .B2(n_653), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_648), .B(n_666), .Y(n_707) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI21xp5_ASAP7_75t_SL g654 ( .A1(n_655), .A2(n_656), .B(n_658), .Y(n_654) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OAI211xp5_ASAP7_75t_SL g670 ( .A1(n_671), .A2(n_673), .B(n_676), .C(n_689), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g704 ( .A(n_675), .Y(n_704) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_681), .B1(n_682), .B2(n_685), .C1(n_687), .C2(n_688), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND4xp25_ASAP7_75t_SL g713 ( .A(n_686), .B(n_714), .C(n_715), .D(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND3xp33_ASAP7_75t_SL g694 ( .A(n_695), .B(n_703), .C(n_712), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_718), .B1(n_719), .B2(n_720), .Y(n_712) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
endmodule