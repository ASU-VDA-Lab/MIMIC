module fake_ariane_684_n_2065 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2065);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2065;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_2),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_47),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_26),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_11),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_77),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_149),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_79),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_34),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_32),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_95),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_48),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_170),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_85),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_40),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_56),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_70),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_30),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_120),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_169),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_62),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_33),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_64),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_174),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_152),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_160),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_132),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_175),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_72),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_189),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_113),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_57),
.Y(n_253)
);

BUFx8_ASAP7_75t_SL g254 ( 
.A(n_75),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_96),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_204),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_61),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_62),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_39),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_25),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_164),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_124),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_200),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_73),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_180),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_145),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_119),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_5),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_54),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_22),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_8),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_206),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_32),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_33),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_157),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_188),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_134),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_22),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_93),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_76),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_203),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_137),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_123),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_10),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_142),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_53),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_148),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_19),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_99),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_19),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_54),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_118),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_125),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_41),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_135),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_36),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_64),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_37),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_37),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_130),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_82),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_186),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_71),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_179),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_143),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_154),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_112),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_117),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_2),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_35),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_94),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_7),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_48),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_177),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_197),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_91),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_144),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_136),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_16),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_183),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_50),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_156),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_153),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_201),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_17),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_58),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_176),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_52),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_42),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_81),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_52),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_47),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_0),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_98),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_114),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_88),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_104),
.Y(n_342)
);

BUFx5_ASAP7_75t_L g343 ( 
.A(n_53),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_60),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_162),
.Y(n_345)
);

INVxp33_ASAP7_75t_R g346 ( 
.A(n_35),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_51),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_18),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_109),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_17),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_74),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_129),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_155),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_51),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_58),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_50),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_102),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_45),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_108),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_205),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_168),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_69),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_111),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_89),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_128),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_115),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_107),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_181),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_6),
.Y(n_369)
);

BUFx8_ASAP7_75t_SL g370 ( 
.A(n_198),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_1),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_23),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_56),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_147),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_34),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_139),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_110),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_46),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_61),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_103),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_161),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_138),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_28),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_43),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_18),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_39),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_41),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_24),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_171),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_44),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_67),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_4),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_184),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_1),
.Y(n_394)
);

BUFx10_ASAP7_75t_L g395 ( 
.A(n_28),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_24),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_126),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_173),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_6),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_13),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_29),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_191),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_26),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_131),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_46),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_87),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_92),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_16),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_106),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_57),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_42),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_116),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_15),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_68),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_254),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_343),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_343),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_375),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_343),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_343),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_233),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_343),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_370),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_252),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_302),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_249),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_229),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_229),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_229),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_349),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_229),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_229),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_210),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_376),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_258),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_378),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_247),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_379),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_260),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_261),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_210),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_271),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_375),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_371),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_211),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_211),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_272),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_223),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_213),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_223),
.Y(n_459)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_379),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_303),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_214),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_215),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_399),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_217),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_303),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_314),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_314),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_275),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_276),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_318),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_222),
.Y(n_473)
);

CKINVDCx14_ASAP7_75t_R g474 ( 
.A(n_269),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_318),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_214),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_324),
.Y(n_477)
);

INVxp67_ASAP7_75t_SL g478 ( 
.A(n_324),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_279),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_358),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_395),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_293),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_225),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_395),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_383),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_383),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_264),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_264),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_269),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_216),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_308),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_216),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_295),
.Y(n_494)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_237),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_269),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_308),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_310),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_310),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_299),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_225),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_380),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_321),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_321),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_363),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_395),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_245),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_241),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_363),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_245),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_301),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_304),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_315),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_402),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_317),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_406),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_406),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_242),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_262),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_380),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_330),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_418),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_418),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_478),
.B(n_234),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_452),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_419),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_465),
.A2(n_435),
.B1(n_439),
.B2(n_427),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_422),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_340),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_422),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_425),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_425),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_430),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_430),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_467),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_462),
.B(n_351),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_474),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_432),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_417),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_432),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_473),
.B(n_421),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_433),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_433),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_434),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_434),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_436),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_436),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_441),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_441),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_431),
.B(n_451),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_442),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_462),
.B(n_249),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_443),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_443),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_447),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_447),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_453),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_453),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_420),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_488),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_476),
.B(n_332),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_488),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_489),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_440),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_489),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_492),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_492),
.A2(n_332),
.B(n_219),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_497),
.Y(n_580)
);

INVxp33_ASAP7_75t_SL g581 ( 
.A(n_426),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_467),
.B(n_380),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_431),
.B(n_476),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_497),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_498),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_498),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_446),
.B(n_332),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_491),
.B(n_218),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_491),
.B(n_221),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_416),
.A2(n_253),
.B1(n_356),
.B2(n_348),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_503),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_448),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_504),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_504),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_493),
.B(n_262),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_505),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_514),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_514),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_515),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_493),
.B(n_243),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_520),
.B(n_259),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_424),
.Y(n_608)
);

AND2x4_ASAP7_75t_L g609 ( 
.A(n_520),
.B(n_273),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g610 ( 
.A(n_583),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_576),
.B(n_444),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_550),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_534),
.A2(n_438),
.B1(n_484),
.B2(n_449),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_548),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

AOI21x1_ASAP7_75t_L g616 ( 
.A1(n_533),
.A2(n_517),
.B(n_515),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_544),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_544),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_582),
.B(n_463),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_526),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_575),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_526),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_431),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_526),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_L g625 ( 
.A(n_525),
.B(n_389),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_576),
.B(n_450),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_550),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_L g628 ( 
.A(n_525),
.B(n_389),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_561),
.A2(n_333),
.B1(n_348),
.B2(n_253),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_526),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_523),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_550),
.B(n_482),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_525),
.B(n_389),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_582),
.B(n_495),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_523),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_588),
.B(n_470),
.C(n_456),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_523),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_571),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_527),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_582),
.B(n_508),
.Y(n_640)
);

BUFx10_ASAP7_75t_L g641 ( 
.A(n_595),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_527),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_576),
.B(n_471),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_525),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_561),
.B(n_479),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_530),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_588),
.A2(n_494),
.B1(n_500),
.B2(n_483),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_576),
.B(n_511),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_530),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_525),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_530),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_538),
.B(n_431),
.Y(n_653)
);

INVxp33_ASAP7_75t_L g654 ( 
.A(n_571),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_548),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_525),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_576),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_531),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_540),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_595),
.B(n_512),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_531),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_525),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_536),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_531),
.Y(n_664)
);

INVx5_ASAP7_75t_L g665 ( 
.A(n_536),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_534),
.B(n_445),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_535),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_534),
.B(n_513),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_546),
.B(n_516),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_528),
.B(n_522),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_546),
.B(n_460),
.Y(n_671)
);

NOR3xp33_ASAP7_75t_L g672 ( 
.A(n_593),
.B(n_362),
.C(n_356),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_575),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_535),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_535),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_540),
.B(n_518),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_549),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_536),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_549),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_552),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_552),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_529),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_564),
.A2(n_501),
.B1(n_510),
.B2(n_507),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_554),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_553),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_541),
.B(n_464),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_541),
.B(n_485),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_524),
.B(n_506),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_553),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_542),
.B(n_519),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_529),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_554),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_542),
.B(n_353),
.Y(n_694)
);

BUFx2_ASAP7_75t_L g695 ( 
.A(n_524),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_524),
.B(n_564),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_578),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_606),
.B(n_607),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_543),
.B(n_353),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_543),
.B(n_466),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_536),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_578),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_580),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_564),
.B(n_212),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_564),
.B(n_212),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_536),
.B(n_389),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_564),
.B(n_220),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_545),
.B(n_490),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_558),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_536),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_581),
.B(n_220),
.Y(n_712)
);

AO21x2_ASAP7_75t_L g713 ( 
.A1(n_579),
.A2(n_230),
.B(n_227),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_558),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_554),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_599),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_606),
.B(n_467),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_556),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_581),
.B(n_226),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_608),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

CKINVDCx6p67_ASAP7_75t_R g722 ( 
.A(n_608),
.Y(n_722)
);

AND3x4_ASAP7_75t_L g723 ( 
.A(n_606),
.B(n_346),
.C(n_413),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_536),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_556),
.Y(n_725)
);

BUFx10_ASAP7_75t_L g726 ( 
.A(n_573),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_560),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_556),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_562),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_545),
.B(n_226),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_606),
.B(n_454),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_556),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_606),
.B(n_228),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_607),
.B(n_454),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_537),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_562),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_537),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_532),
.Y(n_738)
);

AOI21x1_ASAP7_75t_L g739 ( 
.A1(n_579),
.A2(n_248),
.B(n_232),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_593),
.A2(n_369),
.B1(n_373),
.B2(n_362),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_607),
.B(n_228),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_532),
.A2(n_496),
.B1(n_521),
.B2(n_502),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_580),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_556),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_589),
.B(n_257),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_584),
.Y(n_746)
);

BUFx4f_ASAP7_75t_L g747 ( 
.A(n_572),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_567),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_607),
.B(n_455),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_599),
.B(n_224),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_607),
.B(n_231),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_565),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_565),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_599),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_584),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_567),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_566),
.Y(n_757)
);

AO21x2_ASAP7_75t_L g758 ( 
.A1(n_579),
.A2(n_280),
.B(n_274),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_726),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_651),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_657),
.B(n_369),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_638),
.Y(n_762)
);

OR2x6_ASAP7_75t_L g763 ( 
.A(n_695),
.B(n_609),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_657),
.B(n_609),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_670),
.B(n_283),
.C(n_278),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_610),
.B(n_599),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_648),
.B(n_609),
.Y(n_767)
);

O2A1O1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_617),
.A2(n_596),
.B(n_291),
.C(n_296),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_612),
.B(n_609),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_631),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_615),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_651),
.B(n_537),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_646),
.B(n_596),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_612),
.A2(n_596),
.B1(n_574),
.B2(n_577),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_627),
.B(n_596),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_619),
.A2(n_573),
.B1(n_596),
.B2(n_590),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_615),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_651),
.B(n_537),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_651),
.B(n_537),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_627),
.B(n_573),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_631),
.Y(n_781)
);

AO22x2_ASAP7_75t_L g782 ( 
.A1(n_723),
.A2(n_573),
.B1(n_590),
.B2(n_585),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_634),
.B(n_591),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_662),
.B(n_539),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_659),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_618),
.B(n_591),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_619),
.A2(n_592),
.B1(n_594),
.B2(n_585),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_619),
.A2(n_594),
.B1(n_597),
.B2(n_592),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_614),
.B(n_413),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_634),
.B(n_597),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_659),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_677),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_663),
.A2(n_539),
.B(n_567),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_623),
.B(n_539),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_731),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_686),
.B(n_539),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_636),
.B(n_231),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_687),
.B(n_539),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_640),
.B(n_235),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_598),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_619),
.B(n_745),
.Y(n_801)
);

NOR2xp67_ASAP7_75t_SL g802 ( 
.A(n_626),
.B(n_373),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_639),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_645),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_691),
.B(n_600),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_666),
.B(n_600),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_716),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_726),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_632),
.B(n_601),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_641),
.B(n_235),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_694),
.A2(n_601),
.B1(n_236),
.B2(n_239),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_672),
.A2(n_574),
.B1(n_602),
.B2(n_577),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_632),
.B(n_574),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_701),
.A2(n_326),
.B(n_337),
.C(n_289),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_695),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_645),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_668),
.B(n_539),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_662),
.B(n_539),
.Y(n_818)
);

AND2x2_ASAP7_75t_SL g819 ( 
.A(n_699),
.B(n_281),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_662),
.B(n_572),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_731),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_700),
.B(n_577),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_696),
.B(n_605),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_638),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_SL g825 ( 
.A1(n_692),
.A2(n_385),
.B1(n_391),
.B2(n_390),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_754),
.B(n_602),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_679),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_658),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_709),
.A2(n_313),
.B1(n_412),
.B2(n_409),
.Y(n_829)
);

AND2x6_ASAP7_75t_L g830 ( 
.A(n_699),
.B(n_586),
.Y(n_830)
);

BUFx3_ASAP7_75t_L g831 ( 
.A(n_614),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_692),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_653),
.A2(n_385),
.B1(n_390),
.B2(n_388),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_658),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_717),
.B(n_350),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_730),
.B(n_602),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_716),
.B(n_604),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_621),
.B(n_604),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_680),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_635),
.A2(n_586),
.B(n_568),
.C(n_567),
.Y(n_840)
);

AND2x2_ASAP7_75t_SL g841 ( 
.A(n_717),
.B(n_284),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_662),
.B(n_572),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_680),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_673),
.B(n_604),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_697),
.B(n_605),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_661),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_643),
.B(n_605),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_703),
.B(n_586),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_649),
.B(n_586),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_661),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_664),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_704),
.B(n_572),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_743),
.B(n_746),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_678),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_755),
.B(n_572),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_664),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_681),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_641),
.B(n_236),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_750),
.B(n_572),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_667),
.Y(n_860)
);

NOR2x1p5_ASAP7_75t_L g861 ( 
.A(n_655),
.B(n_384),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_733),
.B(n_572),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_666),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_678),
.B(n_587),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_587),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_734),
.B(n_587),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_641),
.B(n_238),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_741),
.B(n_751),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_726),
.A2(n_352),
.B1(n_239),
.B2(n_412),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_705),
.B(n_587),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_654),
.B(n_413),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_734),
.B(n_587),
.Y(n_872)
);

OAI22xp33_ASAP7_75t_L g873 ( 
.A1(n_740),
.A2(n_386),
.B1(n_411),
.B2(n_410),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_613),
.B(n_387),
.C(n_384),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_678),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_731),
.A2(n_352),
.B1(n_240),
.B2(n_409),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_681),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_L g878 ( 
.A(n_660),
.B(n_355),
.C(n_354),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_616),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_635),
.B(n_587),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_637),
.B(n_587),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_685),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_637),
.B(n_642),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_667),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_674),
.Y(n_885)
);

INVx2_ASAP7_75t_SL g886 ( 
.A(n_682),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_642),
.B(n_603),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_731),
.B(n_372),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_749),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_678),
.B(n_603),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_678),
.B(n_603),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_647),
.B(n_603),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_690),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_702),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_647),
.B(n_603),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_650),
.B(n_603),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_702),
.B(n_238),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_749),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_655),
.B(n_455),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_749),
.B(n_394),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_710),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_652),
.A2(n_569),
.B1(n_566),
.B2(n_551),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_720),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_710),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_652),
.B(n_567),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_714),
.Y(n_906)
);

BUFx6f_ASAP7_75t_SL g907 ( 
.A(n_722),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_706),
.B(n_331),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_611),
.B(n_240),
.Y(n_909)
);

INVxp67_ASAP7_75t_SL g910 ( 
.A(n_702),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_714),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_R g912 ( 
.A(n_720),
.B(n_387),
.Y(n_912)
);

OAI22xp33_ASAP7_75t_L g913 ( 
.A1(n_749),
.A2(n_400),
.B1(n_403),
.B2(n_408),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_683),
.B(n_244),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_712),
.B(n_244),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_688),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_719),
.B(n_246),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_708),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_629),
.B(n_457),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_762),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_819),
.A2(n_723),
.B1(n_738),
.B2(n_675),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_783),
.B(n_674),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_786),
.A2(n_721),
.B(n_729),
.C(n_727),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_792),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_831),
.Y(n_925)
);

AO22x1_ASAP7_75t_L g926 ( 
.A1(n_832),
.A2(n_738),
.B1(n_722),
.B2(n_742),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_786),
.B(n_675),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_790),
.B(n_620),
.Y(n_928)
);

AND2x6_ASAP7_75t_L g929 ( 
.A(n_759),
.B(n_808),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_800),
.B(n_620),
.Y(n_930)
);

OAI21xp33_ASAP7_75t_SL g931 ( 
.A1(n_819),
.A2(n_729),
.B(n_727),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_813),
.B(n_809),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_795),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_762),
.B(n_671),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_801),
.B(n_669),
.Y(n_935)
);

AO21x1_ASAP7_75t_L g936 ( 
.A1(n_794),
.A2(n_676),
.B(n_736),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_815),
.B(n_457),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_907),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_795),
.B(n_736),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_821),
.B(n_889),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_770),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_841),
.B(n_622),
.Y(n_942)
);

AO22x1_ASAP7_75t_L g943 ( 
.A1(n_903),
.A2(n_388),
.B1(n_391),
.B2(n_334),
.Y(n_943)
);

AND2x6_ASAP7_75t_SL g944 ( 
.A(n_763),
.B(n_396),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_841),
.B(n_624),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_899),
.B(n_459),
.Y(n_946)
);

NOR2x2_ASAP7_75t_L g947 ( 
.A(n_763),
.B(n_684),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_916),
.B(n_724),
.Y(n_948)
);

INVxp67_ASAP7_75t_SL g949 ( 
.A(n_898),
.Y(n_949)
);

INVxp67_ASAP7_75t_SL g950 ( 
.A(n_898),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_821),
.B(n_702),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_773),
.A2(n_752),
.B1(n_757),
.B2(n_753),
.Y(n_952)
);

OR2x6_ASAP7_75t_L g953 ( 
.A(n_889),
.B(n_752),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_827),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_886),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_830),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_822),
.B(n_919),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_830),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_824),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_839),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_763),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_912),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_781),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_830),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_766),
.B(n_624),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_843),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_805),
.B(n_630),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_912),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_873),
.A2(n_753),
.B(n_757),
.C(n_756),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_780),
.B(n_823),
.Y(n_970)
);

NAND3xp33_ASAP7_75t_SL g971 ( 
.A(n_789),
.B(n_338),
.C(n_336),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_R g972 ( 
.A(n_907),
.B(n_616),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_830),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_830),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_823),
.B(n_630),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_857),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_759),
.B(n_724),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_782),
.A2(n_569),
.B1(n_570),
.B2(n_551),
.Y(n_978)
);

INVxp67_ASAP7_75t_SL g979 ( 
.A(n_807),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_803),
.Y(n_980)
);

AO22x1_ASAP7_75t_L g981 ( 
.A1(n_765),
.A2(n_863),
.B1(n_900),
.B2(n_888),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_877),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_760),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_888),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_769),
.B(n_684),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_808),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_882),
.B(n_689),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_871),
.B(n_459),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_782),
.A2(n_563),
.B1(n_551),
.B2(n_559),
.Y(n_989)
);

INVx4_ASAP7_75t_L g990 ( 
.A(n_760),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_806),
.Y(n_991)
);

NOR2x1p5_ASAP7_75t_L g992 ( 
.A(n_874),
.B(n_344),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_893),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_901),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_900),
.B(n_693),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_782),
.A2(n_570),
.B1(n_559),
.B2(n_563),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_804),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_760),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_835),
.B(n_698),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_799),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_904),
.B(n_698),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_906),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_911),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_853),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_835),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_868),
.B(n_644),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_760),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_816),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_873),
.A2(n_913),
.B1(n_774),
.B2(n_825),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_868),
.Y(n_1010)
);

O2A1O1Ixp5_ASAP7_75t_L g1011 ( 
.A1(n_897),
.A2(n_747),
.B(n_711),
.C(n_735),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_829),
.B(n_461),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_854),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_838),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_774),
.B(n_715),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_828),
.Y(n_1016)
);

AND3x2_ASAP7_75t_SL g1017 ( 
.A(n_913),
.B(n_563),
.C(n_559),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_854),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_854),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_875),
.B(n_718),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_844),
.Y(n_1021)
);

AND2x2_ASAP7_75t_SL g1022 ( 
.A(n_776),
.B(n_625),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_918),
.B(n_718),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_796),
.B(n_725),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_875),
.B(n_725),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_875),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_845),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_768),
.A2(n_756),
.B(n_748),
.C(n_728),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_875),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_834),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_861),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_866),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_865),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_846),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_872),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_787),
.B(n_728),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_771),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_848),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_788),
.B(n_817),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_777),
.B(n_732),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_SL g1041 ( 
.A1(n_794),
.A2(n_644),
.B(n_711),
.C(n_735),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_775),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_850),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_851),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_826),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_852),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_796),
.B(n_732),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_914),
.A2(n_570),
.B1(n_748),
.B2(n_744),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_798),
.B(n_744),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_856),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_798),
.B(n_644),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_855),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_810),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_785),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_767),
.A2(n_711),
.B1(n_735),
.B2(n_737),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_908),
.A2(n_737),
.B1(n_625),
.B2(n_707),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_860),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_858),
.Y(n_1058)
);

NOR2x2_ASAP7_75t_L g1059 ( 
.A(n_876),
.B(n_347),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_867),
.Y(n_1060)
);

AOI21xp33_ASAP7_75t_L g1061 ( 
.A1(n_908),
.A2(n_737),
.B(n_633),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_791),
.B(n_656),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_884),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_878),
.B(n_461),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_909),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_905),
.Y(n_1066)
);

NOR2x2_ASAP7_75t_L g1067 ( 
.A(n_802),
.B(n_405),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_797),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_885),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_817),
.B(n_656),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_883),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_772),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_811),
.B(n_656),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_836),
.B(n_656),
.Y(n_1074)
);

OAI22xp5_ASAP7_75t_L g1075 ( 
.A1(n_764),
.A2(n_747),
.B1(n_414),
.B2(n_665),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_837),
.A2(n_555),
.B1(n_557),
.B2(n_469),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_836),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_879),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_915),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_879),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_917),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_869),
.B(n_468),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_880),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_881),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_887),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_892),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_L g1087 ( 
.A(n_833),
.B(n_568),
.C(n_298),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_895),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_894),
.B(n_665),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_847),
.B(n_665),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_847),
.B(n_665),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_910),
.B(n_812),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_896),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_849),
.B(n_665),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_772),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_812),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_849),
.B(n_468),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_859),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_820),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_840),
.Y(n_1100)
);

AND2x6_ASAP7_75t_SL g1101 ( 
.A(n_870),
.B(n_469),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_761),
.B(n_747),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_1096),
.A2(n_902),
.B1(n_870),
.B2(n_862),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_931),
.A2(n_862),
.B(n_814),
.C(n_793),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_932),
.B(n_1004),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_956),
.B(n_820),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_973),
.B(n_778),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_927),
.A2(n_779),
.B(n_778),
.Y(n_1108)
);

INVx2_ASAP7_75t_SL g1109 ( 
.A(n_925),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_957),
.B(n_1032),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_973),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_973),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_933),
.B(n_779),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_956),
.B(n_958),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_1009),
.B(n_897),
.C(n_902),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_991),
.B(n_472),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_920),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1035),
.B(n_784),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_973),
.B(n_246),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_952),
.A2(n_818),
.B(n_891),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_958),
.B(n_891),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1024),
.A2(n_818),
.B(n_842),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1047),
.A2(n_890),
.B(n_864),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_920),
.B(n_472),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_933),
.Y(n_1125)
);

O2A1O1Ixp5_ASAP7_75t_L g1126 ( 
.A1(n_936),
.A2(n_890),
.B(n_864),
.C(n_842),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_SL g1127 ( 
.A1(n_923),
.A2(n_381),
.B(n_382),
.C(n_397),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_925),
.B(n_475),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_964),
.B(n_974),
.Y(n_1129)
);

OA22x2_ASAP7_75t_L g1130 ( 
.A1(n_1005),
.A2(n_480),
.B1(n_475),
.B2(n_477),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_964),
.Y(n_1131)
);

INVx5_ASAP7_75t_L g1132 ( 
.A(n_939),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_998),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_935),
.A2(n_628),
.B(n_707),
.C(n_633),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_984),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_938),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_924),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_974),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_1010),
.B(n_286),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_998),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1096),
.B(n_568),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1009),
.A2(n_568),
.B1(n_739),
.B2(n_327),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_941),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_935),
.B(n_250),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_998),
.Y(n_1145)
);

AO32x1_ASAP7_75t_L g1146 ( 
.A1(n_1099),
.A2(n_557),
.A3(n_555),
.B1(n_480),
.B2(n_481),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_963),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_923),
.A2(n_628),
.B(n_713),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_963),
.Y(n_1149)
);

AO31x2_ASAP7_75t_L g1150 ( 
.A1(n_1098),
.A2(n_557),
.A3(n_555),
.B(n_486),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_940),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_984),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_959),
.B(n_288),
.Y(n_1153)
);

NAND3xp33_ASAP7_75t_L g1154 ( 
.A(n_1006),
.B(n_568),
.C(n_547),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1049),
.A2(n_758),
.B(n_713),
.Y(n_1155)
);

AND2x6_ASAP7_75t_L g1156 ( 
.A(n_1092),
.B(n_294),
.Y(n_1156)
);

AO21x2_ASAP7_75t_L g1157 ( 
.A1(n_1041),
.A2(n_758),
.B(n_713),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_981),
.B(n_250),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_L g1159 ( 
.A(n_971),
.B(n_486),
.C(n_477),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_968),
.B(n_251),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_1077),
.B(n_251),
.Y(n_1161)
);

BUFx4f_ASAP7_75t_SL g1162 ( 
.A(n_962),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1039),
.A2(n_758),
.B(n_481),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1018),
.B(n_555),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_955),
.B(n_312),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_955),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_998),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_940),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_980),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_961),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1000),
.B(n_312),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_939),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_954),
.A2(n_361),
.B1(n_300),
.B2(n_341),
.Y(n_1173)
);

BUFx12f_ASAP7_75t_L g1174 ( 
.A(n_944),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_934),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_921),
.B(n_946),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_947),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_L g1178 ( 
.A1(n_1006),
.A2(n_313),
.B(n_357),
.Y(n_1178)
);

OAI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_357),
.B1(n_366),
.B2(n_359),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1014),
.B(n_547),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1021),
.B(n_547),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_948),
.A2(n_359),
.B1(n_360),
.B2(n_364),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_949),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_948),
.B(n_360),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_997),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1071),
.B(n_365),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1071),
.B(n_365),
.Y(n_1187)
);

INVxp67_ASAP7_75t_L g1188 ( 
.A(n_937),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1018),
.Y(n_1189)
);

INVx2_ASAP7_75t_SL g1190 ( 
.A(n_1031),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_988),
.B(n_487),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_997),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1051),
.A2(n_311),
.B(n_407),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_947),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1027),
.B(n_547),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_939),
.Y(n_1196)
);

OAI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1087),
.A2(n_367),
.B(n_368),
.Y(n_1197)
);

OR2x6_ASAP7_75t_SL g1198 ( 
.A(n_1059),
.B(n_367),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_950),
.B(n_374),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_960),
.Y(n_1200)
);

BUFx2_ASAP7_75t_SL g1201 ( 
.A(n_1018),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1008),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1067),
.B(n_374),
.C(n_377),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1101),
.B(n_255),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_1042),
.A2(n_307),
.B(n_404),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_966),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_970),
.A2(n_306),
.B(n_398),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1008),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1012),
.B(n_547),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1033),
.B(n_256),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1053),
.B(n_263),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1082),
.B(n_0),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1018),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1078),
.A2(n_389),
.B(n_209),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_976),
.A2(n_305),
.B1(n_345),
.B2(n_342),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_995),
.Y(n_1216)
);

NOR3xp33_ASAP7_75t_SL g1217 ( 
.A(n_1067),
.B(n_393),
.C(n_339),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_967),
.A2(n_297),
.B(n_335),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1058),
.B(n_265),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1016),
.Y(n_1220)
);

O2A1O1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_969),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_1221)
);

INVx4_ASAP7_75t_L g1222 ( 
.A(n_953),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1091),
.A2(n_292),
.B(n_329),
.C(n_328),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1019),
.B(n_209),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1064),
.B(n_3),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1016),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1030),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1019),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_995),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1033),
.B(n_266),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_1091),
.A2(n_389),
.B(n_319),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1038),
.B(n_7),
.Y(n_1232)
);

O2A1O1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1028),
.A2(n_8),
.B(n_9),
.C(n_12),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_953),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_982),
.A2(n_287),
.B1(n_323),
.B2(n_322),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_993),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_994),
.A2(n_325),
.B1(n_320),
.B2(n_267),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1080),
.A2(n_319),
.B(n_290),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1030),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_995),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_943),
.B(n_9),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_926),
.B(n_12),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1061),
.A2(n_282),
.B(n_316),
.C(n_309),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1019),
.Y(n_1244)
);

O2A1O1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1028),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_942),
.A2(n_285),
.B(n_277),
.C(n_270),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_945),
.A2(n_268),
.B(n_290),
.C(n_319),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1068),
.B(n_14),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_922),
.B(n_20),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1041),
.A2(n_319),
.B(n_290),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1045),
.B(n_20),
.Y(n_1251)
);

INVx3_ASAP7_75t_SL g1252 ( 
.A(n_1059),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_999),
.B(n_21),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1033),
.B(n_319),
.Y(n_1254)
);

INVx6_ASAP7_75t_L g1255 ( 
.A(n_1128),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1238),
.A2(n_1011),
.B(n_1080),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1137),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1105),
.B(n_1045),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1105),
.A2(n_1094),
.B(n_1090),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1136),
.Y(n_1260)
);

BUFx4f_ASAP7_75t_L g1261 ( 
.A(n_1189),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1104),
.A2(n_1056),
.B(n_1100),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1110),
.B(n_1092),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1139),
.A2(n_953),
.B1(n_1065),
.B2(n_1079),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1148),
.A2(n_965),
.B(n_928),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1188),
.B(n_999),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1250),
.A2(n_1074),
.B(n_975),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1162),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1120),
.A2(n_930),
.B(n_1102),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1214),
.A2(n_1025),
.B(n_1020),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1117),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1148),
.A2(n_1015),
.B(n_1022),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1110),
.B(n_1098),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1250),
.A2(n_1099),
.B(n_951),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1103),
.A2(n_1070),
.B(n_979),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1129),
.B(n_999),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1155),
.A2(n_1052),
.B(n_1046),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_SL g1278 ( 
.A1(n_1223),
.A2(n_1066),
.B(n_1001),
.C(n_987),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1115),
.B(n_1036),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1176),
.B(n_1175),
.Y(n_1280)
);

NAND2x1_ASAP7_75t_L g1281 ( 
.A(n_1111),
.B(n_929),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1189),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1143),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1147),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1231),
.A2(n_1086),
.B(n_1083),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1212),
.B(n_1097),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1200),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1109),
.B(n_1081),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1103),
.A2(n_1002),
.B1(n_1003),
.B2(n_1022),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1122),
.A2(n_1123),
.B(n_1108),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1206),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1236),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1135),
.B(n_1023),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1124),
.B(n_1152),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1156),
.B(n_1036),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1221),
.A2(n_1037),
.B(n_992),
.C(n_1036),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1163),
.A2(n_1088),
.B(n_1093),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1163),
.A2(n_1073),
.B(n_1062),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1241),
.A2(n_978),
.B(n_1017),
.Y(n_1299)
);

AO32x2_ASAP7_75t_L g1300 ( 
.A1(n_1142),
.A2(n_1017),
.A3(n_990),
.B1(n_1075),
.B2(n_978),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1170),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1191),
.B(n_1023),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1149),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1134),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1183),
.B(n_1023),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1157),
.A2(n_1085),
.B(n_1084),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1153),
.B(n_1054),
.Y(n_1307)
);

AO21x2_ASAP7_75t_L g1308 ( 
.A1(n_1157),
.A2(n_1084),
.B(n_985),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1156),
.B(n_1033),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1249),
.A2(n_1070),
.B(n_1007),
.Y(n_1310)
);

A2O1A1Ixp33_ASAP7_75t_L g1311 ( 
.A1(n_1197),
.A2(n_1070),
.B(n_1040),
.C(n_996),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1247),
.A2(n_1044),
.A3(n_1050),
.B(n_1034),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1169),
.Y(n_1313)
);

INVxp67_ASAP7_75t_SL g1314 ( 
.A(n_1216),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1142),
.A2(n_1055),
.B(n_1048),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1249),
.A2(n_1026),
.B(n_1007),
.Y(n_1316)
);

O2A1O1Ixp5_ASAP7_75t_SL g1317 ( 
.A1(n_1254),
.A2(n_1069),
.B(n_986),
.C(n_1013),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1189),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1131),
.B(n_972),
.Y(n_1319)
);

OAI22x1_ASAP7_75t_L g1320 ( 
.A1(n_1252),
.A2(n_1040),
.B1(n_986),
.B2(n_1050),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1232),
.A2(n_1118),
.B(n_1180),
.Y(n_1321)
);

AND4x1_ASAP7_75t_L g1322 ( 
.A(n_1203),
.B(n_989),
.C(n_996),
.D(n_1048),
.Y(n_1322)
);

NOR3xp33_ASAP7_75t_SL g1323 ( 
.A(n_1160),
.B(n_972),
.C(n_23),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1161),
.B(n_989),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1204),
.B(n_1095),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1190),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1213),
.Y(n_1327)
);

AO32x2_ASAP7_75t_L g1328 ( 
.A1(n_1173),
.A2(n_990),
.A3(n_1072),
.B1(n_1095),
.B2(n_1076),
.Y(n_1328)
);

O2A1O1Ixp5_ASAP7_75t_L g1329 ( 
.A1(n_1184),
.A2(n_1144),
.B(n_1119),
.C(n_1210),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1232),
.A2(n_977),
.B(n_1089),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1224),
.A2(n_1141),
.B(n_1107),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1127),
.A2(n_1118),
.B(n_1141),
.Y(n_1332)
);

INVx1_ASAP7_75t_SL g1333 ( 
.A(n_1253),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1185),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1180),
.A2(n_977),
.B(n_1089),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1192),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1156),
.B(n_929),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1178),
.A2(n_1245),
.B(n_1233),
.C(n_1248),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1166),
.B(n_983),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1156),
.B(n_929),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1202),
.Y(n_1341)
);

BUFx8_ASAP7_75t_L g1342 ( 
.A(n_1174),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1128),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1181),
.A2(n_1089),
.B(n_983),
.Y(n_1344)
);

O2A1O1Ixp5_ASAP7_75t_L g1345 ( 
.A1(n_1230),
.A2(n_1043),
.B(n_1034),
.C(n_1057),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1114),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1195),
.A2(n_1243),
.B(n_1251),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1208),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1114),
.A2(n_1029),
.B(n_1095),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1199),
.B(n_929),
.Y(n_1350)
);

AND3x1_ASAP7_75t_L g1351 ( 
.A(n_1217),
.B(n_21),
.C(n_25),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1220),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1226),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1225),
.A2(n_1029),
.B(n_1072),
.C(n_1095),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1234),
.A2(n_1072),
.B(n_1063),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1251),
.A2(n_1072),
.B(n_1063),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1114),
.A2(n_1063),
.B(n_290),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1227),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1239),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1246),
.A2(n_27),
.B(n_29),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1164),
.A2(n_90),
.B(n_199),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1164),
.A2(n_84),
.B(n_192),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1106),
.A2(n_209),
.B(n_83),
.Y(n_1363)
);

O2A1O1Ixp5_ASAP7_75t_L g1364 ( 
.A1(n_1186),
.A2(n_27),
.B(n_30),
.C(n_31),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1111),
.A2(n_97),
.B(n_190),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1207),
.A2(n_31),
.B(n_36),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_L g1367 ( 
.A(n_1182),
.B(n_209),
.C(n_43),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1179),
.A2(n_38),
.B(n_44),
.C(n_49),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1131),
.B(n_38),
.Y(n_1369)
);

OAI22x1_ASAP7_75t_L g1370 ( 
.A1(n_1242),
.A2(n_49),
.B1(n_55),
.B2(n_59),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1112),
.A2(n_121),
.B(n_187),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1106),
.A2(n_209),
.B(n_105),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1121),
.A2(n_101),
.B(n_182),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1158),
.A2(n_55),
.B(n_59),
.C(n_60),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1112),
.A2(n_133),
.B(n_178),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1193),
.A2(n_63),
.B(n_65),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1218),
.A2(n_63),
.B(n_65),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_R g1378 ( 
.A(n_1213),
.B(n_140),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1151),
.A2(n_127),
.B(n_172),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1116),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1173),
.A2(n_80),
.B(n_159),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1150),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1171),
.B(n_66),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1121),
.A2(n_78),
.B(n_150),
.Y(n_1384)
);

O2A1O1Ixp5_ASAP7_75t_SL g1385 ( 
.A1(n_1187),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1151),
.A2(n_141),
.B(n_146),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1129),
.B(n_185),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1150),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1229),
.B(n_69),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1177),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1168),
.A2(n_1138),
.B(n_1130),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1138),
.B(n_1240),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1194),
.B(n_1215),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1209),
.B(n_1196),
.Y(n_1394)
);

INVx5_ASAP7_75t_L g1395 ( 
.A(n_1213),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1133),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1130),
.Y(n_1397)
);

AO21x1_ASAP7_75t_L g1398 ( 
.A1(n_1172),
.A2(n_1222),
.B(n_1159),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1146),
.A2(n_1235),
.A3(n_1215),
.B(n_1237),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1132),
.B(n_1196),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1172),
.A2(n_1222),
.B(n_1125),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1132),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1132),
.B(n_1196),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1228),
.B(n_1244),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1132),
.A2(n_1196),
.B1(n_1198),
.B2(n_1125),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1235),
.A2(n_1237),
.B1(n_1165),
.B2(n_1205),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1113),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1211),
.B(n_1219),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1168),
.B(n_1133),
.Y(n_1409)
);

NAND3x1_ASAP7_75t_L g1410 ( 
.A(n_1201),
.B(n_1228),
.C(n_1244),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1268),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1383),
.A2(n_1228),
.B1(n_1244),
.B2(n_1145),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1342),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1257),
.Y(n_1414)
);

CKINVDCx16_ASAP7_75t_R g1415 ( 
.A(n_1260),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1262),
.A2(n_1259),
.B(n_1275),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1258),
.B(n_1380),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1290),
.A2(n_1146),
.B(n_1140),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1382),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1255),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_L g1421 ( 
.A(n_1374),
.B(n_1133),
.C(n_1140),
.Y(n_1421)
);

CKINVDCx16_ASAP7_75t_R g1422 ( 
.A(n_1390),
.Y(n_1422)
);

BUFx2_ASAP7_75t_L g1423 ( 
.A(n_1301),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1346),
.B(n_1140),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1324),
.A2(n_1145),
.B1(n_1167),
.B2(n_1397),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1270),
.A2(n_1145),
.B(n_1167),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1306),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1370),
.A2(n_1406),
.B1(n_1286),
.B2(n_1280),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1317),
.A2(n_1331),
.B(n_1332),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1304),
.A2(n_1265),
.B(n_1272),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1261),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1408),
.A2(n_1406),
.B1(n_1338),
.B2(n_1393),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_SL g1433 ( 
.A1(n_1350),
.A2(n_1366),
.B(n_1360),
.C(n_1296),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1294),
.B(n_1273),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_SL g1435 ( 
.A(n_1326),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1346),
.B(n_1407),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1273),
.B(n_1333),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1333),
.B(n_1263),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1368),
.B(n_1360),
.C(n_1366),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1306),
.Y(n_1440)
);

BUFx4_ASAP7_75t_SL g1441 ( 
.A(n_1343),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1267),
.A2(n_1316),
.B(n_1355),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1255),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1271),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1261),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1263),
.B(n_1307),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1321),
.A2(n_1347),
.B(n_1279),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1299),
.B(n_1302),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1287),
.Y(n_1449)
);

OA21x2_ASAP7_75t_L g1450 ( 
.A1(n_1321),
.A2(n_1347),
.B(n_1279),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1346),
.B(n_1276),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1367),
.A2(n_1376),
.B(n_1377),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1289),
.A2(n_1315),
.B1(n_1295),
.B2(n_1264),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1396),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1346),
.B(n_1276),
.Y(n_1455)
);

O2A1O1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1377),
.A2(n_1376),
.B(n_1278),
.C(n_1289),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1356),
.A2(n_1310),
.B(n_1362),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1329),
.A2(n_1330),
.B(n_1344),
.Y(n_1458)
);

AO21x2_ASAP7_75t_L g1459 ( 
.A1(n_1356),
.A2(n_1298),
.B(n_1315),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1308),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1361),
.A2(n_1277),
.B(n_1363),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1291),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1293),
.B(n_1305),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_SL g1464 ( 
.A(n_1342),
.B(n_1325),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1322),
.B(n_1319),
.Y(n_1465)
);

INVx5_ASAP7_75t_L g1466 ( 
.A(n_1395),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1292),
.B(n_1266),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1311),
.A2(n_1372),
.B(n_1364),
.C(n_1373),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1314),
.B(n_1389),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1323),
.A2(n_1330),
.B(n_1369),
.C(n_1335),
.Y(n_1470)
);

AOI21xp33_ASAP7_75t_L g1471 ( 
.A1(n_1320),
.A2(n_1309),
.B(n_1394),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1378),
.Y(n_1472)
);

AOI221xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1369),
.A2(n_1405),
.B1(n_1351),
.B2(n_1354),
.C(n_1384),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1282),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1313),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_1277),
.Y(n_1476)
);

OAI222xp33_ASAP7_75t_L g1477 ( 
.A1(n_1295),
.A2(n_1309),
.B1(n_1352),
.B2(n_1334),
.C1(n_1353),
.C2(n_1348),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1387),
.B(n_1392),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1394),
.A2(n_1391),
.B(n_1337),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1381),
.A2(n_1358),
.B1(n_1341),
.B2(n_1359),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1285),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1365),
.A2(n_1375),
.B(n_1371),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1345),
.A2(n_1386),
.B(n_1379),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1285),
.A2(n_1357),
.B(n_1349),
.Y(n_1484)
);

OAI222xp33_ASAP7_75t_L g1485 ( 
.A1(n_1337),
.A2(n_1340),
.B1(n_1303),
.B2(n_1283),
.C1(n_1284),
.C2(n_1336),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1387),
.A2(n_1340),
.B(n_1300),
.C(n_1328),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1281),
.A2(n_1297),
.B(n_1410),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1312),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1381),
.A2(n_1398),
.B1(n_1300),
.B2(n_1392),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1288),
.B(n_1282),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1312),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1400),
.A2(n_1403),
.B(n_1401),
.Y(n_1492)
);

O2A1O1Ixp5_ASAP7_75t_L g1493 ( 
.A1(n_1404),
.A2(n_1318),
.B(n_1327),
.C(n_1409),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1339),
.A2(n_1395),
.B1(n_1318),
.B2(n_1327),
.Y(n_1494)
);

INVx6_ASAP7_75t_L g1495 ( 
.A(n_1402),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1312),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1399),
.B(n_1385),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1399),
.B(n_1328),
.Y(n_1498)
);

AO21x2_ASAP7_75t_L g1499 ( 
.A1(n_1328),
.A2(n_1300),
.B(n_1399),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1257),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1268),
.Y(n_1501)
);

BUFx2_ASAP7_75t_SL g1502 ( 
.A(n_1268),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1257),
.Y(n_1504)
);

AOI21xp33_ASAP7_75t_L g1505 ( 
.A1(n_1406),
.A2(n_1338),
.B(n_1408),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1306),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1346),
.B(n_1132),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1256),
.Y(n_1508)
);

INVx2_ASAP7_75t_SL g1509 ( 
.A(n_1268),
.Y(n_1509)
);

NOR4xp25_ASAP7_75t_L g1510 ( 
.A(n_1374),
.B(n_1383),
.C(n_1368),
.D(n_1408),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1410),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1256),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1258),
.B(n_1105),
.Y(n_1513)
);

BUFx2_ASAP7_75t_R g1514 ( 
.A(n_1343),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1257),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1383),
.A2(n_1096),
.B(n_931),
.C(n_1115),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1410),
.Y(n_1517)
);

INVxp67_ASAP7_75t_SL g1518 ( 
.A(n_1382),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1262),
.A2(n_1259),
.B(n_1275),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_SL g1522 ( 
.A(n_1408),
.B(n_789),
.C(n_655),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1346),
.B(n_1407),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1290),
.A2(n_1304),
.B(n_1265),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1265),
.A2(n_1388),
.B(n_1382),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1256),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1408),
.A2(n_1383),
.B(n_646),
.Y(n_1527)
);

AOI21xp5_ASAP7_75t_L g1528 ( 
.A1(n_1262),
.A2(n_1259),
.B(n_1275),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1294),
.B(n_1280),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1306),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1268),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1257),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1294),
.B(n_1280),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1268),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1290),
.A2(n_1304),
.B(n_1265),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1261),
.Y(n_1538)
);

OA21x2_ASAP7_75t_L g1539 ( 
.A1(n_1290),
.A2(n_1304),
.B(n_1265),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1257),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1257),
.Y(n_1541)
);

NAND2x1p5_ASAP7_75t_L g1542 ( 
.A(n_1346),
.B(n_1132),
.Y(n_1542)
);

AO31x2_ASAP7_75t_L g1543 ( 
.A1(n_1382),
.A2(n_936),
.A3(n_1231),
.B(n_1388),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1383),
.B(n_1408),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1324),
.A2(n_1096),
.B1(n_1115),
.B2(n_1299),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1268),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1301),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1256),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1301),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1290),
.A2(n_1274),
.B(n_1256),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_SL g1552 ( 
.A1(n_1383),
.A2(n_782),
.B1(n_1156),
.B2(n_1176),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1257),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_SL g1555 ( 
.A1(n_1330),
.A2(n_1360),
.B(n_1398),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_SL g1556 ( 
.A1(n_1338),
.A2(n_1350),
.B(n_923),
.C(n_1406),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1257),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1290),
.A2(n_1269),
.B(n_1256),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1383),
.A2(n_1176),
.B1(n_819),
.B2(n_782),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1383),
.B(n_1374),
.C(n_1408),
.Y(n_1561)
);

OR2x6_ASAP7_75t_L g1562 ( 
.A(n_1275),
.B(n_1295),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1294),
.B(n_1280),
.Y(n_1563)
);

NAND3xp33_ASAP7_75t_L g1564 ( 
.A(n_1383),
.B(n_1374),
.C(n_1408),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1383),
.A2(n_1009),
.B1(n_1408),
.B2(n_1406),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1268),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1257),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1416),
.A2(n_1528),
.B(n_1521),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1454),
.Y(n_1569)
);

AOI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1516),
.A2(n_1456),
.B(n_1556),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1423),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1535),
.Y(n_1572)
);

NOR2xp67_ASAP7_75t_R g1573 ( 
.A(n_1511),
.B(n_1517),
.Y(n_1573)
);

O2A1O1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1565),
.A2(n_1527),
.B(n_1505),
.C(n_1432),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1544),
.B(n_1564),
.C(n_1561),
.Y(n_1575)
);

AOI21x1_ASAP7_75t_SL g1576 ( 
.A1(n_1497),
.A2(n_1469),
.B(n_1490),
.Y(n_1576)
);

AOI21x1_ASAP7_75t_SL g1577 ( 
.A1(n_1498),
.A2(n_1513),
.B(n_1478),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1454),
.B(n_1451),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1446),
.B(n_1434),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1563),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1516),
.A2(n_1556),
.B(n_1433),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1438),
.B(n_1437),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1550),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1468),
.A2(n_1452),
.B(n_1439),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1544),
.A2(n_1510),
.B(n_1522),
.C(n_1433),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1468),
.A2(n_1453),
.B(n_1470),
.C(n_1555),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1474),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1560),
.A2(n_1552),
.B1(n_1428),
.B2(n_1465),
.Y(n_1588)
);

INVxp67_ASAP7_75t_SL g1589 ( 
.A(n_1481),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1448),
.B(n_1444),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1560),
.A2(n_1428),
.B1(n_1465),
.B2(n_1448),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1417),
.B(n_1467),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1453),
.B(n_1447),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1451),
.B(n_1455),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1447),
.B(n_1450),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1449),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1545),
.A2(n_1430),
.B1(n_1474),
.B2(n_1421),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1463),
.B(n_1567),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1447),
.B(n_1450),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1462),
.B(n_1500),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1504),
.B(n_1515),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1533),
.B(n_1540),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1450),
.B(n_1541),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1554),
.B(n_1558),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1545),
.A2(n_1430),
.B1(n_1486),
.B2(n_1422),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1476),
.A2(n_1430),
.B(n_1539),
.Y(n_1606)
);

AOI21x1_ASAP7_75t_SL g1607 ( 
.A1(n_1424),
.A2(n_1481),
.B(n_1415),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1495),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1486),
.A2(n_1412),
.B1(n_1472),
.B2(n_1489),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1473),
.A2(n_1458),
.B(n_1489),
.C(n_1480),
.Y(n_1610)
);

O2A1O1Ixp5_ASAP7_75t_L g1611 ( 
.A1(n_1493),
.A2(n_1471),
.B(n_1494),
.C(n_1511),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1475),
.Y(n_1612)
);

O2A1O1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1464),
.A2(n_1445),
.B(n_1509),
.C(n_1532),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1420),
.B(n_1443),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1429),
.A2(n_1503),
.B(n_1546),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1413),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1499),
.B(n_1562),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1472),
.A2(n_1435),
.B1(n_1425),
.B2(n_1562),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1451),
.B(n_1455),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1419),
.B(n_1499),
.Y(n_1620)
);

AOI21x1_ASAP7_75t_SL g1621 ( 
.A1(n_1424),
.A2(n_1502),
.B(n_1441),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1419),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1435),
.A2(n_1425),
.B1(n_1562),
.B2(n_1514),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1459),
.B(n_1524),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1413),
.Y(n_1625)
);

AOI21x1_ASAP7_75t_SL g1626 ( 
.A1(n_1424),
.A2(n_1441),
.B(n_1491),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1455),
.B(n_1517),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1459),
.B(n_1537),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1536),
.Y(n_1629)
);

OAI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1547),
.A2(n_1480),
.B1(n_1566),
.B2(n_1536),
.Y(n_1630)
);

OA22x2_ASAP7_75t_L g1631 ( 
.A1(n_1436),
.A2(n_1523),
.B1(n_1492),
.B2(n_1487),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1495),
.B(n_1523),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1411),
.A2(n_1501),
.B1(n_1431),
.B2(n_1538),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1479),
.B(n_1518),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1436),
.B(n_1523),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1537),
.A2(n_1477),
.B(n_1485),
.C(n_1491),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1503),
.A2(n_1519),
.B(n_1534),
.Y(n_1637)
);

AOI21x1_ASAP7_75t_SL g1638 ( 
.A1(n_1436),
.A2(n_1418),
.B(n_1482),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1520),
.A2(n_1559),
.B(n_1530),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1525),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1543),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1466),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1431),
.B(n_1538),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1538),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1546),
.A2(n_1557),
.B(n_1553),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1538),
.B(n_1466),
.Y(n_1646)
);

AOI221x1_ASAP7_75t_SL g1647 ( 
.A1(n_1488),
.A2(n_1506),
.B1(n_1531),
.B2(n_1427),
.C(n_1440),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1507),
.A2(n_1542),
.B1(n_1483),
.B2(n_1496),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1484),
.B(n_1426),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1483),
.A2(n_1460),
.B1(n_1427),
.B2(n_1440),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1543),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1483),
.A2(n_1460),
.B1(n_1506),
.B2(n_1531),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1457),
.B(n_1461),
.Y(n_1653)
);

AOI221x1_ASAP7_75t_SL g1654 ( 
.A1(n_1508),
.A2(n_1512),
.B1(n_1526),
.B2(n_1549),
.C(n_1551),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_L g1655 ( 
.A1(n_1457),
.A2(n_1527),
.B(n_1565),
.C(n_1505),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1442),
.A2(n_1527),
.B(n_1565),
.C(n_1505),
.Y(n_1656)
);

NOR2xp67_ASAP7_75t_L g1657 ( 
.A(n_1442),
.B(n_1511),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1446),
.B(n_1434),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1416),
.A2(n_1528),
.B(n_1521),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1414),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1529),
.B(n_1535),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1516),
.A2(n_1565),
.B(n_1456),
.Y(n_1662)
);

OAI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1527),
.A2(n_1565),
.B1(n_1009),
.B2(n_1564),
.C(n_1561),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1414),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1414),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1544),
.A2(n_1527),
.B1(n_1565),
.B2(n_1564),
.Y(n_1666)
);

AND2x4_ASAP7_75t_SL g1667 ( 
.A(n_1547),
.B(n_1268),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1544),
.A2(n_1527),
.B1(n_1565),
.B2(n_1564),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1544),
.B(n_614),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1516),
.A2(n_1565),
.B(n_1456),
.Y(n_1670)
);

AOI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1416),
.A2(n_1528),
.B(n_1521),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1527),
.A2(n_1383),
.B(n_1564),
.C(n_1561),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1529),
.B(n_1535),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1414),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1414),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1529),
.B(n_1535),
.Y(n_1676)
);

BUFx3_ASAP7_75t_L g1677 ( 
.A(n_1547),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1414),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1527),
.A2(n_1565),
.B(n_1505),
.C(n_1383),
.Y(n_1679)
);

AOI21x1_ASAP7_75t_SL g1680 ( 
.A1(n_1497),
.A2(n_1408),
.B(n_899),
.Y(n_1680)
);

CKINVDCx6p67_ASAP7_75t_R g1681 ( 
.A(n_1413),
.Y(n_1681)
);

NOR2xp67_ASAP7_75t_L g1682 ( 
.A(n_1511),
.B(n_1517),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1446),
.B(n_1434),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1529),
.B(n_1535),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1414),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1446),
.B(n_1434),
.Y(n_1686)
);

O2A1O1Ixp33_ASAP7_75t_L g1687 ( 
.A1(n_1565),
.A2(n_1527),
.B(n_1505),
.C(n_1432),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1416),
.A2(n_1528),
.B(n_1521),
.Y(n_1688)
);

OR2x6_ASAP7_75t_L g1689 ( 
.A(n_1568),
.B(n_1659),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1657),
.B(n_1568),
.Y(n_1690)
);

BUFx3_ASAP7_75t_L g1691 ( 
.A(n_1627),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1603),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1659),
.B(n_1671),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1593),
.B(n_1600),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1603),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1612),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1572),
.B(n_1580),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_R g1698 ( 
.A(n_1616),
.B(n_1625),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1602),
.B(n_1604),
.Y(n_1699)
);

BUFx2_ASAP7_75t_SL g1700 ( 
.A(n_1682),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1579),
.B(n_1658),
.Y(n_1701)
);

NOR2xp67_ASAP7_75t_L g1702 ( 
.A(n_1671),
.B(n_1688),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1590),
.B(n_1596),
.Y(n_1703)
);

BUFx12f_ASAP7_75t_L g1704 ( 
.A(n_1677),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1587),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1688),
.A2(n_1606),
.B(n_1645),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1622),
.B(n_1661),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1673),
.B(n_1620),
.Y(n_1708)
);

OA21x2_ASAP7_75t_L g1709 ( 
.A1(n_1606),
.A2(n_1628),
.B(n_1624),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1650),
.A2(n_1652),
.B(n_1628),
.Y(n_1710)
);

INVx1_ASAP7_75t_SL g1711 ( 
.A(n_1667),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1660),
.B(n_1664),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1588),
.A2(n_1591),
.B1(n_1663),
.B2(n_1668),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1569),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1665),
.B(n_1674),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1579),
.B(n_1658),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1649),
.B(n_1635),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1675),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1683),
.B(n_1686),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1678),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1685),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1601),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1676),
.B(n_1684),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1624),
.A2(n_1640),
.B(n_1610),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1641),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1595),
.B(n_1599),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1669),
.B(n_1575),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1651),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1617),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1617),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1683),
.B(n_1686),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1649),
.B(n_1632),
.Y(n_1732)
);

BUFx6f_ASAP7_75t_L g1733 ( 
.A(n_1642),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1592),
.B(n_1582),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1595),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1589),
.B(n_1599),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1605),
.B(n_1583),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1634),
.Y(n_1738)
);

XNOR2x2_ASAP7_75t_L g1739 ( 
.A(n_1663),
.B(n_1666),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1631),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1631),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_L g1742 ( 
.A(n_1672),
.B(n_1687),
.C(n_1574),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1598),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1582),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1653),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1571),
.B(n_1581),
.Y(n_1746)
);

AND2x4_ASAP7_75t_L g1747 ( 
.A(n_1578),
.B(n_1619),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1636),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1636),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1574),
.B(n_1687),
.C(n_1679),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1609),
.A2(n_1630),
.B1(n_1570),
.B2(n_1623),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1597),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1648),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1570),
.A2(n_1581),
.B1(n_1618),
.B2(n_1633),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1584),
.B(n_1670),
.Y(n_1755)
);

INVx2_ASAP7_75t_SL g1756 ( 
.A(n_1608),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1647),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1608),
.B(n_1656),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1662),
.B(n_1629),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1726),
.B(n_1689),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1726),
.B(n_1655),
.Y(n_1761)
);

CKINVDCx20_ASAP7_75t_R g1762 ( 
.A(n_1711),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1689),
.B(n_1615),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_L g1764 ( 
.A(n_1755),
.Y(n_1764)
);

AOI322xp5_ASAP7_75t_L g1765 ( 
.A1(n_1713),
.A2(n_1585),
.A3(n_1586),
.B1(n_1614),
.B2(n_1613),
.C1(n_1680),
.C2(n_1577),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1725),
.Y(n_1766)
);

CKINVDCx20_ASAP7_75t_R g1767 ( 
.A(n_1704),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1733),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1725),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1708),
.B(n_1639),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1691),
.B(n_1717),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1689),
.B(n_1637),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1696),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1696),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1694),
.B(n_1637),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1692),
.B(n_1586),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1692),
.B(n_1585),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1693),
.B(n_1594),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1693),
.B(n_1594),
.Y(n_1780)
);

INVxp67_ASAP7_75t_L g1781 ( 
.A(n_1740),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_SL g1782 ( 
.A(n_1755),
.B(n_1646),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1694),
.B(n_1654),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1695),
.B(n_1573),
.Y(n_1784)
);

OAI33xp33_ASAP7_75t_L g1785 ( 
.A1(n_1742),
.A2(n_1576),
.A3(n_1607),
.B1(n_1681),
.B2(n_1621),
.B3(n_1626),
.Y(n_1785)
);

NOR2x1_ASAP7_75t_L g1786 ( 
.A(n_1700),
.B(n_1644),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1709),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1699),
.B(n_1643),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1699),
.B(n_1611),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1735),
.B(n_1638),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1709),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1736),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1740),
.B(n_1741),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1709),
.Y(n_1794)
);

NAND2xp33_ASAP7_75t_SL g1795 ( 
.A(n_1767),
.B(n_1714),
.Y(n_1795)
);

OAI31xp33_ASAP7_75t_L g1796 ( 
.A1(n_1783),
.A2(n_1742),
.A3(n_1750),
.B(n_1752),
.Y(n_1796)
);

INVx4_ASAP7_75t_L g1797 ( 
.A(n_1764),
.Y(n_1797)
);

CKINVDCx16_ASAP7_75t_R g1798 ( 
.A(n_1762),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1777),
.B(n_1746),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1764),
.A2(n_1750),
.B1(n_1751),
.B2(n_1754),
.Y(n_1800)
);

AO21x2_ASAP7_75t_L g1801 ( 
.A1(n_1787),
.A2(n_1749),
.B(n_1757),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1765),
.B(n_1727),
.C(n_1757),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1778),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1771),
.B(n_1779),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1761),
.A2(n_1748),
.B1(n_1744),
.B2(n_1737),
.C(n_1729),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1777),
.B(n_1746),
.Y(n_1806)
);

OAI33xp33_ASAP7_75t_L g1807 ( 
.A1(n_1761),
.A2(n_1744),
.A3(n_1731),
.B1(n_1719),
.B2(n_1716),
.B3(n_1701),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1778),
.B(n_1723),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1766),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1784),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1760),
.B(n_1723),
.Y(n_1811)
);

INVx4_ASAP7_75t_L g1812 ( 
.A(n_1764),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1789),
.B(n_1703),
.Y(n_1813)
);

NAND4xp25_ASAP7_75t_SL g1814 ( 
.A(n_1765),
.B(n_1783),
.C(n_1760),
.D(n_1739),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1768),
.Y(n_1815)
);

NOR4xp25_ASAP7_75t_SL g1816 ( 
.A(n_1769),
.B(n_1698),
.C(n_1700),
.D(n_1753),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1792),
.B(n_1697),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1793),
.A2(n_1739),
.B1(n_1737),
.B2(n_1753),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1793),
.A2(n_1758),
.B1(n_1730),
.B2(n_1729),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1793),
.A2(n_1730),
.B1(n_1724),
.B2(n_1710),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1781),
.A2(n_1759),
.B1(n_1738),
.B2(n_1743),
.C(n_1702),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1766),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1776),
.B(n_1707),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1772),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1760),
.B(n_1717),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_SL g1826 ( 
.A1(n_1783),
.A2(n_1710),
.B1(n_1724),
.B2(n_1690),
.Y(n_1826)
);

AOI21xp33_ASAP7_75t_L g1827 ( 
.A1(n_1784),
.A2(n_1724),
.B(n_1710),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1790),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1788),
.B(n_1703),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1776),
.B(n_1707),
.Y(n_1830)
);

AOI33xp33_ASAP7_75t_L g1831 ( 
.A1(n_1790),
.A2(n_1721),
.A3(n_1718),
.B1(n_1705),
.B2(n_1715),
.B3(n_1712),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1785),
.A2(n_1690),
.B(n_1706),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1791),
.A2(n_1736),
.B1(n_1722),
.B2(n_1743),
.C(n_1734),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1788),
.B(n_1732),
.Y(n_1834)
);

NAND4xp25_ASAP7_75t_SL g1835 ( 
.A(n_1786),
.B(n_1704),
.C(n_1721),
.D(n_1722),
.Y(n_1835)
);

AND2x6_ASAP7_75t_SL g1836 ( 
.A(n_1771),
.B(n_1747),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1785),
.A2(n_1720),
.B1(n_1715),
.B2(n_1712),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1768),
.Y(n_1838)
);

OAI211xp5_ASAP7_75t_L g1839 ( 
.A1(n_1773),
.A2(n_1706),
.B(n_1756),
.C(n_1745),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1801),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1809),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1828),
.Y(n_1842)
);

AOI21xp33_ASAP7_75t_L g1843 ( 
.A1(n_1796),
.A2(n_1794),
.B(n_1791),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1809),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1836),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1796),
.B(n_1775),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1822),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1836),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1802),
.A2(n_1786),
.B(n_1782),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1824),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1802),
.B(n_1814),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1823),
.B(n_1770),
.Y(n_1854)
);

OA21x2_ASAP7_75t_L g1855 ( 
.A1(n_1832),
.A2(n_1827),
.B(n_1839),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1799),
.B(n_1775),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1811),
.B(n_1780),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1797),
.Y(n_1858)
);

NAND3xp33_ASAP7_75t_SL g1859 ( 
.A(n_1826),
.B(n_1816),
.C(n_1800),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1815),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1823),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_SL g1862 ( 
.A(n_1797),
.B(n_1782),
.Y(n_1862)
);

BUFx2_ASAP7_75t_L g1863 ( 
.A(n_1815),
.Y(n_1863)
);

INVx2_ASAP7_75t_SL g1864 ( 
.A(n_1815),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1830),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1801),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1797),
.B(n_1812),
.Y(n_1867)
);

BUFx2_ASAP7_75t_L g1868 ( 
.A(n_1838),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1838),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1849),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1849),
.Y(n_1871)
);

NAND2x1p5_ASAP7_75t_L g1872 ( 
.A(n_1858),
.B(n_1797),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1853),
.B(n_1798),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1859),
.A2(n_1807),
.B1(n_1801),
.B2(n_1805),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1846),
.B(n_1804),
.Y(n_1875)
);

INVx1_ASAP7_75t_SL g1876 ( 
.A(n_1846),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1846),
.B(n_1804),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1850),
.B(n_1804),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1859),
.B(n_1812),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1849),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1852),
.Y(n_1881)
);

NAND4xp25_ASAP7_75t_L g1882 ( 
.A(n_1853),
.B(n_1795),
.C(n_1831),
.D(n_1763),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1850),
.B(n_1825),
.Y(n_1883)
);

AOI31xp33_ASAP7_75t_L g1884 ( 
.A1(n_1851),
.A2(n_1818),
.A3(n_1806),
.B(n_1810),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1850),
.B(n_1825),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1848),
.B(n_1808),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1841),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1841),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1857),
.B(n_1834),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1848),
.B(n_1813),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1845),
.B(n_1810),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1845),
.B(n_1837),
.Y(n_1892)
);

BUFx2_ASAP7_75t_L g1893 ( 
.A(n_1851),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1857),
.B(n_1834),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1847),
.B(n_1837),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1844),
.Y(n_1896)
);

HB1xp67_ASAP7_75t_L g1897 ( 
.A(n_1847),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1844),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1863),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1856),
.B(n_1829),
.Y(n_1900)
);

AOI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1843),
.A2(n_1833),
.B(n_1816),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1840),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1840),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1855),
.A2(n_1820),
.B1(n_1821),
.B2(n_1819),
.Y(n_1904)
);

NOR3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1867),
.B(n_1798),
.C(n_1835),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1840),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1842),
.B(n_1843),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1861),
.B(n_1817),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1886),
.B(n_1861),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1887),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1893),
.A2(n_1862),
.B1(n_1855),
.B2(n_1812),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1887),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1893),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1888),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1883),
.B(n_1863),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1888),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1883),
.B(n_1863),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1885),
.B(n_1875),
.Y(n_1918)
);

INVx1_ASAP7_75t_SL g1919 ( 
.A(n_1876),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_SL g1920 ( 
.A(n_1905),
.B(n_1868),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1897),
.B(n_1865),
.Y(n_1921)
);

INVx4_ASAP7_75t_L g1922 ( 
.A(n_1899),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1876),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1885),
.B(n_1868),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1896),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1890),
.B(n_1865),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1890),
.B(n_1854),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1896),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1898),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1873),
.B(n_1855),
.Y(n_1930)
);

INVx6_ASAP7_75t_L g1931 ( 
.A(n_1875),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1874),
.B(n_1855),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1879),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1877),
.B(n_1868),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1898),
.Y(n_1935)
);

OAI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1884),
.A2(n_1879),
.B1(n_1904),
.B2(n_1895),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1892),
.B(n_1855),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1899),
.B(n_1855),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1908),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1884),
.A2(n_1862),
.B1(n_1812),
.B2(n_1858),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1870),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1877),
.B(n_1860),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1870),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1902),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1871),
.Y(n_1945)
);

NAND2x2_ASAP7_75t_L g1946 ( 
.A(n_1907),
.B(n_1860),
.Y(n_1946)
);

NAND2x1p5_ASAP7_75t_L g1947 ( 
.A(n_1878),
.B(n_1858),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1941),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1933),
.B(n_1878),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1936),
.A2(n_1840),
.B1(n_1882),
.B2(n_1901),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1922),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1913),
.B(n_1900),
.Y(n_1952)
);

OR2x2_ASAP7_75t_L g1953 ( 
.A(n_1932),
.B(n_1937),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1913),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1943),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1922),
.Y(n_1956)
);

INVx4_ASAP7_75t_L g1957 ( 
.A(n_1922),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1931),
.Y(n_1958)
);

AO21x2_ASAP7_75t_L g1959 ( 
.A1(n_1938),
.A2(n_1906),
.B(n_1902),
.Y(n_1959)
);

INVx1_ASAP7_75t_SL g1960 ( 
.A(n_1919),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1931),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1931),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1945),
.Y(n_1963)
);

NOR2x1p5_ASAP7_75t_L g1964 ( 
.A(n_1930),
.B(n_1858),
.Y(n_1964)
);

BUFx3_ASAP7_75t_L g1965 ( 
.A(n_1923),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1911),
.A2(n_1872),
.B(n_1906),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1918),
.B(n_1889),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1910),
.Y(n_1968)
);

AO21x2_ASAP7_75t_L g1969 ( 
.A1(n_1944),
.A2(n_1906),
.B(n_1902),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1918),
.B(n_1889),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1927),
.B(n_1882),
.Y(n_1971)
);

INVx3_ASAP7_75t_SL g1972 ( 
.A(n_1931),
.Y(n_1972)
);

AND3x2_ASAP7_75t_L g1973 ( 
.A(n_1944),
.B(n_1866),
.C(n_1903),
.Y(n_1973)
);

HB1xp67_ASAP7_75t_L g1974 ( 
.A(n_1912),
.Y(n_1974)
);

AND2x4_ASAP7_75t_L g1975 ( 
.A(n_1942),
.B(n_1903),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1915),
.Y(n_1976)
);

AOI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1950),
.A2(n_1946),
.B1(n_1920),
.B2(n_1940),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1967),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1974),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1960),
.B(n_1915),
.Y(n_1980)
);

AOI221xp5_ASAP7_75t_L g1981 ( 
.A1(n_1950),
.A2(n_1903),
.B1(n_1920),
.B2(n_1866),
.C(n_1909),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1953),
.A2(n_1946),
.B1(n_1942),
.B2(n_1917),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1960),
.B(n_1926),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1971),
.A2(n_1947),
.B1(n_1927),
.B2(n_1924),
.Y(n_1984)
);

NAND3xp33_ASAP7_75t_L g1985 ( 
.A(n_1953),
.B(n_1934),
.C(n_1924),
.Y(n_1985)
);

OAI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1966),
.A2(n_1917),
.B(n_1934),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1960),
.B(n_1939),
.Y(n_1987)
);

AOI322xp5_ASAP7_75t_L g1988 ( 
.A1(n_1949),
.A2(n_1921),
.A3(n_1935),
.B1(n_1929),
.B2(n_1928),
.C1(n_1914),
.C2(n_1925),
.Y(n_1988)
);

AOI221xp5_ASAP7_75t_L g1989 ( 
.A1(n_1953),
.A2(n_1916),
.B1(n_1926),
.B2(n_1891),
.C(n_1881),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1967),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1965),
.B(n_1894),
.Y(n_1991)
);

A2O1A1Ixp33_ASAP7_75t_L g1992 ( 
.A1(n_1971),
.A2(n_1953),
.B(n_1966),
.C(n_1949),
.Y(n_1992)
);

O2A1O1Ixp33_ASAP7_75t_SL g1993 ( 
.A1(n_1971),
.A2(n_1860),
.B(n_1869),
.C(n_1864),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1974),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1965),
.B(n_1976),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1965),
.B(n_1976),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1954),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1954),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1965),
.B(n_1894),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1978),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1990),
.B(n_1976),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1996),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1991),
.B(n_1949),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1997),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1999),
.B(n_1949),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1980),
.B(n_1972),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1988),
.B(n_1954),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1983),
.B(n_1976),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1987),
.B(n_1958),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1995),
.B(n_1971),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1998),
.B(n_1958),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1988),
.B(n_1954),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1979),
.Y(n_2013)
);

AOI221xp5_ASAP7_75t_SL g2014 ( 
.A1(n_2007),
.A2(n_1992),
.B1(n_1981),
.B2(n_1986),
.C(n_1984),
.Y(n_2014)
);

AOI221xp5_ASAP7_75t_L g2015 ( 
.A1(n_2007),
.A2(n_1989),
.B1(n_1985),
.B2(n_1977),
.C(n_1994),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_2009),
.B(n_1982),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_2012),
.A2(n_1993),
.B(n_1966),
.Y(n_2017)
);

AOI221xp5_ASAP7_75t_L g2018 ( 
.A1(n_2012),
.A2(n_2010),
.B1(n_2002),
.B2(n_2005),
.C(n_2013),
.Y(n_2018)
);

NOR3xp33_ASAP7_75t_L g2019 ( 
.A(n_2006),
.B(n_1961),
.C(n_1958),
.Y(n_2019)
);

NOR3xp33_ASAP7_75t_L g2020 ( 
.A(n_2011),
.B(n_1961),
.C(n_1958),
.Y(n_2020)
);

OAI22xp33_ASAP7_75t_L g2021 ( 
.A1(n_2008),
.A2(n_1972),
.B1(n_1961),
.B2(n_1962),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_2001),
.A2(n_1972),
.B1(n_1962),
.B2(n_1961),
.Y(n_2022)
);

AOI211xp5_ASAP7_75t_L g2023 ( 
.A1(n_2003),
.A2(n_1972),
.B(n_1966),
.C(n_1962),
.Y(n_2023)
);

AOI221xp5_ASAP7_75t_L g2024 ( 
.A1(n_2004),
.A2(n_1959),
.B1(n_1952),
.B2(n_1968),
.C(n_1955),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2020),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_2015),
.A2(n_1962),
.B1(n_1972),
.B2(n_2000),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_2022),
.Y(n_2027)
);

NOR4xp25_ASAP7_75t_L g2028 ( 
.A(n_2018),
.B(n_1956),
.C(n_1951),
.D(n_1968),
.Y(n_2028)
);

NOR4xp25_ASAP7_75t_SL g2029 ( 
.A(n_2016),
.B(n_1968),
.C(n_1948),
.D(n_1955),
.Y(n_2029)
);

AOI221xp5_ASAP7_75t_SL g2030 ( 
.A1(n_2017),
.A2(n_2023),
.B1(n_2021),
.B2(n_2024),
.C(n_1951),
.Y(n_2030)
);

OAI322xp33_ASAP7_75t_L g2031 ( 
.A1(n_2014),
.A2(n_1951),
.A3(n_1956),
.B1(n_1948),
.B2(n_1963),
.C1(n_1955),
.C2(n_1952),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_2027),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_2025),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_2031),
.B(n_1951),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2029),
.B(n_1967),
.Y(n_2035)
);

XNOR2xp5_ASAP7_75t_L g2036 ( 
.A(n_2026),
.B(n_2019),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2030),
.B(n_1967),
.Y(n_2037)
);

XNOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2028),
.B(n_1964),
.Y(n_2038)
);

OAI21xp5_ASAP7_75t_SL g2039 ( 
.A1(n_2025),
.A2(n_1956),
.B(n_1973),
.Y(n_2039)
);

AND2x2_ASAP7_75t_SL g2040 ( 
.A(n_2035),
.B(n_1957),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_2037),
.A2(n_1959),
.B1(n_1964),
.B2(n_1969),
.Y(n_2041)
);

OAI321xp33_ASAP7_75t_L g2042 ( 
.A1(n_2034),
.A2(n_2033),
.A3(n_2038),
.B1(n_1956),
.B2(n_2039),
.C(n_2036),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_2032),
.Y(n_2043)
);

NAND4xp25_ASAP7_75t_SL g2044 ( 
.A(n_2039),
.B(n_1970),
.C(n_1948),
.D(n_1963),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2035),
.B(n_1970),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_2043),
.Y(n_2046)
);

OAI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_2045),
.A2(n_1963),
.B1(n_1947),
.B2(n_1957),
.Y(n_2047)
);

NOR2x1_ASAP7_75t_L g2048 ( 
.A(n_2044),
.B(n_1957),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_2040),
.Y(n_2049)
);

NAND2x1_ASAP7_75t_L g2050 ( 
.A(n_2046),
.B(n_1957),
.Y(n_2050)
);

OAI221xp5_ASAP7_75t_L g2051 ( 
.A1(n_2049),
.A2(n_2041),
.B1(n_2042),
.B2(n_1957),
.C(n_1872),
.Y(n_2051)
);

OAI211xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2051),
.A2(n_2048),
.B(n_2047),
.C(n_1957),
.Y(n_2052)
);

AOI322xp5_ASAP7_75t_L g2053 ( 
.A1(n_2050),
.A2(n_1975),
.A3(n_1973),
.B1(n_1959),
.B2(n_1969),
.C1(n_1964),
.C2(n_1970),
.Y(n_2053)
);

OAI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_2053),
.A2(n_1975),
.B(n_1970),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2052),
.Y(n_2055)
);

NAND3xp33_ASAP7_75t_L g2056 ( 
.A(n_2055),
.B(n_1975),
.C(n_1959),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2054),
.B(n_1959),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_2057),
.Y(n_2058)
);

XOR2xp5_ASAP7_75t_L g2059 ( 
.A(n_2056),
.B(n_1975),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_2059),
.A2(n_1959),
.B1(n_1969),
.B2(n_1975),
.Y(n_2060)
);

AOI21xp5_ASAP7_75t_SL g2061 ( 
.A1(n_2060),
.A2(n_2058),
.B(n_1975),
.Y(n_2061)
);

OAI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2061),
.A2(n_1969),
.B(n_1872),
.Y(n_2062)
);

INVxp67_ASAP7_75t_L g2063 ( 
.A(n_2062),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2063),
.A2(n_1969),
.B1(n_1880),
.B2(n_1871),
.Y(n_2064)
);

AOI211xp5_ASAP7_75t_L g2065 ( 
.A1(n_2064),
.A2(n_1969),
.B(n_1867),
.C(n_1864),
.Y(n_2065)
);


endmodule