module real_jpeg_25859_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_1),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_1),
.B(n_73),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_1),
.B(n_28),
.C(n_40),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_162),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_1),
.B(n_86),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_1),
.A2(n_25),
.B1(n_31),
.B2(n_236),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_59),
.B1(n_60),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_80),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_80),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_3),
.A2(n_49),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_5),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_5),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_7),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_119),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_119),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_119),
.Y(n_259)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_9),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_166),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_166),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_166),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_14),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_158),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_158),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_158),
.Y(n_229)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_140),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_121),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_20),
.B(n_121),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_96),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_21),
.A2(n_75),
.B1(n_76),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_21),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_50),
.B2(n_74),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_22),
.A2(n_51),
.B(n_53),
.Y(n_138)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_24),
.A2(n_34),
.B1(n_51),
.B2(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_25),
.A2(n_148),
.B(n_150),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_25),
.A2(n_101),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_25),
.A2(n_229),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_25),
.A2(n_32),
.B(n_150),
.Y(n_254)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_26),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_26),
.A2(n_149),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_26),
.A2(n_196),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_241),
.Y(n_240)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_29),
.Y(n_184)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_30),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_43),
.B(n_46),
.Y(n_34)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_35),
.A2(n_42),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_35),
.A2(n_42),
.B1(n_215),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_35),
.A2(n_89),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_38),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_37),
.A2(n_84),
.B(n_250),
.C(n_252),
.Y(n_249)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_38),
.B(n_211),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_L g252 ( 
.A(n_38),
.B(n_59),
.C(n_83),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_42),
.A2(n_92),
.B(n_109),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_42),
.B(n_162),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_44),
.A2(n_91),
.B1(n_93),
.B2(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_90),
.B(n_93),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_67),
.B(n_69),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_54),
.A2(n_117),
.B(n_120),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_54),
.A2(n_56),
.B1(n_165),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_55),
.B(n_70),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_55),
.A2(n_73),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_55),
.A2(n_73),
.B1(n_118),
.B2(n_172),
.Y(n_291)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_57),
.A2(n_60),
.B(n_163),
.C(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_58),
.B(n_59),
.C(n_66),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_60),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g251 ( 
.A(n_60),
.B(n_162),
.CON(n_251),
.SN(n_251)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_66),
.A2(n_162),
.B(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_73),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_71),
.B(n_162),
.Y(n_163)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_88),
.B(n_95),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_88),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_85),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_81),
.A2(n_87),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_86),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_81),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_81),
.A2(n_86),
.B1(n_201),
.B2(n_251),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_81),
.A2(n_135),
.B(n_177),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_85),
.B(n_114),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_85),
.A2(n_175),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_86),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_90),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_91),
.A2(n_93),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_91),
.A2(n_93),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_123),
.B1(n_136),
.B2(n_137),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_96),
.A2(n_97),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_110),
.C(n_115),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_98),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_99),
.A2(n_100),
.B1(n_106),
.B2(n_107),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_104),
.A2(n_182),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_105),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_302)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_138),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_307),
.B(n_313),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_295),
.B(n_306),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_203),
.B(n_283),
.C(n_294),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_188),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_144),
.B(n_188),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_167),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_146),
.B(n_154),
.C(n_167),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_153),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_147),
.B(n_153),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_151),
.Y(n_237)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_152),
.B(n_162),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_160),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_178),
.B2(n_187),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_170),
.B(n_173),
.C(n_187),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_180),
.B1(n_185),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_189),
.B(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_191),
.B(n_193),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_282),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_277),
.B(n_281),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_262),
.B(n_276),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_245),
.B(n_261),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_225),
.B(n_244),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_216),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_212),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_220),
.C(n_223),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_243),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_231),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_238),
.B(n_242),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_260),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_260),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_255),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_256),
.C(n_257),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_272),
.C(n_274),
.Y(n_280)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_280),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_285),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_288),
.C(n_293),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_291),
.C(n_292),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_297),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_305),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_304),
.C(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_301),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_310),
.Y(n_312)
);


endmodule