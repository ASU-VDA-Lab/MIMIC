module real_jpeg_13042_n_17 (n_338, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_338;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_2),
.A2(n_53),
.B1(n_54),
.B2(n_62),
.Y(n_265)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_4),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_76),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_76),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_4),
.A2(n_63),
.B1(n_65),
.B2(n_76),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_6),
.A2(n_34),
.B1(n_53),
.B2(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_6),
.A2(n_34),
.B1(n_63),
.B2(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_7),
.A2(n_38),
.B1(n_63),
.B2(n_65),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_7),
.A2(n_38),
.B1(n_53),
.B2(n_54),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_8),
.A2(n_53),
.B1(n_54),
.B2(n_133),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_8),
.A2(n_63),
.B1(n_65),
.B2(n_133),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_133),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_10),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_10),
.A2(n_63),
.B1(n_65),
.B2(n_80),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_10),
.A2(n_53),
.B1(n_54),
.B2(n_80),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_80),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_11),
.A2(n_63),
.B1(n_65),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_11),
.B(n_54),
.C(n_68),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_11),
.B(n_89),
.Y(n_169)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_11),
.A2(n_124),
.B(n_177),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_23),
.B(n_88),
.C(n_204),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_161),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_11),
.B(n_21),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_11),
.B(n_30),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_12),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_13),
.A2(n_63),
.B1(n_65),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_13),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_173),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_13),
.A2(n_23),
.B1(n_24),
.B2(n_173),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_173),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_63),
.B1(n_65),
.B2(n_91),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_91),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_15),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_15),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_15),
.B(n_24),
.Y(n_261)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_21),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_21),
.A2(n_27),
.B1(n_37),
.B2(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_22),
.A2(n_75),
.B(n_77),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_22),
.A2(n_28),
.B1(n_75),
.B2(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_22),
.B(n_79),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_22),
.A2(n_28),
.B1(n_100),
.B2(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_22),
.A2(n_77),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_22),
.A2(n_28),
.B1(n_132),
.B2(n_275),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_23),
.A2(n_24),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

AOI32xp33_ASAP7_75t_L g260 ( 
.A1(n_23),
.A2(n_26),
.A3(n_31),
.B1(n_248),
.B2(n_261),
.Y(n_260)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_27),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_28),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_28),
.A2(n_31),
.B(n_161),
.C(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_35),
.B(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_36),
.B(n_333),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_332),
.B(n_334),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_320),
.B(n_331),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_149),
.B(n_317),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_136),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_111),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_46),
.B(n_111),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_81),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_47),
.B(n_82),
.C(n_97),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B(n_74),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_48),
.A2(n_49),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_59),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_50),
.A2(n_51),
.B1(n_74),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_50),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_57),
.Y(n_51)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_52),
.A2(n_56),
.B1(n_182),
.B2(n_184),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_52),
.B(n_178),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_52),
.A2(n_56),
.B1(n_123),
.B2(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_53),
.B(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_56),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_56),
.B(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_71),
.B2(n_73),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_61),
.A2(n_66),
.B1(n_73),
.B2(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_65),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g89 ( 
.A1(n_63),
.A2(n_65),
.B1(n_87),
.B2(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_63),
.B(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_65),
.A2(n_87),
.B(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_66),
.A2(n_73),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_66),
.B(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_66),
.A2(n_73),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_66),
.A2(n_73),
.B1(n_128),
.B2(n_254),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_68),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_72),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_70),
.A2(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_70),
.B(n_161),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_70),
.A2(n_174),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_73),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_97),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_83),
.B(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_94),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_90),
.B1(n_92),
.B2(n_93),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_84),
.A2(n_90),
.B1(n_92),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_84),
.A2(n_92),
.B1(n_105),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_84),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_84),
.A2(n_92),
.B1(n_224),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_84),
.A2(n_210),
.B(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_89),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_85),
.B(n_211),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_85),
.A2(n_89),
.B(n_324),
.Y(n_323)
);

NOR2x1_ASAP7_75t_R g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_92),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_92),
.A2(n_130),
.B(n_225),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_160),
.B(n_162),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_95),
.A2(n_162),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_110),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_99),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_99),
.B(n_102),
.C(n_107),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_99),
.B(n_140),
.C(n_147),
.Y(n_330)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_109),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_107),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_107),
.B(n_141),
.C(n_145),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.C(n_118),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_112),
.A2(n_113),
.B1(n_117),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_117),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_118),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_131),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_119),
.A2(n_120),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_121),
.A2(n_126),
.B1(n_127),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_121),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_124),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_124),
.A2(n_125),
.B1(n_206),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_124),
.A2(n_125),
.B1(n_231),
.B2(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_125),
.A2(n_183),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_161),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_125),
.A2(n_191),
.B(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_129),
.B(n_131),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_135),
.B(n_246),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g317 ( 
.A1(n_136),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_148),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_137),
.B(n_148),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_147),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_142),
.Y(n_326)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_146),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_311),
.B(n_316),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_299),
.B(n_310),
.Y(n_150)
);

OAI321xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_267),
.A3(n_292),
.B1(n_297),
.B2(n_298),
.C(n_338),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_240),
.B(n_266),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_218),
.B(n_239),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_199),
.B(n_217),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_179),
.B(n_198),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_166),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_157),
.B(n_166),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_164),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_171),
.C(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_176),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_187),
.B(n_197),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_181),
.B(n_185),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_192),
.B(n_196),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_212),
.C(n_216),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_214),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_220),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_232),
.B2(n_233),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_235),
.C(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_227),
.C(n_230),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_241),
.B(n_242),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_256),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_243),
.B(n_257),
.C(n_258),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_249),
.B2(n_255),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_244),
.B(n_250),
.C(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_282),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_282),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_278),
.C(n_281),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_269),
.A2(n_270),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_272),
.B(n_276),
.C(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_281),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_280),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_291),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_284),
.B(n_286),
.C(n_291),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_290),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_309),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_304),
.C(n_305),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_330),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_330),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_323),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_325),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_327),
.C(n_329),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_333),
.Y(n_336)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);


endmodule