module fake_jpeg_18318_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_67;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_24),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_2),
.Y(n_39)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_20),
.B1(n_15),
.B2(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_20),
.B1(n_15),
.B2(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_21),
.A2(n_25),
.B1(n_13),
.B2(n_24),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_16),
.C(n_3),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_5),
.B(n_6),
.Y(n_49)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_28),
.Y(n_46)
);

NOR3xp33_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_29),
.C(n_31),
.Y(n_51)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_36),
.B(n_33),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_26),
.C(n_7),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_42),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.C(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_44),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_61),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_48),
.C(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_55),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g64 ( 
.A(n_60),
.B(n_46),
.Y(n_64)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_65),
.A3(n_67),
.B1(n_62),
.B2(n_43),
.C1(n_56),
.C2(n_26),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_69),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_43),
.Y(n_69)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_70),
.A2(n_41),
.B(n_45),
.Y(n_71)
);


endmodule