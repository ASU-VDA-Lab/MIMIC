module real_aes_15795_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_1252;
wire n_430;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_340;
wire n_483;
wire n_1280;
wire n_1352;
wire n_394;
wire n_1323;
wire n_729;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_0), .A2(n_6), .B1(n_267), .B2(n_270), .Y(n_266) );
OAI22xp33_ASAP7_75t_SL g929 ( .A1(n_1), .A2(n_114), .B1(n_789), .B2(n_841), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g942 ( .A1(n_1), .A2(n_27), .B1(n_533), .B2(n_554), .Y(n_942) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_2), .A2(n_28), .B1(n_571), .B2(n_582), .Y(n_970) );
OAI22xp5_ASAP7_75t_SL g978 ( .A1(n_2), .A2(n_117), .B1(n_533), .B2(n_556), .Y(n_978) );
AOI22xp33_ASAP7_75t_SL g1150 ( .A1(n_3), .A2(n_7), .B1(n_616), .B2(n_1151), .Y(n_1150) );
AOI22xp33_ASAP7_75t_SL g1188 ( .A1(n_3), .A2(n_213), .B1(n_1072), .B2(n_1189), .Y(n_1188) );
INVx1_ASAP7_75t_L g858 ( .A(n_4), .Y(n_858) );
INVx1_ASAP7_75t_L g1075 ( .A(n_5), .Y(n_1075) );
AOI22xp33_ASAP7_75t_L g1192 ( .A1(n_7), .A2(n_217), .B1(n_520), .B2(n_1189), .Y(n_1192) );
AOI22xp33_ASAP7_75t_SL g1279 ( .A1(n_8), .A2(n_234), .B1(n_621), .B2(n_1280), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_8), .A2(n_160), .B1(n_505), .B2(n_1289), .Y(n_1288) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_9), .A2(n_645), .B(n_649), .C(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g664 ( .A(n_9), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g973 ( .A(n_10), .Y(n_973) );
INVx1_ASAP7_75t_L g1058 ( .A(n_11), .Y(n_1058) );
INVx1_ASAP7_75t_L g1333 ( .A(n_12), .Y(n_1333) );
OAI22xp33_ASAP7_75t_L g1374 ( .A1(n_12), .A2(n_83), .B1(n_1375), .B2(n_1378), .Y(n_1374) );
AOI22xp33_ASAP7_75t_SL g1273 ( .A1(n_13), .A2(n_214), .B1(n_621), .B2(n_1274), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_13), .A2(n_196), .B1(n_488), .B2(n_1241), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_14), .Y(n_949) );
INVx1_ASAP7_75t_L g465 ( .A(n_15), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_15), .B(n_475), .Y(n_614) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_15), .B(n_576), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_15), .B(n_201), .Y(n_1311) );
OAI22xp33_ASAP7_75t_L g774 ( .A1(n_16), .A2(n_185), .B1(n_467), .B2(n_657), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_16), .A2(n_185), .B1(n_796), .B2(n_798), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_17), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g887 ( .A(n_18), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g896 ( .A(n_19), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_20), .A2(n_208), .B1(n_621), .B2(n_1017), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_20), .A2(n_61), .B1(n_523), .B2(n_1037), .Y(n_1036) );
OAI222xp33_ASAP7_75t_L g992 ( .A1(n_21), .A2(n_188), .B1(n_572), .B2(n_925), .C1(n_993), .C2(n_994), .Y(n_992) );
OAI222xp33_ASAP7_75t_L g1023 ( .A1(n_21), .A2(n_129), .B1(n_188), .B2(n_1024), .C1(n_1025), .C2(n_1026), .Y(n_1023) );
INVx1_ASAP7_75t_L g670 ( .A(n_22), .Y(n_670) );
INVx2_ASAP7_75t_L g263 ( .A(n_23), .Y(n_263) );
AND2x2_ASAP7_75t_L g265 ( .A(n_23), .B(n_106), .Y(n_265) );
AND2x2_ASAP7_75t_L g271 ( .A(n_23), .B(n_269), .Y(n_271) );
INVx1_ASAP7_75t_L g549 ( .A(n_24), .Y(n_549) );
OAI211xp5_ASAP7_75t_L g1098 ( .A1(n_25), .A2(n_542), .B(n_756), .C(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1108 ( .A(n_25), .Y(n_1108) );
INVx1_ASAP7_75t_L g1173 ( .A(n_26), .Y(n_1173) );
OAI22xp33_ASAP7_75t_SL g926 ( .A1(n_27), .A2(n_216), .B1(n_571), .B2(n_927), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_28), .B(n_535), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_29), .A2(n_194), .B1(n_533), .B2(n_1077), .Y(n_1076) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_29), .A2(n_244), .B1(n_571), .B2(n_657), .Y(n_1088) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_30), .A2(n_206), .B1(n_267), .B2(n_270), .Y(n_288) );
INVx1_ASAP7_75t_L g1117 ( .A(n_31), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1250 ( .A1(n_32), .A2(n_1251), .B1(n_1252), .B2(n_1254), .Y(n_1250) );
CKINVDCx5p33_ASAP7_75t_R g1251 ( .A(n_32), .Y(n_1251) );
INVx1_ASAP7_75t_L g1008 ( .A(n_33), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_33), .A2(n_208), .B1(n_493), .B2(n_1037), .Y(n_1043) );
XOR2xp5_ASAP7_75t_L g882 ( .A(n_34), .B(n_883), .Y(n_882) );
XNOR2x2_ASAP7_75t_SL g1094 ( .A(n_35), .B(n_1095), .Y(n_1094) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_36), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_37), .A2(n_105), .B1(n_1348), .B2(n_1352), .Y(n_1347) );
INVx1_ASAP7_75t_L g1170 ( .A(n_38), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_38), .A2(n_168), .B1(n_980), .B2(n_1025), .Y(n_1178) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_39), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_40), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_41), .A2(n_238), .B1(n_259), .B2(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g1101 ( .A(n_42), .Y(n_1101) );
OAI211xp5_ASAP7_75t_L g1105 ( .A1(n_42), .A2(n_687), .B(n_1106), .C(n_1107), .Y(n_1105) );
INVx1_ASAP7_75t_L g848 ( .A(n_43), .Y(n_848) );
INVx1_ASAP7_75t_L g1201 ( .A(n_44), .Y(n_1201) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_45), .A2(n_86), .B1(n_621), .B2(n_1232), .Y(n_1231) );
AOI22xp33_ASAP7_75t_SL g1245 ( .A1(n_45), .A2(n_224), .B1(n_520), .B2(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1312 ( .A(n_46), .Y(n_1312) );
INVx1_ASAP7_75t_L g1174 ( .A(n_47), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g643 ( .A1(n_48), .A2(n_116), .B1(n_581), .B2(n_582), .Y(n_643) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_48), .A2(n_58), .B1(n_554), .B2(n_556), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_49), .A2(n_219), .B1(n_267), .B2(n_270), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_50), .Y(n_957) );
AO22x1_ASAP7_75t_L g285 ( .A1(n_51), .A2(n_65), .B1(n_259), .B2(n_264), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_52), .A2(n_247), .B1(n_533), .B2(n_535), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_52), .A2(n_53), .B1(n_581), .B2(n_582), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_53), .A2(n_154), .B1(n_554), .B2(n_556), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_54), .A2(n_131), .B1(n_1025), .B2(n_1208), .Y(n_1207) );
INVxp67_ASAP7_75t_SL g1220 ( .A(n_54), .Y(n_1220) );
INVx1_ASAP7_75t_L g1258 ( .A(n_55), .Y(n_1258) );
INVx1_ASAP7_75t_L g491 ( .A(n_56), .Y(n_491) );
INVx1_ASAP7_75t_L g499 ( .A(n_56), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_57), .A2(n_124), .B1(n_796), .B2(n_820), .Y(n_819) );
OAI22xp33_ASAP7_75t_L g840 ( .A1(n_57), .A2(n_124), .B1(n_467), .B2(n_841), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_58), .A2(n_182), .B1(n_571), .B2(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g748 ( .A(n_59), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_60), .Y(n_951) );
INVx1_ASAP7_75t_L g1009 ( .A(n_61), .Y(n_1009) );
XOR2xp5_ASAP7_75t_L g1044 ( .A(n_62), .B(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g732 ( .A(n_63), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_64), .A2(n_85), .B1(n_616), .B2(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1187 ( .A(n_64), .Y(n_1187) );
INVx1_ASAP7_75t_L g261 ( .A(n_66), .Y(n_261) );
XOR2x2_ASAP7_75t_L g1197 ( .A(n_67), .B(n_1198), .Y(n_1197) );
INVx2_ASAP7_75t_L g514 ( .A(n_68), .Y(n_514) );
XNOR2x2_ASAP7_75t_L g720 ( .A(n_69), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_70), .A2(n_220), .B1(n_488), .B2(n_493), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_70), .A2(n_159), .B1(n_624), .B2(n_626), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_71), .A2(n_200), .B1(n_788), .B2(n_790), .Y(n_787) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_71), .A2(n_200), .B1(n_810), .B2(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g1050 ( .A(n_72), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1205 ( .A(n_73), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_73), .A2(n_131), .B1(n_783), .B2(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g545 ( .A(n_74), .Y(n_545) );
INVx1_ASAP7_75t_L g654 ( .A(n_75), .Y(n_654) );
INVx1_ASAP7_75t_L g539 ( .A(n_76), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_77), .A2(n_157), .B1(n_259), .B2(n_264), .Y(n_282) );
INVx1_ASAP7_75t_L g1127 ( .A(n_78), .Y(n_1127) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_79), .A2(n_177), .B1(n_1171), .B2(n_1323), .C(n_1324), .Y(n_1322) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_79), .A2(n_123), .B1(n_1037), .B2(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g734 ( .A(n_80), .Y(n_734) );
INVx1_ASAP7_75t_L g678 ( .A(n_81), .Y(n_678) );
AO221x2_ASAP7_75t_L g352 ( .A1(n_82), .A2(n_192), .B1(n_267), .B2(n_270), .C(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g1329 ( .A(n_83), .Y(n_1329) );
INVx1_ASAP7_75t_L g1163 ( .A(n_84), .Y(n_1163) );
INVxp67_ASAP7_75t_SL g1191 ( .A(n_85), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_86), .A2(n_94), .B1(n_520), .B2(n_1241), .Y(n_1240) );
XOR2xp5_ASAP7_75t_L g984 ( .A(n_87), .B(n_985), .Y(n_984) );
AOI221xp5_ASAP7_75t_L g500 ( .A1(n_88), .A2(n_245), .B1(n_501), .B2(n_505), .C(n_510), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_88), .A2(n_121), .B1(n_632), .B2(n_635), .Y(n_631) );
AOI21xp33_ASAP7_75t_L g1315 ( .A1(n_89), .A2(n_1276), .B(n_1316), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_89), .A2(n_151), .B1(n_1126), .B2(n_1239), .Y(n_1369) );
INVx1_ASAP7_75t_L g922 ( .A(n_90), .Y(n_922) );
OAI211xp5_ASAP7_75t_SL g933 ( .A1(n_90), .A2(n_802), .B(n_934), .C(n_936), .Y(n_933) );
INVx1_ASAP7_75t_L g1263 ( .A(n_91), .Y(n_1263) );
OAI221xp5_ASAP7_75t_L g1268 ( .A1(n_91), .A2(n_225), .B1(n_889), .B2(n_1269), .C(n_1270), .Y(n_1268) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_92), .A2(n_138), .B1(n_581), .B2(n_582), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_92), .A2(n_138), .B1(n_535), .B2(n_556), .Y(n_1267) );
INVx1_ASAP7_75t_L g1168 ( .A(n_93), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_94), .A2(n_224), .B1(n_624), .B2(n_1230), .Y(n_1235) );
OAI211xp5_ASAP7_75t_L g1302 ( .A1(n_95), .A2(n_1303), .B(n_1308), .C(n_1313), .Y(n_1302) );
INVx1_ASAP7_75t_L g1362 ( .A(n_95), .Y(n_1362) );
INVx1_ASAP7_75t_L g726 ( .A(n_96), .Y(n_726) );
OAI211xp5_ASAP7_75t_L g775 ( .A1(n_97), .A2(n_776), .B(n_779), .C(n_785), .Y(n_775) );
INVx1_ASAP7_75t_L g808 ( .A(n_97), .Y(n_808) );
OAI221xp5_ASAP7_75t_L g1070 ( .A1(n_98), .A2(n_244), .B1(n_535), .B2(n_554), .C(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1086 ( .A(n_98), .Y(n_1086) );
INVx1_ASAP7_75t_L g854 ( .A(n_99), .Y(n_854) );
AND2x2_ASAP7_75t_L g260 ( .A(n_100), .B(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_100), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g987 ( .A1(n_101), .A2(n_988), .B(n_989), .C(n_998), .Y(n_987) );
INVx1_ASAP7_75t_L g1030 ( .A(n_101), .Y(n_1030) );
INVx1_ASAP7_75t_L g1052 ( .A(n_102), .Y(n_1052) );
INVx1_ASAP7_75t_L g1124 ( .A(n_103), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g1278 ( .A1(n_104), .A2(n_196), .B1(n_991), .B2(n_1276), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_104), .A2(n_214), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
OAI211xp5_ASAP7_75t_SL g1318 ( .A1(n_105), .A2(n_1319), .B(n_1321), .C(n_1328), .Y(n_1318) );
AND2x2_ASAP7_75t_L g262 ( .A(n_106), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g269 ( .A(n_106), .Y(n_269) );
INVx1_ASAP7_75t_L g1053 ( .A(n_107), .Y(n_1053) );
INVx1_ASAP7_75t_L g1210 ( .A(n_108), .Y(n_1210) );
INVx2_ASAP7_75t_L g512 ( .A(n_109), .Y(n_512) );
INVx1_ASAP7_75t_L g529 ( .A(n_109), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_109), .B(n_514), .Y(n_1342) );
INVx1_ASAP7_75t_L g686 ( .A(n_110), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_111), .A2(n_190), .B1(n_259), .B2(n_264), .Y(n_258) );
INVx1_ASAP7_75t_L g1120 ( .A(n_112), .Y(n_1120) );
AOI22xp33_ASAP7_75t_SL g1236 ( .A1(n_113), .A2(n_236), .B1(n_621), .B2(n_1232), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_113), .A2(n_165), .B1(n_1035), .B2(n_1239), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_114), .A2(n_216), .B1(n_535), .B2(n_556), .Y(n_932) );
OAI22xp33_ASAP7_75t_SL g975 ( .A1(n_115), .A2(n_117), .B1(n_581), .B2(n_657), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_115), .A2(n_120), .B1(n_939), .B2(n_940), .Y(n_982) );
OAI22xp5_ASAP7_75t_SL g659 ( .A1(n_116), .A2(n_182), .B1(n_533), .B2(n_535), .Y(n_659) );
INVx1_ASAP7_75t_L g863 ( .A(n_118), .Y(n_863) );
INVx1_ASAP7_75t_L g691 ( .A(n_119), .Y(n_691) );
INVx1_ASAP7_75t_L g974 ( .A(n_120), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_121), .A2(n_195), .B1(n_501), .B2(n_505), .C(n_518), .Y(n_517) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_122), .A2(n_211), .B1(n_533), .B2(n_1103), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1112 ( .A1(n_122), .A2(n_211), .B1(n_571), .B2(n_841), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_123), .A2(n_183), .B1(n_621), .B2(n_1232), .Y(n_1317) );
INVx1_ASAP7_75t_L g1133 ( .A(n_125), .Y(n_1133) );
INVx1_ASAP7_75t_L g997 ( .A(n_126), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1027 ( .A1(n_126), .A2(n_199), .B1(n_535), .B2(n_556), .Y(n_1027) );
INVx1_ASAP7_75t_L g688 ( .A(n_127), .Y(n_688) );
AO22x1_ASAP7_75t_L g286 ( .A1(n_128), .A2(n_204), .B1(n_267), .B2(n_270), .Y(n_286) );
AOI31xp33_ASAP7_75t_L g485 ( .A1(n_128), .A2(n_486), .A3(n_531), .B(n_567), .Y(n_485) );
NAND2xp33_ASAP7_75t_SL g609 ( .A(n_128), .B(n_610), .Y(n_609) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_128), .Y(n_638) );
INVx1_ASAP7_75t_L g990 ( .A(n_129), .Y(n_990) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_130), .Y(n_1011) );
BUFx3_ASAP7_75t_L g492 ( .A(n_132), .Y(n_492) );
OAI211xp5_ASAP7_75t_SL g971 ( .A1(n_133), .A2(n_649), .B(n_920), .C(n_972), .Y(n_971) );
OAI211xp5_ASAP7_75t_SL g979 ( .A1(n_133), .A2(n_802), .B(n_980), .C(n_981), .Y(n_979) );
INVx1_ASAP7_75t_L g1149 ( .A(n_134), .Y(n_1149) );
INVx1_ASAP7_75t_L g676 ( .A(n_135), .Y(n_676) );
INVx1_ASAP7_75t_L g846 ( .A(n_136), .Y(n_846) );
INVx1_ASAP7_75t_L g728 ( .A(n_137), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_139), .A2(n_152), .B1(n_267), .B2(n_270), .Y(n_313) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_140), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_141), .Y(n_954) );
CKINVDCx5p33_ASAP7_75t_R g1004 ( .A(n_142), .Y(n_1004) );
INVx1_ASAP7_75t_L g1074 ( .A(n_143), .Y(n_1074) );
XOR2x2_ASAP7_75t_L g640 ( .A(n_144), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g852 ( .A(n_145), .Y(n_852) );
INVx1_ASAP7_75t_L g524 ( .A(n_146), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_146), .A2(n_220), .B1(n_616), .B2(n_621), .Y(n_615) );
INVx1_ASAP7_75t_L g741 ( .A(n_147), .Y(n_741) );
INVx1_ASAP7_75t_L g823 ( .A(n_148), .Y(n_823) );
INVx1_ASAP7_75t_L g1130 ( .A(n_149), .Y(n_1130) );
INVx1_ASAP7_75t_L g1134 ( .A(n_150), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1325 ( .A1(n_151), .A2(n_231), .B1(n_621), .B2(n_1326), .Y(n_1325) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_153), .Y(n_891) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_154), .Y(n_573) );
INVx1_ASAP7_75t_L g1164 ( .A(n_155), .Y(n_1164) );
INVx1_ASAP7_75t_L g1061 ( .A(n_156), .Y(n_1061) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_158), .A2(n_218), .B1(n_259), .B2(n_264), .Y(n_289) );
INVx1_ASAP7_75t_L g521 ( .A(n_159), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g1275 ( .A1(n_160), .A2(n_227), .B1(n_1171), .B2(n_1276), .Y(n_1275) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_161), .A2(n_175), .B1(n_535), .B2(n_811), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_161), .A2(n_175), .B1(n_789), .B2(n_1111), .Y(n_1110) );
INVx1_ASAP7_75t_L g1002 ( .A(n_162), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_162), .B(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1203 ( .A(n_163), .Y(n_1203) );
INVx1_ASAP7_75t_L g693 ( .A(n_164), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_165), .A2(n_172), .B1(n_1227), .B2(n_1230), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_166), .B(n_513), .Y(n_1073) );
INVxp67_ASAP7_75t_SL g1082 ( .A(n_166), .Y(n_1082) );
OAI211xp5_ASAP7_75t_SL g821 ( .A1(n_167), .A2(n_801), .B(n_802), .C(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g834 ( .A(n_167), .Y(n_834) );
INVx1_ASAP7_75t_L g1167 ( .A(n_168), .Y(n_1167) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_169), .Y(n_904) );
INVx1_ASAP7_75t_L g1257 ( .A(n_170), .Y(n_1257) );
OAI211xp5_ASAP7_75t_L g919 ( .A1(n_171), .A2(n_649), .B(n_920), .C(n_921), .Y(n_919) );
INVx1_ASAP7_75t_L g941 ( .A(n_171), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g1238 ( .A1(n_172), .A2(n_236), .B1(n_1035), .B2(n_1239), .Y(n_1238) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_173), .A2(n_215), .B1(n_259), .B2(n_264), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_174), .A2(n_239), .B1(n_810), .B2(n_811), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_174), .A2(n_239), .B1(n_836), .B2(n_837), .Y(n_835) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_176), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_177), .A2(n_183), .B1(n_1206), .B2(n_1368), .Y(n_1370) );
INVx1_ASAP7_75t_L g1262 ( .A(n_178), .Y(n_1262) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_179), .Y(n_888) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_180), .Y(n_1314) );
AOI22xp33_ASAP7_75t_SL g1372 ( .A1(n_180), .A2(n_231), .B1(n_893), .B2(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g651 ( .A(n_181), .Y(n_651) );
AO22x1_ASAP7_75t_L g302 ( .A1(n_184), .A2(n_205), .B1(n_259), .B2(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g1131 ( .A(n_186), .Y(n_1131) );
INVx1_ASAP7_75t_L g1056 ( .A(n_187), .Y(n_1056) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_189), .Y(n_354) );
OA22x2_ASAP7_75t_L g1299 ( .A1(n_189), .A2(n_354), .B1(n_1300), .B2(n_1381), .Y(n_1299) );
INVx1_ASAP7_75t_L g784 ( .A(n_191), .Y(n_784) );
OAI211xp5_ASAP7_75t_L g800 ( .A1(n_191), .A2(n_801), .B(n_802), .C(n_803), .Y(n_800) );
INVx1_ASAP7_75t_L g684 ( .A(n_193), .Y(n_684) );
INVxp67_ASAP7_75t_SL g1084 ( .A(n_194), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_195), .A2(n_245), .B1(n_624), .B2(n_626), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_197), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_198), .A2(n_228), .B1(n_267), .B2(n_270), .Y(n_275) );
XOR2xp5_ASAP7_75t_L g944 ( .A(n_198), .B(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g999 ( .A(n_199), .Y(n_999) );
BUFx3_ASAP7_75t_L g475 ( .A(n_201), .Y(n_475) );
INVx1_ASAP7_75t_L g576 ( .A(n_201), .Y(n_576) );
INVx1_ASAP7_75t_L g781 ( .A(n_202), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_203), .Y(n_356) );
XOR2x2_ASAP7_75t_L g816 ( .A(n_206), .B(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_207), .Y(n_923) );
CKINVDCx5p33_ASAP7_75t_R g953 ( .A(n_209), .Y(n_953) );
INVx1_ASAP7_75t_L g1049 ( .A(n_210), .Y(n_1049) );
INVx1_ASAP7_75t_L g859 ( .A(n_212), .Y(n_859) );
INVxp67_ASAP7_75t_SL g1154 ( .A(n_213), .Y(n_1154) );
INVxp67_ASAP7_75t_SL g1155 ( .A(n_217), .Y(n_1155) );
INVx2_ASAP7_75t_L g516 ( .A(n_221), .Y(n_516) );
INVx1_ASAP7_75t_L g566 ( .A(n_221), .Y(n_566) );
INVx1_ASAP7_75t_L g768 ( .A(n_221), .Y(n_768) );
INVx1_ASAP7_75t_L g1100 ( .A(n_222), .Y(n_1100) );
INVx1_ASAP7_75t_L g1148 ( .A(n_223), .Y(n_1148) );
OAI211xp5_ASAP7_75t_L g1260 ( .A1(n_225), .A2(n_600), .B(n_1007), .C(n_1261), .Y(n_1260) );
AO22x1_ASAP7_75t_L g304 ( .A1(n_226), .A2(n_242), .B1(n_267), .B2(n_270), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_227), .A2(n_234), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_229), .Y(n_898) );
XNOR2xp5_ASAP7_75t_L g1144 ( .A(n_230), .B(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1346 ( .A(n_232), .Y(n_1346) );
INVx1_ASAP7_75t_L g1060 ( .A(n_233), .Y(n_1060) );
INVx1_ASAP7_75t_L g749 ( .A(n_235), .Y(n_749) );
INVx1_ASAP7_75t_L g1212 ( .A(n_237), .Y(n_1212) );
INVx1_ASAP7_75t_L g862 ( .A(n_240), .Y(n_862) );
AOI21xp33_ASAP7_75t_L g1013 ( .A1(n_241), .A2(n_624), .B(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1033 ( .A(n_241), .Y(n_1033) );
INVx1_ASAP7_75t_L g824 ( .A(n_243), .Y(n_824) );
OAI211xp5_ASAP7_75t_L g827 ( .A1(n_243), .A2(n_828), .B(n_831), .C(n_832), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g995 ( .A(n_246), .Y(n_995) );
INVx1_ASAP7_75t_L g569 ( .A(n_247), .Y(n_569) );
INVx1_ASAP7_75t_L g739 ( .A(n_248), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_259), .B1(n_452), .B2(n_476), .C(n_1249), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NOR2xp67_ASAP7_75t_SL g251 ( .A(n_252), .B(n_403), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_350), .B(n_358), .Y(n_252) );
NOR4xp25_ASAP7_75t_L g253 ( .A(n_254), .B(n_317), .C(n_329), .D(n_345), .Y(n_253) );
OAI211xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_272), .B(n_290), .C(n_305), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_256), .Y(n_255) );
OAI322xp33_ASAP7_75t_L g329 ( .A1(n_256), .A2(n_274), .A3(n_330), .B1(n_331), .B2(n_336), .C1(n_341), .C2(n_343), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_256), .A2(n_283), .B1(n_371), .B2(n_372), .Y(n_370) );
INVx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g299 ( .A(n_257), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g309 ( .A(n_257), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g335 ( .A(n_257), .Y(n_335) );
AND2x2_ASAP7_75t_L g366 ( .A(n_257), .B(n_319), .Y(n_366) );
OR2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_311), .Y(n_373) );
AND2x2_ASAP7_75t_L g380 ( .A(n_257), .B(n_301), .Y(n_380) );
AND2x2_ASAP7_75t_L g398 ( .A(n_257), .B(n_300), .Y(n_398) );
AND2x2_ASAP7_75t_L g422 ( .A(n_257), .B(n_311), .Y(n_422) );
OR2x2_ASAP7_75t_L g442 ( .A(n_257), .B(n_301), .Y(n_442) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_266), .Y(n_257) );
INVx2_ASAP7_75t_L g355 ( .A(n_259), .Y(n_355) );
AND2x6_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x2_ASAP7_75t_L g264 ( .A(n_260), .B(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g267 ( .A(n_260), .B(n_268), .Y(n_267) );
AND2x6_ASAP7_75t_L g270 ( .A(n_260), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_260), .B(n_265), .Y(n_277) );
AND2x2_ASAP7_75t_L g303 ( .A(n_260), .B(n_265), .Y(n_303) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_261), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g1386 ( .A1(n_262), .A2(n_1387), .B(n_1388), .Y(n_1386) );
AND2x2_ASAP7_75t_L g268 ( .A(n_263), .B(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g357 ( .A(n_264), .Y(n_357) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_278), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_273), .B(n_287), .Y(n_293) );
AND2x2_ASAP7_75t_L g325 ( .A(n_273), .B(n_326), .Y(n_325) );
AND3x1_ASAP7_75t_L g378 ( .A(n_273), .B(n_287), .C(n_297), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_273), .B(n_297), .Y(n_386) );
AND2x2_ASAP7_75t_L g396 ( .A(n_273), .B(n_279), .Y(n_396) );
AND2x2_ASAP7_75t_L g416 ( .A(n_273), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
BUFx2_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
AND2x2_ASAP7_75t_L g342 ( .A(n_274), .B(n_326), .Y(n_342) );
OR2x2_ASAP7_75t_L g348 ( .A(n_274), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g382 ( .A(n_274), .B(n_283), .Y(n_382) );
AND2x2_ASAP7_75t_L g435 ( .A(n_274), .B(n_417), .Y(n_435) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .Y(n_278) );
INVx1_ASAP7_75t_L g308 ( .A(n_279), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_279), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_279), .B(n_326), .Y(n_374) );
AND2x2_ASAP7_75t_L g412 ( .A(n_279), .B(n_334), .Y(n_412) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g291 ( .A(n_280), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g315 ( .A(n_280), .B(n_311), .Y(n_315) );
AND2x2_ASAP7_75t_L g319 ( .A(n_280), .B(n_311), .Y(n_319) );
INVx1_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
AND2x2_ASAP7_75t_L g389 ( .A(n_280), .B(n_301), .Y(n_389) );
AND2x2_ASAP7_75t_L g402 ( .A(n_280), .B(n_295), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_280), .B(n_310), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_280), .B(n_320), .Y(n_440) );
OR2x2_ASAP7_75t_L g443 ( .A(n_280), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g349 ( .A(n_283), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_283), .B(n_396), .Y(n_438) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
INVx2_ASAP7_75t_L g297 ( .A(n_284), .Y(n_297) );
AND2x2_ASAP7_75t_L g326 ( .A(n_284), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_284), .B(n_295), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_284), .B(n_352), .C(n_407), .Y(n_445) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g296 ( .A(n_287), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g327 ( .A(n_287), .Y(n_327) );
OAI211xp5_ASAP7_75t_L g369 ( .A1(n_287), .A2(n_315), .B(n_370), .C(n_374), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_287), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_294), .B(n_298), .Y(n_290) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_293), .B(n_308), .Y(n_371) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_293), .A2(n_348), .B1(n_379), .B2(n_425), .C(n_426), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_293), .A2(n_315), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g364 ( .A(n_294), .B(n_324), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_294), .B(n_325), .Y(n_410) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g316 ( .A(n_295), .B(n_297), .Y(n_316) );
OR2x2_ASAP7_75t_L g320 ( .A(n_295), .B(n_297), .Y(n_320) );
OR2x2_ASAP7_75t_L g330 ( .A(n_296), .B(n_326), .Y(n_330) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_296), .B(n_337), .C(n_340), .Y(n_336) );
AND2x2_ASAP7_75t_L g395 ( .A(n_296), .B(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_297), .A2(n_325), .B1(n_366), .B2(n_367), .C(n_369), .Y(n_365) );
AND2x2_ASAP7_75t_L g417 ( .A(n_297), .B(n_327), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_298), .A2(n_427), .B(n_429), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_298), .B(n_364), .Y(n_431) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_300), .B(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_SL g332 ( .A(n_300), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g344 ( .A(n_300), .B(n_310), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_300), .B(n_352), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_300), .B(n_372), .Y(n_383) );
AND2x2_ASAP7_75t_L g436 ( .A(n_300), .B(n_334), .Y(n_436) );
CKINVDCx6p67_ASAP7_75t_R g300 ( .A(n_301), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_301), .Y(n_328) );
OR2x2_ASAP7_75t_L g346 ( .A(n_301), .B(n_347), .Y(n_346) );
OR2x6_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
OR2x2_ASAP7_75t_L g340 ( .A(n_302), .B(n_304), .Y(n_340) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_314), .B(n_316), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
CKINVDCx6p67_ASAP7_75t_R g347 ( .A(n_309), .Y(n_347) );
INVx2_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g334 ( .A(n_311), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
CKINVDCx14_ASAP7_75t_R g392 ( .A(n_316), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_316), .B(n_412), .Y(n_411) );
O2A1O1Ixp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_320), .B(n_321), .C(n_328), .Y(n_317) );
AOI21xp33_ASAP7_75t_L g449 ( .A1(n_318), .A2(n_450), .B(n_451), .Y(n_449) );
CKINVDCx14_ASAP7_75t_R g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
AND2x2_ASAP7_75t_L g377 ( .A(n_323), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g407 ( .A(n_323), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_323), .B(n_372), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_323), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_325), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g450 ( .A(n_325), .Y(n_450) );
AND2x2_ASAP7_75t_L g401 ( .A(n_326), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g430 ( .A(n_326), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g420 ( .A1(n_328), .A2(n_341), .B(n_421), .C(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_333), .A2(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_334), .B(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_337), .B(n_342), .Y(n_448) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
AND2x2_ASAP7_75t_L g419 ( .A(n_339), .B(n_342), .Y(n_419) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI21xp5_ASAP7_75t_SL g384 ( .A1(n_342), .A2(n_385), .B(n_387), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_343), .A2(n_347), .B1(n_438), .B2(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_347), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_441) );
OAI31xp33_ASAP7_75t_SL g418 ( .A1(n_350), .A2(n_419), .A3(n_420), .B(n_424), .Y(n_418) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g393 ( .A(n_352), .Y(n_393) );
OAI22xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_355), .B1(n_356), .B2(n_357), .Y(n_353) );
OAI222xp33_ASAP7_75t_L g1249 ( .A1(n_354), .A2(n_1250), .B1(n_1293), .B2(n_1297), .C1(n_1382), .C2(n_1385), .Y(n_1249) );
AOI211xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B(n_375), .C(n_390), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .B(n_365), .Y(n_361) );
INVx2_ASAP7_75t_L g368 ( .A(n_362), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_362), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_362), .B(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_366), .Y(n_391) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
OAI321xp33_ASAP7_75t_L g390 ( .A1(n_373), .A2(n_391), .A3(n_392), .B1(n_393), .B2(n_394), .C(n_397), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_381), .B2(n_383), .C(n_384), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_380), .B(n_407), .Y(n_425) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_380), .A2(n_447), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
AOI211xp5_ASAP7_75t_L g404 ( .A1(n_398), .A2(n_405), .B(n_408), .C(n_413), .Y(n_404) );
INVx1_ASAP7_75t_L g414 ( .A(n_398), .Y(n_414) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND5xp2_ASAP7_75t_L g403 ( .A(n_404), .B(n_418), .C(n_431), .D(n_432), .E(n_446), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g423 ( .A(n_416), .Y(n_423) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NOR3xp33_ASAP7_75t_SL g432 ( .A(n_433), .B(n_437), .C(n_441), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g451 ( .A(n_435), .Y(n_451) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_461), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_456), .B(n_464), .Y(n_1384) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g1296 ( .A(n_458), .B(n_460), .Y(n_1296) );
INVx1_ASAP7_75t_L g1387 ( .A(n_458), .Y(n_1387) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g1389 ( .A(n_460), .B(n_1387), .Y(n_1389) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g603 ( .A(n_464), .B(n_604), .Y(n_603) );
AOI21xp5_ASAP7_75t_SL g986 ( .A1(n_464), .A2(n_987), .B(n_1000), .Y(n_986) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x4_ASAP7_75t_L g630 ( .A(n_465), .B(n_475), .Y(n_630) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_465), .B(n_474), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g1172 ( .A1(n_466), .A2(n_574), .B1(n_1173), .B2(n_1174), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1256 ( .A1(n_466), .A2(n_574), .B1(n_1257), .B2(n_1258), .Y(n_1256) );
AND2x4_ASAP7_75t_SL g1383 ( .A(n_466), .B(n_1384), .Y(n_1383) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_468), .B(n_473), .Y(n_467) );
OR2x2_ASAP7_75t_L g581 ( .A(n_468), .B(n_575), .Y(n_581) );
OR2x6_ASAP7_75t_L g789 ( .A(n_468), .B(n_575), .Y(n_789) );
INVx1_ASAP7_75t_L g916 ( .A(n_468), .Y(n_916) );
BUFx4f_ASAP7_75t_L g1003 ( .A(n_468), .Y(n_1003) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g572 ( .A(n_469), .Y(n_572) );
BUFx4f_ASAP7_75t_L g672 ( .A(n_469), .Y(n_672) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x2_ASAP7_75t_L g577 ( .A(n_471), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g586 ( .A(n_471), .Y(n_586) );
INVx1_ASAP7_75t_L g593 ( .A(n_471), .Y(n_593) );
AND2x2_ASAP7_75t_L g599 ( .A(n_471), .B(n_472), .Y(n_599) );
INVx2_ASAP7_75t_L g619 ( .A(n_471), .Y(n_619) );
NAND2x1_ASAP7_75t_L g648 ( .A(n_471), .B(n_472), .Y(n_648) );
INVx2_ASAP7_75t_L g578 ( .A(n_472), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_472), .B(n_586), .Y(n_585) );
BUFx2_ASAP7_75t_L g590 ( .A(n_472), .Y(n_590) );
INVx1_ASAP7_75t_L g620 ( .A(n_472), .Y(n_620) );
AND2x2_ASAP7_75t_L g622 ( .A(n_472), .B(n_586), .Y(n_622) );
OR2x2_ASAP7_75t_L g681 ( .A(n_472), .B(n_619), .Y(n_681) );
OR2x6_ASAP7_75t_L g571 ( .A(n_473), .B(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g994 ( .A1(n_473), .A2(n_995), .B1(n_996), .B2(n_997), .Y(n_994) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g583 ( .A(n_474), .Y(n_583) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x4_ASAP7_75t_L g591 ( .A(n_475), .B(n_592), .Y(n_591) );
BUFx2_ASAP7_75t_L g653 ( .A(n_475), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B1(n_1089), .B2(n_1090), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
XOR2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_879), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_718), .B2(n_878), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
XNOR2x1_ASAP7_75t_L g483 ( .A(n_484), .B(n_640), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_606), .Y(n_484) );
INVx1_ASAP7_75t_L g608 ( .A(n_486), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_500), .B(n_517), .Y(n_486) );
BUFx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g520 ( .A(n_489), .Y(n_520) );
INVx2_ASAP7_75t_L g541 ( .A(n_489), .Y(n_541) );
AND2x4_ASAP7_75t_L g543 ( .A(n_489), .B(n_530), .Y(n_543) );
BUFx2_ASAP7_75t_L g662 ( .A(n_489), .Y(n_662) );
BUFx2_ASAP7_75t_L g1037 ( .A(n_489), .Y(n_1037) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_489), .Y(n_1072) );
BUFx2_ASAP7_75t_L g1206 ( .A(n_489), .Y(n_1206) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g509 ( .A(n_490), .Y(n_509) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g552 ( .A(n_491), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_491), .B(n_492), .Y(n_558) );
INVx2_ASAP7_75t_L g496 ( .A(n_492), .Y(n_496) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_492), .Y(n_508) );
OR2x2_ASAP7_75t_L g534 ( .A(n_492), .B(n_498), .Y(n_534) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g1189 ( .A(n_494), .Y(n_1189) );
INVx8_ASAP7_75t_L g1241 ( .A(n_494), .Y(n_1241) );
INVx8_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx3_ASAP7_75t_L g523 ( .A(n_495), .Y(n_523) );
BUFx3_ASAP7_75t_L g1248 ( .A(n_495), .Y(n_1248) );
NAND2x1p5_ASAP7_75t_L g1353 ( .A(n_495), .B(n_1354), .Y(n_1353) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
AND2x4_ASAP7_75t_L g503 ( .A(n_496), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g504 ( .A(n_499), .Y(n_504) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g555 ( .A(n_502), .B(n_536), .Y(n_555) );
INVx2_ASAP7_75t_L g710 ( .A(n_502), .Y(n_710) );
AND2x4_ASAP7_75t_L g799 ( .A(n_502), .B(n_536), .Y(n_799) );
BUFx6f_ASAP7_75t_L g1035 ( .A(n_502), .Y(n_1035) );
INVx2_ASAP7_75t_L g1186 ( .A(n_502), .Y(n_1186) );
INVx1_ASAP7_75t_L g1290 ( .A(n_502), .Y(n_1290) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_503), .Y(n_705) );
BUFx8_ASAP7_75t_L g893 ( .A(n_503), .Y(n_893) );
INVx2_ASAP7_75t_L g1042 ( .A(n_503), .Y(n_1042) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_R g1287 ( .A(n_506), .Y(n_1287) );
INVx5_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_507), .Y(n_1039) );
BUFx12f_ASAP7_75t_L g1239 ( .A(n_507), .Y(n_1239) );
BUFx3_ASAP7_75t_L g1373 ( .A(n_507), .Y(n_1373) );
AND2x4_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
BUFx2_ASAP7_75t_L g548 ( .A(n_508), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_508), .B(n_552), .Y(n_702) );
INVx2_ASAP7_75t_L g940 ( .A(n_508), .Y(n_940) );
INVx1_ASAP7_75t_L g938 ( .A(n_509), .Y(n_938) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND3xp33_ASAP7_75t_L g1237 ( .A(n_511), .B(n_1238), .C(n_1240), .Y(n_1237) );
AOI33xp33_ASAP7_75t_L g1281 ( .A1(n_511), .A2(n_1282), .A3(n_1285), .B1(n_1288), .B2(n_1291), .B3(n_1292), .Y(n_1281) );
AOI33xp33_ASAP7_75t_L g1366 ( .A1(n_511), .A2(n_1367), .A3(n_1369), .B1(n_1370), .B2(n_1371), .B3(n_1372), .Y(n_1366) );
AND3x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .C(n_515), .Y(n_511) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_512), .Y(n_561) );
NAND2xp33_ASAP7_75t_SL g697 ( .A(n_512), .B(n_514), .Y(n_697) );
INVx1_ASAP7_75t_L g1355 ( .A(n_512), .Y(n_1355) );
INVx3_ASAP7_75t_L g547 ( .A(n_513), .Y(n_547) );
AND2x2_ASAP7_75t_L g937 ( .A(n_513), .B(n_938), .Y(n_937) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g530 ( .A(n_514), .Y(n_530) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g527 ( .A(n_516), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_521), .B1(n_522), .B2(n_524), .C(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
BUFx3_ASAP7_75t_L g1368 ( .A(n_523), .Y(n_1368) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI33xp33_ASAP7_75t_L g1047 ( .A1(n_526), .A2(n_844), .A3(n_1048), .B1(n_1051), .B2(n_1054), .B3(n_1059), .Y(n_1047) );
OAI33xp33_ASAP7_75t_L g1115 ( .A1(n_526), .A2(n_844), .A3(n_1116), .B1(n_1123), .B2(n_1128), .B3(n_1132), .Y(n_1115) );
INVx1_ASAP7_75t_L g1292 ( .A(n_526), .Y(n_1292) );
INVx1_ASAP7_75t_SL g1371 ( .A(n_526), .Y(n_1371) );
OR2x6_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x4_ASAP7_75t_L g613 ( .A(n_527), .B(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g712 ( .A(n_527), .B(n_528), .Y(n_712) );
INVx1_ASAP7_75t_L g1019 ( .A(n_527), .Y(n_1019) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND3x1_ASAP7_75t_L g766 ( .A(n_529), .B(n_530), .C(n_767), .Y(n_766) );
OR2x4_ASAP7_75t_L g533 ( .A(n_530), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g536 ( .A(n_530), .Y(n_536) );
OR2x6_ASAP7_75t_L g556 ( .A(n_530), .B(n_557), .Y(n_556) );
AND2x4_ASAP7_75t_L g1354 ( .A(n_530), .B(n_1355), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_531), .B(n_567), .Y(n_607) );
OAI31xp33_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_537), .A3(n_553), .B(n_559), .Y(n_531) );
INVx2_ASAP7_75t_SL g797 ( .A(n_533), .Y(n_797) );
INVx1_ASAP7_75t_L g1029 ( .A(n_533), .Y(n_1029) );
INVx2_ASAP7_75t_SL g1202 ( .A(n_533), .Y(n_1202) );
OR2x4_ASAP7_75t_L g535 ( .A(n_534), .B(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g700 ( .A(n_534), .Y(n_700) );
BUFx4f_ASAP7_75t_L g714 ( .A(n_534), .Y(n_714) );
BUFx3_ASAP7_75t_L g755 ( .A(n_534), .Y(n_755) );
BUFx3_ASAP7_75t_L g847 ( .A(n_534), .Y(n_847) );
BUFx3_ASAP7_75t_L g810 ( .A(n_535), .Y(n_810) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_535), .Y(n_1182) );
INVx2_ASAP7_75t_SL g1211 ( .A(n_535), .Y(n_1211) );
NAND3xp33_ASAP7_75t_SL g537 ( .A(n_538), .B(n_542), .C(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_539), .A2(n_545), .B1(n_589), .B2(n_591), .Y(n_588) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g1177 ( .A(n_541), .Y(n_1177) );
INVx1_ASAP7_75t_L g1284 ( .A(n_541), .Y(n_1284) );
NAND3xp33_ASAP7_75t_SL g660 ( .A(n_542), .B(n_661), .C(n_663), .Y(n_660) );
CKINVDCx8_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
CKINVDCx8_ASAP7_75t_R g802 ( .A(n_543), .Y(n_802) );
NOR3xp33_ASAP7_75t_L g1022 ( .A(n_543), .B(n_1023), .C(n_1027), .Y(n_1022) );
AOI211xp5_ASAP7_75t_L g1176 ( .A1(n_543), .A2(n_1168), .B(n_1177), .C(n_1178), .Y(n_1176) );
AOI211xp5_ASAP7_75t_L g1204 ( .A1(n_543), .A2(n_1205), .B(n_1206), .C(n_1207), .Y(n_1204) );
NOR3xp33_ASAP7_75t_L g1266 ( .A(n_543), .B(n_1267), .C(n_1268), .Y(n_1266) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_549), .B2(n_550), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_546), .A2(n_550), .B1(n_651), .B2(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_546), .A2(n_937), .B1(n_973), .B2(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1025 ( .A(n_546), .Y(n_1025) );
AOI222xp33_ASAP7_75t_L g1071 ( .A1(n_546), .A2(n_550), .B1(n_1072), .B2(n_1073), .C1(n_1074), .C2(n_1075), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1270 ( .A(n_546), .B(n_1262), .Y(n_1270) );
AND2x4_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
AND2x2_ASAP7_75t_L g550 ( .A(n_547), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g805 ( .A(n_547), .B(n_548), .Y(n_805) );
AND2x4_ASAP7_75t_L g807 ( .A(n_547), .B(n_551), .Y(n_807) );
AND2x4_ASAP7_75t_L g935 ( .A(n_547), .B(n_548), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_549), .B(n_595), .Y(n_594) );
AOI32xp33_ASAP7_75t_L g936 ( .A1(n_550), .A2(n_923), .A3(n_937), .B1(n_939), .B2(n_941), .Y(n_936) );
INVxp67_ASAP7_75t_L g980 ( .A(n_550), .Y(n_980) );
INVxp67_ASAP7_75t_L g1026 ( .A(n_550), .Y(n_1026) );
INVx1_ASAP7_75t_L g1208 ( .A(n_550), .Y(n_1208) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g1028 ( .A1(n_555), .A2(n_995), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
INVx1_ASAP7_75t_L g812 ( .A(n_556), .Y(n_812) );
INVx2_ASAP7_75t_L g1078 ( .A(n_556), .Y(n_1078) );
INVx1_ASAP7_75t_L g1213 ( .A(n_556), .Y(n_1213) );
BUFx3_ASAP7_75t_L g763 ( .A(n_557), .Y(n_763) );
INVx1_ASAP7_75t_L g895 ( .A(n_557), .Y(n_895) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g708 ( .A(n_558), .Y(n_708) );
OAI31xp33_ASAP7_75t_SL g658 ( .A1(n_559), .A2(n_659), .A3(n_660), .B(n_665), .Y(n_658) );
OAI31xp33_ASAP7_75t_L g1096 ( .A1(n_559), .A2(n_1097), .A3(n_1098), .B(n_1102), .Y(n_1096) );
INVx1_ASAP7_75t_L g1183 ( .A(n_559), .Y(n_1183) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x2_ASAP7_75t_SL g814 ( .A(n_560), .B(n_562), .Y(n_814) );
AND2x2_ASAP7_75t_L g943 ( .A(n_560), .B(n_562), .Y(n_943) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_564), .B(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g696 ( .A(n_564), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g745 ( .A(n_564), .Y(n_745) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_564), .B(n_1342), .Y(n_1341) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g605 ( .A(n_565), .Y(n_605) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AO21x1_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_579), .B(n_602), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_573), .B2(n_574), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g1216 ( .A(n_571), .Y(n_1216) );
BUFx3_ASAP7_75t_L g747 ( .A(n_572), .Y(n_747) );
BUFx3_ASAP7_75t_L g963 ( .A(n_572), .Y(n_963) );
BUFx6f_ASAP7_75t_L g1068 ( .A(n_572), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1138 ( .A(n_572), .Y(n_1138) );
INVx4_ASAP7_75t_L g657 ( .A(n_574), .Y(n_657) );
CKINVDCx16_ASAP7_75t_R g841 ( .A(n_574), .Y(n_841) );
INVx3_ASAP7_75t_SL g988 ( .A(n_574), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_574), .A2(n_1201), .B1(n_1203), .B2(n_1216), .Y(n_1215) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_577), .Y(n_625) );
BUFx3_ASAP7_75t_L g1229 ( .A(n_577), .Y(n_1229) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_587), .Y(n_579) );
INVx1_ASAP7_75t_L g1087 ( .A(n_582), .Y(n_1087) );
OR2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x2_ASAP7_75t_L g589 ( .A(n_583), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g601 ( .A(n_583), .B(n_597), .Y(n_601) );
AND2x2_ASAP7_75t_L g786 ( .A(n_583), .B(n_627), .Y(n_786) );
INVx8_ASAP7_75t_L g675 ( .A(n_584), .Y(n_675) );
OR2x2_ASAP7_75t_L g792 ( .A(n_584), .B(n_653), .Y(n_792) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_584), .Y(n_1139) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_594), .C(n_600), .Y(n_587) );
INVx1_ASAP7_75t_L g993 ( .A(n_589), .Y(n_993) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_589), .A2(n_924), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
AOI22xp5_ASAP7_75t_L g1261 ( .A1(n_589), .A2(n_924), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
AND2x4_ASAP7_75t_L g652 ( .A(n_590), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g833 ( .A(n_590), .B(n_653), .Y(n_833) );
BUFx2_ASAP7_75t_L g1310 ( .A(n_590), .Y(n_1310) );
BUFx3_ASAP7_75t_L g655 ( .A(n_591), .Y(n_655) );
INVx2_ASAP7_75t_L g783 ( .A(n_591), .Y(n_783) );
INVx2_ASAP7_75t_L g925 ( .A(n_591), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_592), .B(n_1311), .Y(n_1351) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g1219 ( .A(n_598), .Y(n_1219) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_599), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g1165 ( .A(n_600), .B(n_1166), .C(n_1169), .Y(n_1165) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g649 ( .A(n_601), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g1217 ( .A1(n_601), .A2(n_1218), .B(n_1220), .C(n_1221), .Y(n_1217) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_602), .A2(n_1162), .B(n_1172), .Y(n_1161) );
AO21x1_ASAP7_75t_L g1255 ( .A1(n_602), .A2(n_1256), .B(n_1259), .Y(n_1255) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI31xp33_ASAP7_75t_L g642 ( .A1(n_603), .A2(n_643), .A3(n_644), .B(n_656), .Y(n_642) );
BUFx3_ASAP7_75t_L g793 ( .A(n_603), .Y(n_793) );
BUFx2_ASAP7_75t_L g930 ( .A(n_603), .Y(n_930) );
OAI31xp33_ASAP7_75t_L g969 ( .A1(n_603), .A2(n_970), .A3(n_971), .B(n_975), .Y(n_969) );
OAI21xp5_ASAP7_75t_L g1079 ( .A1(n_603), .A2(n_1080), .B(n_1088), .Y(n_1079) );
BUFx2_ASAP7_75t_SL g1113 ( .A(n_603), .Y(n_1113) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g1350 ( .A(n_605), .B(n_1351), .Y(n_1350) );
INVxp67_ASAP7_75t_L g1356 ( .A(n_605), .Y(n_1356) );
OAI31xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .A3(n_609), .B(n_637), .Y(n_606) );
INVx1_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
AOI33xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_615), .A3(n_623), .B1(n_628), .B2(n_629), .B3(n_631), .Y(n_610) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_611), .Y(n_1233) );
AOI33xp33_ASAP7_75t_L g1272 ( .A1(n_611), .A2(n_629), .A3(n_1273), .B1(n_1275), .B2(n_1278), .B3(n_1279), .Y(n_1272) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
OAI33xp33_ASAP7_75t_L g1135 ( .A1(n_612), .A2(n_689), .A3(n_1136), .B1(n_1140), .B2(n_1142), .B3(n_1143), .Y(n_1135) );
INVx4_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g668 ( .A(n_613), .Y(n_668) );
INVx2_ASAP7_75t_L g724 ( .A(n_613), .Y(n_724) );
INVx2_ASAP7_75t_L g906 ( .A(n_613), .Y(n_906) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g1017 ( .A(n_617), .Y(n_1017) );
INVx1_ASAP7_75t_L g1232 ( .A(n_617), .Y(n_1232) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_618), .Y(n_634) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_618), .B(n_1307), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_618), .B(n_1311), .Y(n_1345) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
BUFx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g636 ( .A(n_622), .Y(n_636) );
BUFx6f_ASAP7_75t_L g1159 ( .A(n_622), .Y(n_1159) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g1277 ( .A(n_625), .Y(n_1277) );
AND2x4_ASAP7_75t_L g1335 ( .A(n_625), .B(n_1307), .Y(n_1335) );
BUFx3_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx3_ASAP7_75t_L g991 ( .A(n_627), .Y(n_991) );
BUFx6f_ASAP7_75t_L g1171 ( .A(n_627), .Y(n_1171) );
BUFx3_ASAP7_75t_L g1230 ( .A(n_627), .Y(n_1230) );
AND2x4_ASAP7_75t_SL g1306 ( .A(n_627), .B(n_1307), .Y(n_1306) );
AND2x6_ASAP7_75t_L g1327 ( .A(n_627), .B(n_1311), .Y(n_1327) );
INVx2_ASAP7_75t_L g689 ( .A(n_629), .Y(n_689) );
INVx2_ASAP7_75t_L g917 ( .A(n_629), .Y(n_917) );
AND2x4_ASAP7_75t_L g743 ( .A(n_630), .B(n_744), .Y(n_743) );
OAI221xp5_ASAP7_75t_L g1006 ( .A1(n_630), .A2(n_869), .B1(n_1007), .B2(n_1008), .C(n_1009), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_630), .B(n_744), .Y(n_1160) );
INVx4_ASAP7_75t_L g1324 ( .A(n_630), .Y(n_1324) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g1280 ( .A(n_633), .Y(n_1280) );
INVx2_ASAP7_75t_L g1326 ( .A(n_633), .Y(n_1326) );
INVx3_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_634), .B(n_653), .Y(n_1085) );
BUFx6f_ASAP7_75t_L g1274 ( .A(n_634), .Y(n_1274) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g1151 ( .A(n_636), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
NAND3xp33_ASAP7_75t_SL g641 ( .A(n_642), .B(n_658), .C(n_666), .Y(n_641) );
INVx5_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_647), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
BUFx2_ASAP7_75t_SL g740 ( .A(n_647), .Y(n_740) );
BUFx3_ASAP7_75t_L g830 ( .A(n_647), .Y(n_830) );
BUFx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_648), .Y(n_683) );
NAND3xp33_ASAP7_75t_SL g1080 ( .A(n_649), .B(n_1081), .C(n_1083), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_654), .B2(n_655), .Y(n_650) );
BUFx3_ASAP7_75t_L g780 ( .A(n_652), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_652), .A2(n_655), .B1(n_973), .B2(n_974), .Y(n_972) );
INVx1_ASAP7_75t_L g1222 ( .A(n_652), .Y(n_1222) );
O2A1O1Ixp33_ASAP7_75t_L g989 ( .A1(n_653), .A2(n_990), .B(n_991), .C(n_992), .Y(n_989) );
INVx1_ASAP7_75t_L g996 ( .A(n_653), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_654), .B(n_662), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g1081 ( .A1(n_655), .A2(n_833), .B1(n_991), .B2(n_1074), .C1(n_1075), .C2(n_1082), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_694), .Y(n_666) );
OAI33xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .A3(n_677), .B1(n_685), .B2(n_689), .B3(n_690), .Y(n_667) );
OAI33xp33_ASAP7_75t_L g961 ( .A1(n_668), .A2(n_917), .A3(n_962), .B1(n_964), .B2(n_965), .B3(n_968), .Y(n_961) );
BUFx6f_ASAP7_75t_L g1152 ( .A(n_668), .Y(n_1152) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B1(n_673), .B2(n_676), .Y(n_669) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_670), .A2(n_686), .B1(n_699), .B2(n_701), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_671), .A2(n_691), .B1(n_692), .B2(n_693), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_671), .A2(n_887), .B1(n_903), .B2(n_908), .Y(n_907) );
INVx4_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx3_ASAP7_75t_L g727 ( .A(n_672), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g962 ( .A1(n_673), .A2(n_949), .B1(n_959), .B2(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_673), .A2(n_1053), .B1(n_1058), .B2(n_1068), .Y(n_1067) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g692 ( .A(n_675), .Y(n_692) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_675), .Y(n_730) );
INVx4_ASAP7_75t_L g908 ( .A(n_675), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g713 ( .A1(n_676), .A2(n_688), .B1(n_714), .B2(n_715), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_682), .B2(n_684), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_678), .A2(n_691), .B1(n_704), .B2(n_706), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_679), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_685) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g733 ( .A(n_680), .Y(n_733) );
BUFx2_ASAP7_75t_L g870 ( .A(n_680), .Y(n_870) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g738 ( .A(n_681), .Y(n_738) );
INVx1_ASAP7_75t_L g911 ( .A(n_681), .Y(n_911) );
BUFx3_ASAP7_75t_L g966 ( .A(n_681), .Y(n_966) );
BUFx2_ASAP7_75t_L g1141 ( .A(n_681), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_682), .A2(n_1050), .B1(n_1061), .B2(n_1066), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1153 ( .A1(n_682), .A2(n_736), .B1(n_1154), .B2(n_1155), .C(n_1156), .Y(n_1153) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
BUFx4f_ASAP7_75t_L g687 ( .A(n_683), .Y(n_687) );
BUFx4f_ASAP7_75t_L g778 ( .A(n_683), .Y(n_778) );
INVx4_ASAP7_75t_L g872 ( .A(n_683), .Y(n_872) );
BUFx4f_ASAP7_75t_L g920 ( .A(n_683), .Y(n_920) );
BUFx4f_ASAP7_75t_L g1012 ( .A(n_683), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_684), .A2(n_693), .B1(n_710), .B2(n_711), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g964 ( .A1(n_687), .A2(n_910), .B1(n_953), .B2(n_956), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g1147 ( .A1(n_687), .A2(n_1066), .B1(n_1148), .B2(n_1149), .C(n_1150), .Y(n_1147) );
OAI211xp5_ASAP7_75t_L g1313 ( .A1(n_687), .A2(n_1314), .B(n_1315), .C(n_1317), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_692), .A2(n_1127), .B1(n_1131), .B2(n_1137), .Y(n_1143) );
OAI33xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_698), .A3(n_703), .B1(n_709), .B2(n_712), .B3(n_713), .Y(n_694) );
OAI33xp33_ASAP7_75t_L g885 ( .A1(n_695), .A2(n_712), .A3(n_886), .B1(n_890), .B2(n_897), .B3(n_902), .Y(n_885) );
OAI33xp33_ASAP7_75t_L g947 ( .A1(n_695), .A2(n_712), .A3(n_948), .B1(n_952), .B2(n_955), .B3(n_958), .Y(n_947) );
BUFx4f_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx4f_ASAP7_75t_L g751 ( .A(n_696), .Y(n_751) );
BUFx2_ASAP7_75t_L g844 ( .A(n_696), .Y(n_844) );
OR2x6_ASAP7_75t_L g1375 ( .A(n_699), .B(n_1376), .Y(n_1375) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx3_ASAP7_75t_L g1119 ( .A(n_700), .Y(n_1119) );
INVx2_ASAP7_75t_L g757 ( .A(n_701), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_701), .A2(n_714), .B1(n_903), .B2(n_904), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g958 ( .A1(n_701), .A2(n_714), .B1(n_959), .B2(n_960), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g1132 ( .A1(n_701), .A2(n_1119), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
BUFx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_702), .Y(n_717) );
BUFx2_ASAP7_75t_L g772 ( .A(n_702), .Y(n_772) );
INVx2_ASAP7_75t_L g857 ( .A(n_704), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g897 ( .A1(n_704), .A2(n_898), .B1(n_899), .B2(n_901), .Y(n_897) );
INVx3_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx5_ASAP7_75t_L g759 ( .A(n_705), .Y(n_759) );
INVx2_ASAP7_75t_SL g762 ( .A(n_705), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g952 ( .A1(n_706), .A2(n_710), .B1(n_953), .B2(n_954), .Y(n_952) );
INVx3_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g711 ( .A(n_707), .Y(n_711) );
CKINVDCx8_ASAP7_75t_R g760 ( .A(n_707), .Y(n_760) );
INVx3_ASAP7_75t_L g1057 ( .A(n_707), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g900 ( .A(n_708), .Y(n_900) );
OAI221xp5_ASAP7_75t_L g1190 ( .A1(n_710), .A2(n_711), .B1(n_1149), .B2(n_1191), .C(n_1192), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_711), .A2(n_762), .B1(n_956), .B2(n_957), .Y(n_955) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_714), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_886) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_714), .A2(n_949), .B1(n_950), .B2(n_951), .Y(n_948) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_714), .A2(n_1024), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_714), .A2(n_889), .B1(n_1060), .B2(n_1061), .Y(n_1059) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g801 ( .A(n_716), .Y(n_801) );
INVx2_ASAP7_75t_L g1024 ( .A(n_716), .Y(n_1024) );
INVx4_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx3_ASAP7_75t_L g850 ( .A(n_717), .Y(n_850) );
BUFx6f_ASAP7_75t_L g889 ( .A(n_717), .Y(n_889) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_717), .B(n_1341), .Y(n_1349) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_815), .B(n_877), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g878 ( .A1(n_719), .A2(n_815), .B(n_877), .Y(n_878) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g877 ( .A(n_720), .B(n_816), .Y(n_877) );
NAND3xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_773), .C(n_794), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_750), .Y(n_722) );
OAI33xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .A3(n_731), .B1(n_735), .B2(n_742), .B3(n_746), .Y(n_723) );
OAI33xp33_ASAP7_75t_L g864 ( .A1(n_724), .A2(n_865), .A3(n_868), .B1(n_873), .B2(n_875), .B3(n_876), .Y(n_864) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_726), .A2(n_739), .B1(n_753), .B2(n_756), .Y(n_752) );
INVx2_ASAP7_75t_SL g867 ( .A(n_727), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g769 ( .A1(n_728), .A2(n_741), .B1(n_753), .B2(n_770), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_729), .A2(n_747), .B1(n_748), .B2(n_749), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_729), .A2(n_846), .B1(n_862), .B2(n_866), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_729), .A2(n_854), .B1(n_859), .B2(n_866), .Y(n_876) );
INVx6_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx5_ASAP7_75t_L g1005 ( .A(n_730), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_732), .A2(n_748), .B1(n_759), .B2(n_760), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_734), .A2(n_749), .B1(n_762), .B2(n_763), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_739), .B1(n_740), .B2(n_741), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx4_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_743), .Y(n_875) );
NAND3xp33_ASAP7_75t_L g1234 ( .A(n_743), .B(n_1235), .C(n_1236), .Y(n_1234) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI33xp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .A3(n_758), .B1(n_761), .B2(n_764), .B3(n_769), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
BUFx3_ASAP7_75t_L g853 ( .A(n_759), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_760), .A2(n_852), .B1(n_853), .B2(n_854), .Y(n_851) );
OAI221xp5_ASAP7_75t_L g1040 ( .A1(n_760), .A2(n_1004), .B1(n_1011), .B2(n_1041), .C(n_1043), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_763), .A2(n_856), .B1(n_858), .B2(n_859), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g1185 ( .A1(n_763), .A2(n_1148), .B1(n_1186), .B2(n_1187), .C(n_1188), .Y(n_1185) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g860 ( .A(n_765), .Y(n_860) );
INVx3_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx3_ASAP7_75t_L g1195 ( .A(n_766), .Y(n_1195) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g1344 ( .A(n_768), .Y(n_1344) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_770), .A2(n_847), .B1(n_862), .B2(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g1122 ( .A(n_772), .Y(n_1122) );
OAI31xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .A3(n_787), .B(n_793), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_782), .B2(n_784), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_781), .A2(n_804), .B1(n_806), .B2(n_808), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_782), .A2(n_823), .B1(n_833), .B2(n_834), .Y(n_832) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g1109 ( .A(n_783), .Y(n_1109) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g831 ( .A(n_786), .Y(n_831) );
INVx3_ASAP7_75t_L g1106 ( .A(n_786), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
BUFx2_ASAP7_75t_L g836 ( .A(n_789), .Y(n_836) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_SL g1111 ( .A(n_791), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_791), .A2(n_1085), .B1(n_1210), .B2(n_1212), .Y(n_1223) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g839 ( .A(n_792), .Y(n_839) );
INVx1_ASAP7_75t_L g928 ( .A(n_792), .Y(n_928) );
OAI31xp33_ASAP7_75t_L g826 ( .A1(n_793), .A2(n_827), .A3(n_835), .B(n_840), .Y(n_826) );
OAI31xp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_800), .A3(n_809), .B(n_813), .Y(n_794) );
INVx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_797), .A2(n_799), .B1(n_1173), .B2(n_1174), .Y(n_1179) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g820 ( .A(n_799), .Y(n_820) );
INVx2_ASAP7_75t_L g1103 ( .A(n_799), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g1200 ( .A1(n_799), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_799), .A2(n_1202), .B1(n_1257), .B2(n_1258), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_804), .A2(n_806), .B1(n_823), .B2(n_824), .Y(n_822) );
BUFx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_807), .A2(n_935), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
INVx1_ASAP7_75t_L g1269 ( .A(n_807), .Y(n_1269) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
OAI31xp33_ASAP7_75t_L g818 ( .A1(n_813), .A2(n_819), .A3(n_821), .B(n_825), .Y(n_818) );
BUFx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g1020 ( .A1(n_814), .A2(n_1021), .B(n_1031), .Y(n_1020) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_814), .A2(n_1113), .B1(n_1199), .B2(n_1214), .C(n_1224), .Y(n_1198) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_826), .C(n_842), .Y(n_817) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_830), .A2(n_1124), .B1(n_1130), .B2(n_1141), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_830), .A2(n_1120), .B1(n_1134), .B2(n_1141), .Y(n_1142) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_833), .A2(n_922), .B1(n_923), .B2(n_924), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_833), .A2(n_1100), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_838), .A2(n_1085), .B1(n_1163), .B2(n_1164), .C(n_1165), .Y(n_1162) );
INVx2_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_864), .Y(n_842) );
OAI33xp33_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .A3(n_851), .B1(n_855), .B2(n_860), .B3(n_861), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_844), .A2(n_860), .B1(n_1032), .B2(n_1040), .Y(n_1031) );
OAI22xp33_ASAP7_75t_L g1184 ( .A1(n_844), .A2(n_1185), .B1(n_1190), .B2(n_1193), .Y(n_1184) );
OAI22xp33_ASAP7_75t_L g845 ( .A1(n_846), .A2(n_847), .B1(n_848), .B2(n_849), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_848), .A2(n_863), .B1(n_869), .B2(n_874), .Y(n_873) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx3_ASAP7_75t_L g950 ( .A(n_850), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_852), .A2(n_858), .B1(n_869), .B2(n_871), .Y(n_868) );
INVx2_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx4_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g874 ( .A(n_872), .Y(n_874) );
INVx2_ASAP7_75t_L g912 ( .A(n_872), .Y(n_912) );
INVx2_ASAP7_75t_L g967 ( .A(n_872), .Y(n_967) );
INVx1_ASAP7_75t_L g1007 ( .A(n_872), .Y(n_1007) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
XNOR2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_983), .Y(n_880) );
XNOR2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_944), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_918), .C(n_931), .Y(n_883) );
NOR2xp33_ASAP7_75t_SL g884 ( .A(n_885), .B(n_905), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_888), .A2(n_904), .B1(n_910), .B2(n_912), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B1(n_894), .B2(n_896), .Y(n_890) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_891), .A2(n_898), .B1(n_910), .B2(n_912), .Y(n_909) );
INVx2_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
INVx3_ASAP7_75t_L g1055 ( .A(n_893), .Y(n_1055) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_893), .Y(n_1129) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g914 ( .A1(n_896), .A2(n_901), .B1(n_908), .B2(n_915), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_899), .A2(n_1041), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g1128 ( .A1(n_899), .A2(n_1129), .B1(n_1130), .B2(n_1131), .Y(n_1128) );
BUFx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
OR2x2_ASAP7_75t_L g1340 ( .A(n_900), .B(n_1341), .Y(n_1340) );
OAI33xp33_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_907), .A3(n_909), .B1(n_913), .B2(n_914), .B3(n_917), .Y(n_905) );
OAI33xp33_ASAP7_75t_L g1062 ( .A1(n_906), .A2(n_917), .A3(n_1063), .B1(n_1064), .B2(n_1065), .B3(n_1067), .Y(n_1062) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_908), .A2(n_954), .B1(n_957), .B2(n_963), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_908), .A2(n_963), .B1(n_1049), .B2(n_1060), .Y(n_1063) );
INVx2_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g1066 ( .A(n_911), .Y(n_1066) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
OAI31xp33_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_926), .A3(n_929), .B(n_930), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_920), .A2(n_966), .B1(n_1052), .B2(n_1056), .Y(n_1064) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
NAND2xp5_ASAP7_75t_SL g998 ( .A(n_928), .B(n_999), .Y(n_998) );
OAI31xp33_ASAP7_75t_SL g931 ( .A1(n_932), .A2(n_933), .A3(n_942), .B(n_943), .Y(n_931) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1365 ( .A(n_938), .Y(n_1365) );
AND2x4_ASAP7_75t_SL g1360 ( .A(n_939), .B(n_1361), .Y(n_1360) );
INVx3_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
OAI31xp33_ASAP7_75t_SL g976 ( .A1(n_943), .A2(n_977), .A3(n_978), .B(n_979), .Y(n_976) );
OAI21xp5_ASAP7_75t_L g1069 ( .A1(n_943), .A2(n_1070), .B(n_1076), .Y(n_1069) );
NAND3xp33_ASAP7_75t_L g945 ( .A(n_946), .B(n_969), .C(n_976), .Y(n_945) );
NOR2xp33_ASAP7_75t_SL g946 ( .A(n_947), .B(n_961), .Y(n_946) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_951), .A2(n_960), .B1(n_966), .B2(n_967), .Y(n_965) );
XOR2xp5_ASAP7_75t_L g983 ( .A(n_984), .B(n_1044), .Y(n_983) );
OAI21xp5_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_1018), .B(n_1020), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1006), .B(n_1010), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1003), .B1(n_1004), .B2(n_1005), .Y(n_1001) );
OAI211xp5_ASAP7_75t_SL g1010 ( .A1(n_1011), .A2(n_1012), .B(n_1013), .C(n_1016), .Y(n_1010) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1015), .Y(n_1316) );
INVx2_ASAP7_75t_L g1336 ( .A(n_1018), .Y(n_1336) );
BUFx2_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
NAND2xp5_ASAP7_75t_SL g1021 ( .A(n_1022), .B(n_1028), .Y(n_1021) );
OAI211xp5_ASAP7_75t_L g1032 ( .A1(n_1033), .A2(n_1034), .B(n_1036), .C(n_1038), .Y(n_1032) );
INVx2_ASAP7_75t_SL g1034 ( .A(n_1035), .Y(n_1034) );
AND2x4_ASAP7_75t_L g1380 ( .A(n_1037), .B(n_1361), .Y(n_1380) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx3_ASAP7_75t_L g1126 ( .A(n_1042), .Y(n_1126) );
NAND3xp33_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1069), .C(n_1079), .Y(n_1045) );
NOR2xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1062), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_1057), .A2(n_1124), .B1(n_1125), .B2(n_1127), .Y(n_1123) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_1078), .A2(n_1163), .B1(n_1164), .B2(n_1181), .Y(n_1180) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_1084), .A2(n_1085), .B1(n_1086), .B2(n_1087), .Y(n_1083) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_1091), .A2(n_1092), .B1(n_1196), .B2(n_1197), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
XNOR2xp5_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1144), .Y(n_1093) );
NAND3xp33_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1104), .C(n_1114), .Y(n_1095) );
OAI31xp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1110), .A3(n_1112), .B(n_1113), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1135), .Y(n_1114) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1118), .B1(n_1120), .B2(n_1121), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_1117), .A2(n_1133), .B1(n_1137), .B2(n_1139), .Y(n_1136) );
BUFx4f_ASAP7_75t_SL g1118 ( .A(n_1119), .Y(n_1118) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_1122), .Y(n_1121) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1126), .B(n_1377), .Y(n_1379) );
INVx2_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
NOR4xp25_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1161), .C(n_1175), .D(n_1184), .Y(n_1145) );
OAI22xp33_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1152), .B1(n_1153), .B2(n_1160), .Y(n_1146) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
AND2x4_ASAP7_75t_L g1320 ( .A(n_1159), .B(n_1307), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
AOI31xp33_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1179), .A3(n_1180), .B(n_1183), .Y(n_1175) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
AO21x1_ASAP7_75t_L g1265 ( .A1(n_1183), .A2(n_1266), .B(n_1271), .Y(n_1265) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1186), .Y(n_1286) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
BUFx2_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1244 ( .A(n_1195), .Y(n_1244) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
NAND3xp33_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1204), .C(n_1209), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1211), .B1(n_1212), .B2(n_1213), .Y(n_1209) );
NAND3xp33_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1217), .C(n_1223), .Y(n_1214) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NAND4xp25_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1234), .C(n_1237), .D(n_1242), .Y(n_1224) );
NAND3xp33_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1231), .C(n_1233), .Y(n_1225) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1323 ( .A(n_1229), .Y(n_1323) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .C(n_1245), .Y(n_1242) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
BUFx2_ASAP7_75t_L g1283 ( .A(n_1248), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
NAND4xp75_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1265), .C(n_1272), .D(n_1281), .Y(n_1254) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1260), .B(n_1264), .Y(n_1259) );
INVx2_ASAP7_75t_SL g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
CKINVDCx5p33_ASAP7_75t_R g1293 ( .A(n_1294), .Y(n_1293) );
HB1xp67_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
BUFx3_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1300), .Y(n_1381) );
NAND3xp33_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1337), .C(n_1357), .Y(n_1300) );
OAI21xp5_ASAP7_75t_SL g1301 ( .A1(n_1302), .A2(n_1318), .B(n_1336), .Y(n_1301) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx4_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1312), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1310), .B(n_1311), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1359 ( .A1(n_1312), .A2(n_1360), .B1(n_1362), .B2(n_1363), .Y(n_1359) );
INVx3_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
AOI21xp5_ASAP7_75t_L g1321 ( .A1(n_1322), .A2(n_1325), .B(n_1327), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_1329), .A2(n_1330), .B1(n_1333), .B2(n_1334), .Y(n_1328) );
INVx2_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
BUFx6f_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
AOI21xp5_ASAP7_75t_L g1337 ( .A1(n_1338), .A2(n_1346), .B(n_1347), .Y(n_1337) );
INVx8_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
AND2x4_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1343), .Y(n_1339) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1341), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1345), .Y(n_1343) );
AND2x4_ASAP7_75t_L g1361 ( .A(n_1344), .B(n_1354), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1348 ( .A(n_1349), .B(n_1350), .Y(n_1348) );
OR2x6_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1356), .Y(n_1352) );
NOR3xp33_ASAP7_75t_L g1357 ( .A(n_1358), .B(n_1374), .C(n_1380), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1366), .Y(n_1358) );
AND2x4_ASAP7_75t_SL g1363 ( .A(n_1361), .B(n_1364), .Y(n_1363) );
INVx2_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
INVxp67_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx2_ASAP7_75t_SL g1378 ( .A(n_1379), .Y(n_1378) );
INVx3_ASAP7_75t_L g1382 ( .A(n_1383), .Y(n_1382) );
INVxp67_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
endmodule