module fake_jpeg_19759_n_296 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_296);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_10),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_39),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_0),
.C(n_1),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_14),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_33),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_49),
.A2(n_17),
.B1(n_32),
.B2(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_51),
.A2(n_55),
.B1(n_64),
.B2(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_52),
.B(n_70),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_17),
.B1(n_32),
.B2(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_39),
.B1(n_48),
.B2(n_32),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_56),
.A2(n_60),
.B1(n_82),
.B2(n_83),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_17),
.B1(n_15),
.B2(n_26),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_25),
.B1(n_18),
.B2(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_67),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_75),
.Y(n_113)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_19),
.B1(n_30),
.B2(n_22),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_73),
.Y(n_129)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_77),
.B(n_79),
.Y(n_118)
);

CKINVDCx12_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_80),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_24),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_15),
.B1(n_26),
.B2(n_27),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_34),
.B1(n_33),
.B2(n_21),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_86),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_93),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_16),
.B1(n_23),
.B2(n_33),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_21),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_38),
.B(n_27),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_97),
.Y(n_126)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_49),
.A2(n_23),
.B1(n_34),
.B2(n_27),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_29),
.B1(n_25),
.B2(n_35),
.Y(n_128)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_59),
.B(n_18),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_53),
.C(n_72),
.Y(n_139)
);

NAND2x1_ASAP7_75t_L g102 ( 
.A(n_59),
.B(n_25),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_51),
.B(n_92),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_70),
.A2(n_29),
.B(n_18),
.C(n_25),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_104),
.A2(n_116),
.B(n_126),
.Y(n_157)
);

OR2x2_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_18),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g146 ( 
.A1(n_119),
.A2(n_99),
.B(n_95),
.Y(n_146)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_84),
.B(n_34),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_76),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_23),
.B1(n_29),
.B2(n_18),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_125),
.A2(n_128),
.B1(n_130),
.B2(n_55),
.Y(n_136)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_133),
.B(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_129),
.A2(n_57),
.B(n_64),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_143),
.B(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_124),
.A2(n_64),
.B1(n_71),
.B2(n_88),
.Y(n_137)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_125),
.B(n_116),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_12),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_155),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_161),
.Y(n_166)
);

INVx5_ASAP7_75t_SL g141 ( 
.A(n_120),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_145),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_159),
.C(n_103),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_129),
.A2(n_81),
.B1(n_71),
.B2(n_58),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

XOR2x1_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_115),
.Y(n_194)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_53),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_81),
.B1(n_74),
.B2(n_85),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_94),
.B1(n_69),
.B2(n_76),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_102),
.A2(n_92),
.B(n_90),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_111),
.A2(n_69),
.B1(n_90),
.B2(n_91),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_101),
.B(n_62),
.C(n_35),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_160),
.B(n_100),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_102),
.A2(n_1),
.B(n_2),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_130),
.B1(n_118),
.B2(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_6),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_109),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_122),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_174),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_179),
.B(n_180),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_104),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_155),
.C(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_186),
.B1(n_141),
.B2(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_185),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_104),
.B1(n_118),
.B2(n_115),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_122),
.B(n_114),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_132),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_184),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_107),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_136),
.A2(n_108),
.B1(n_107),
.B2(n_120),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_6),
.C(n_8),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_188),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_138),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_123),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_189),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_192),
.A2(n_194),
.B(n_149),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_140),
.B(n_108),
.Y(n_195)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_201),
.C(n_206),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_199),
.A2(n_202),
.B(n_213),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_150),
.C(n_154),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_168),
.A2(n_137),
.B(n_134),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_182),
.A2(n_137),
.B1(n_152),
.B2(n_144),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_210),
.B1(n_212),
.B2(n_186),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_147),
.C(n_161),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_176),
.B(n_162),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_214),
.Y(n_233)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_173),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_151),
.B1(n_148),
.B2(n_141),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_100),
.B(n_117),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_131),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_194),
.B(n_179),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_232),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_169),
.B(n_192),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_229),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_185),
.C(n_177),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_231),
.C(n_234),
.Y(n_245)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_177),
.B(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_196),
.B(n_188),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_227),
.B(n_172),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_230),
.B1(n_204),
.B2(n_203),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_198),
.A2(n_177),
.B(n_166),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_211),
.B(n_205),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_166),
.C(n_195),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g232 ( 
.A1(n_205),
.A2(n_178),
.B1(n_172),
.B2(n_174),
.C(n_183),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_193),
.C(n_190),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_193),
.C(n_190),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_213),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

BUFx12f_ASAP7_75t_SL g238 ( 
.A(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_238),
.A2(n_220),
.B(n_229),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_244),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_215),
.B1(n_203),
.B2(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_242),
.B1(n_252),
.B2(n_228),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_211),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_223),
.B(n_196),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_237),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_215),
.B1(n_217),
.B2(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_221),
.C(n_234),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_260),
.C(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_257),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_238),
.A2(n_158),
.B1(n_208),
.B2(n_218),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_255),
.A2(n_249),
.B1(n_184),
.B2(n_250),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_241),
.B(n_230),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_258),
.B(n_263),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_221),
.C(n_235),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_233),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_244),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_181),
.Y(n_263)
);

AOI31xp67_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_218),
.A3(n_231),
.B(n_220),
.Y(n_264)
);

AOI321xp33_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_219),
.A3(n_200),
.B1(n_209),
.B2(n_164),
.C(n_171),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_243),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_268),
.C(n_262),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_273),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_253),
.C(n_256),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_274),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_249),
.B1(n_252),
.B2(n_164),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_259),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_256),
.Y(n_276)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_276),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_280),
.Y(n_286)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_265),
.B(n_248),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_158),
.B(n_115),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_275),
.Y(n_290)
);

NOR4xp25_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_278),
.C(n_277),
.D(n_270),
.Y(n_288)
);

OAI21xp33_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_290),
.B(n_291),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_287),
.C(n_106),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_6),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_106),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_287),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_295),
.Y(n_296)
);


endmodule