module fake_jpeg_15186_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_65),
.Y(n_88)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_52),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_81),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_54),
.B1(n_60),
.B2(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_49),
.B1(n_50),
.B2(n_2),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_87),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_93),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_95),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_44),
.A3(n_63),
.B1(n_59),
.B2(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_98),
.B(n_58),
.Y(n_121)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_83),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_0),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_62),
.B1(n_64),
.B2(n_3),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_64),
.B1(n_1),
.B2(n_3),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_107),
.B(n_108),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_99),
.B(n_51),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_122),
.C(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_5),
.C(n_7),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_126),
.B(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_127),
.B(n_129),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_125),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_112),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_111),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_140),
.A2(n_116),
.B1(n_113),
.B2(n_120),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_106),
.B(n_90),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_142),
.C(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_143),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_150),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_147),
.B(n_9),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g153 ( 
.A(n_152),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_8),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_11),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_155),
.B(n_13),
.Y(n_156)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_14),
.B(n_15),
.Y(n_157)
);

OAI311xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_17),
.A3(n_18),
.B1(n_19),
.C1(n_20),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_21),
.B(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_24),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_26),
.B(n_29),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_32),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_34),
.Y(n_163)
);


endmodule