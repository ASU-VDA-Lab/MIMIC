module real_jpeg_3394_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_4),
.A2(n_30),
.B1(n_32),
.B2(n_56),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_5),
.A2(n_30),
.B1(n_32),
.B2(n_59),
.Y(n_99)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_7),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_34),
.B1(n_50),
.B2(n_51),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_7),
.B(n_25),
.C(n_38),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_7),
.B(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_7),
.B(n_23),
.C(n_30),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_7),
.B(n_51),
.C(n_62),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_7),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_54),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_7),
.B(n_61),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_106),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_104),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_86),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_14),
.B(n_86),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_68),
.C(n_78),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_15),
.A2(n_16),
.B1(n_68),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_46),
.B2(n_67),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_17),
.A2(n_18),
.B1(n_112),
.B2(n_118),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_17),
.A2(n_18),
.B1(n_81),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_35),
.B2(n_45),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_19),
.B(n_45),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_19),
.A2(n_20),
.B1(n_60),
.B2(n_120),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_19),
.A2(n_20),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_19),
.A2(n_60),
.B(n_124),
.C(n_190),
.Y(n_193)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_35),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_20),
.A2(n_96),
.B(n_100),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_20),
.B(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_120),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_20),
.B(n_117),
.C(n_143),
.Y(n_142)
);

AO21x2_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_29),
.B(n_33),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_22)
);

INVx3_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

OA22x2_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_24),
.A2(n_25),
.B1(n_38),
.B2(n_42),
.Y(n_43)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_25),
.B(n_158),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_29),
.Y(n_175)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_30),
.A2(n_32),
.B1(n_62),
.B2(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_30),
.B(n_169),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_35),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_35),
.A2(n_45),
.B1(n_69),
.B2(n_77),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_35),
.A2(n_45),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

AO21x2_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_44),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_40),
.B(n_115),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_43),
.Y(n_144)
);

AOI211xp5_ASAP7_75t_SL g123 ( 
.A1(n_45),
.A2(n_60),
.B(n_85),
.C(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_46),
.A2(n_80),
.B(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_60),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_47),
.A2(n_60),
.B1(n_120),
.B2(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_47),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_48),
.A2(n_55),
.B1(n_57),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_51),
.B(n_180),
.Y(n_179)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_60),
.A2(n_82),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_60),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_60),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_60),
.A2(n_120),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_60),
.A2(n_120),
.B1(n_167),
.B2(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_60),
.A2(n_120),
.B1(n_155),
.B2(n_196),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B(n_66),
.Y(n_60)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_64),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_68),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_72),
.B2(n_77),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_83),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_78),
.A2(n_79),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B(n_84),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_84),
.B(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_94),
.B2(n_95),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI21x1_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_199),
.B(n_205),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_146),
.Y(n_107)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_132),
.B(n_145),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_147),
.C(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_125),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_125),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.C(n_122),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_117),
.B1(n_143),
.B2(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_117),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_116),
.A2(n_117),
.B1(n_156),
.B2(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_117),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_117),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_117),
.B(n_120),
.C(n_174),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_151),
.C(n_155),
.Y(n_150)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_128),
.C(n_130),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_136),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.C(n_142),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_138),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_139),
.A2(n_140),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_162),
.B(n_198),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_159),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_159),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_155),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_192),
.B(n_197),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_186),
.B(n_191),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_176),
.B(n_185),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_170),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_194),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_200),
.B(n_201),
.Y(n_205)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);


endmodule