module fake_jpeg_23045_n_318 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_27),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_39),
.CON(n_50),
.SN(n_50)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.Y(n_57)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_24),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_31),
.B(n_19),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_67),
.B(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_22),
.B1(n_33),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_59),
.B1(n_66),
.B2(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_33),
.B1(n_34),
.B2(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_64),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_22),
.B1(n_32),
.B2(n_28),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_67)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_21),
.B1(n_19),
.B2(n_28),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_32),
.B1(n_19),
.B2(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_37),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_74),
.B(n_8),
.C(n_15),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_35),
.B1(n_24),
.B2(n_26),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_76),
.A2(n_92),
.B1(n_98),
.B2(n_100),
.Y(n_121)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_107),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_35),
.B1(n_26),
.B2(n_20),
.Y(n_92)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_102),
.Y(n_134)
);

INVx2_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_97),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_39),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_46),
.A2(n_20),
.B1(n_34),
.B2(n_23),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_10),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_41),
.B1(n_29),
.B2(n_23),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_46),
.A2(n_60),
.B1(n_56),
.B2(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_0),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_10),
.C(n_15),
.Y(n_123)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_8),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_128),
.Y(n_159)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_60),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_117),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_116),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_75),
.Y(n_117)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_120),
.A2(n_125),
.B1(n_4),
.B2(n_5),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_126),
.B1(n_94),
.B2(n_82),
.Y(n_146)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_8),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_83),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_4),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_99),
.A2(n_2),
.B(n_4),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_81),
.B(n_73),
.Y(n_143)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_84),
.C(n_78),
.Y(n_162)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_138),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_121),
.A2(n_99),
.B1(n_85),
.B2(n_91),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_146),
.B1(n_157),
.B2(n_167),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_130),
.B(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_150),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_91),
.B1(n_105),
.B2(n_73),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_149),
.B1(n_154),
.B2(n_155),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_105),
.B1(n_82),
.B2(n_79),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_87),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_162),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_80),
.B1(n_78),
.B2(n_77),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_109),
.A2(n_95),
.B1(n_89),
.B2(n_88),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_88),
.B1(n_103),
.B2(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_124),
.B(n_84),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_103),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_164),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_86),
.B(n_77),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_166),
.B(n_137),
.Y(n_176)
);

NAND2x1_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_5),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_173),
.B(n_177),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_176),
.A2(n_199),
.B(n_202),
.Y(n_228)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_189),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_191),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_149),
.B1(n_141),
.B2(n_118),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_187),
.B1(n_194),
.B2(n_158),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_128),
.B1(n_110),
.B2(n_122),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_195),
.B1(n_154),
.B2(n_138),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_126),
.B1(n_122),
.B2(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_166),
.B(n_122),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_159),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_120),
.B1(n_111),
.B2(n_114),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_111),
.B1(n_136),
.B2(n_112),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_114),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_154),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_143),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_129),
.B(n_132),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_114),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_170),
.A2(n_5),
.B(n_6),
.Y(n_202)
);

XNOR2x2_ASAP7_75t_SL g204 ( 
.A(n_191),
.B(n_159),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_225),
.B(n_227),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_206),
.B1(n_216),
.B2(n_217),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_150),
.B1(n_153),
.B2(n_158),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_156),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_209),
.C(n_215),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_218),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_132),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_214),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_140),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_187),
.B1(n_198),
.B2(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_148),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_154),
.B1(n_111),
.B2(n_125),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_194),
.B1(n_216),
.B2(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_193),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_192),
.B(n_182),
.C(n_176),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_226),
.C(n_182),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_125),
.Y(n_226)
);

OR2x2_ASAP7_75t_SL g227 ( 
.A(n_199),
.B(n_7),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_203),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_230),
.B(n_241),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_208),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_233),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_237),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_171),
.B(n_199),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_249),
.C(n_229),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_195),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_213),
.A2(n_171),
.B1(n_188),
.B2(n_184),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_248),
.B1(n_220),
.B2(n_225),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_243),
.A2(n_247),
.B1(n_250),
.B2(n_222),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_246),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_211),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_183),
.B1(n_174),
.B2(n_190),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_185),
.C(n_174),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_227),
.B(n_226),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_232),
.B(n_237),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_254),
.B(n_243),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_186),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_266),
.C(n_242),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_203),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_259),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_215),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_228),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_248),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_200),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_223),
.B1(n_222),
.B2(n_228),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_265),
.A2(n_236),
.B1(n_244),
.B2(n_245),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_249),
.C(n_250),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_236),
.B1(n_233),
.B2(n_234),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_272),
.Y(n_283)
);

AOI321xp33_ASAP7_75t_L g286 ( 
.A1(n_270),
.A2(n_261),
.A3(n_260),
.B1(n_196),
.B2(n_202),
.C(n_185),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_235),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_247),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_278),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_256),
.C(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_186),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_197),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_282),
.A2(n_266),
.B1(n_257),
.B2(n_259),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_270),
.B(n_265),
.CI(n_254),
.CON(n_284),
.SN(n_284)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_285),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_268),
.CI(n_262),
.CON(n_285),
.SN(n_285)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_276),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_258),
.B(n_256),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_293),
.B(n_16),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_6),
.C(n_288),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_277),
.A2(n_5),
.B1(n_6),
.B2(n_12),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_283),
.CI(n_285),
.CON(n_309),
.SN(n_309)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_294),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_294),
.B(n_272),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_299),
.B(n_300),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_279),
.B(n_16),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_279),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_303),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_292),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

AOI31xp33_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_286),
.A3(n_290),
.B(n_284),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_309),
.B(n_283),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_304),
.B(n_308),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_313),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_314),
.B(n_292),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_284),
.Y(n_318)
);


endmodule