module fake_jpeg_6072_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVxp33_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_57),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_28),
.B1(n_36),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_52),
.B1(n_58),
.B2(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_60),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_28),
.B1(n_35),
.B2(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_13),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_46),
.B(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_46),
.B(n_13),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_66),
.Y(n_77)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_28),
.B1(n_35),
.B2(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_41),
.A2(n_26),
.B1(n_20),
.B2(n_23),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_65),
.B1(n_19),
.B2(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_64),
.B(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_21),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_29),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_70),
.A2(n_82),
.B(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_74),
.B1(n_83),
.B2(n_49),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_44),
.B1(n_39),
.B2(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_80),
.B1(n_57),
.B2(n_60),
.Y(n_88)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_66),
.A2(n_44),
.B1(n_39),
.B2(n_29),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_82),
.A2(n_61),
.B1(n_56),
.B2(n_63),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_29),
.B1(n_36),
.B2(n_34),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_89),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_99),
.B1(n_100),
.B2(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_64),
.C(n_40),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_92),
.C(n_72),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_66),
.C(n_49),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_97),
.B1(n_68),
.B2(n_78),
.Y(n_105)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_102),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_55),
.B1(n_62),
.B2(n_60),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_77),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_77),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_55),
.B1(n_62),
.B2(n_34),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_84),
.A2(n_55),
.B1(n_36),
.B2(n_30),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_77),
.B(n_67),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_115),
.B1(n_19),
.B2(n_23),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_98),
.B(n_70),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_110),
.C(n_31),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_94),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_112),
.B(n_116),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_125),
.B(n_121),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_86),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_74),
.B1(n_79),
.B2(n_75),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_80),
.B1(n_104),
.B2(n_76),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_122),
.B(n_19),
.Y(n_147)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_125),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_97),
.A2(n_30),
.B1(n_76),
.B2(n_42),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_96),
.B1(n_89),
.B2(n_103),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_23),
.B(n_20),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_104),
.B(n_21),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_101),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_124),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_91),
.B1(n_90),
.B2(n_92),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_145),
.B1(n_25),
.B2(n_17),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_139),
.B1(n_147),
.B2(n_112),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_140),
.C(n_106),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_18),
.B(n_17),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_22),
.B1(n_17),
.B2(n_25),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_31),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_166),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_111),
.B1(n_119),
.B2(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_168),
.C(n_170),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_152),
.A2(n_154),
.B1(n_155),
.B2(n_156),
.Y(n_183)
);

AOI22x1_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_124),
.B1(n_122),
.B2(n_120),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_135),
.A2(n_110),
.B1(n_109),
.B2(n_123),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_114),
.B1(n_25),
.B2(n_24),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_31),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_148),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_135),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_167),
.B1(n_171),
.B2(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_127),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_132),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_130),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_129),
.C(n_126),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_133),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_31),
.C(n_30),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_25),
.B1(n_24),
.B2(n_22),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_18),
.B1(n_17),
.B2(n_16),
.Y(n_172)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_172),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_16),
.B1(n_15),
.B2(n_42),
.Y(n_173)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_175),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_161),
.A2(n_138),
.B1(n_141),
.B2(n_137),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_176),
.A2(n_160),
.B1(n_162),
.B2(n_164),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_179),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_16),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_128),
.C(n_144),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_189),
.C(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_155),
.B(n_131),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_158),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_147),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_195),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_139),
.C(n_145),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_14),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_132),
.C(n_31),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_15),
.B1(n_16),
.B2(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_193),
.A2(n_172),
.B1(n_153),
.B2(n_166),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_16),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_177),
.A2(n_154),
.B(n_167),
.C(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_189),
.B(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_201),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_212),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_8),
.B(n_12),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_204),
.A2(n_21),
.B(n_7),
.Y(n_226)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_209),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_16),
.C(n_14),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_211),
.C(n_215),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_176),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_14),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_198),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_14),
.C(n_0),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_216),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_184),
.C(n_179),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_227),
.C(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_194),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_186),
.B1(n_195),
.B2(n_178),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_224),
.A2(n_226),
.B1(n_204),
.B2(n_211),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_232),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_205),
.C(n_213),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_21),
.B1(n_7),
.B2(n_2),
.Y(n_242)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_205),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_241),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_220),
.B(n_223),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_239),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_246),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_240),
.C(n_217),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_208),
.C(n_200),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_7),
.Y(n_241)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_6),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_221),
.B(n_222),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_5),
.B1(n_11),
.B2(n_2),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_8),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_229),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_254),
.B(n_255),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_256),
.C(n_251),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_219),
.B(n_224),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_8),
.Y(n_255)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_237),
.Y(n_256)
);

AOI21x1_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_233),
.B(n_5),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_240),
.A2(n_5),
.B1(n_11),
.B2(n_3),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_238),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_264),
.B(n_9),
.Y(n_275)
);

NAND2x1_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_4),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_253),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_3),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_269),
.B(n_259),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_281)
);

OAI321xp33_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_273),
.A3(n_267),
.B1(n_10),
.B2(n_12),
.C(n_1),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_4),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_4),
.B(n_9),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_277),
.C(n_9),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_262),
.B(n_9),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_279),
.B(n_280),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_266),
.B(n_267),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_10),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_281),
.C(n_0),
.Y(n_285)
);

OAI21x1_ASAP7_75t_SL g286 ( 
.A1(n_285),
.A2(n_283),
.B(n_0),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_0),
.B1(n_1),
.B2(n_242),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_287),
.B(n_1),
.Y(n_288)
);


endmodule