module fake_jpeg_24912_n_38 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_38);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_38;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx6_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_1),
.C(n_2),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_21),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_25),
.A2(n_18),
.B1(n_10),
.B2(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_8),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_20),
.B(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_18),
.B1(n_3),
.B2(n_6),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_31),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_32),
.C(n_30),
.Y(n_35)
);

AOI31xp67_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_34),
.A3(n_29),
.B(n_13),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B1(n_12),
.B2(n_16),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_9),
.Y(n_38)
);


endmodule