module fake_jpeg_9206_n_147 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_147);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_20),
.Y(n_30)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_13),
.B(n_15),
.C(n_22),
.Y(n_45)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_46),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_28),
.B1(n_25),
.B2(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_26),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_48),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_14),
.B1(n_25),
.B2(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_14),
.B1(n_25),
.B2(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_32),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_SL g57 ( 
.A(n_42),
.B(n_45),
.C(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_62),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_46),
.B(n_31),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_38),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_50),
.B1(n_37),
.B2(n_35),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_64),
.B1(n_52),
.B2(n_58),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_61),
.B1(n_63),
.B2(n_37),
.Y(n_84)
);

XNOR2x1_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_24),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_24),
.C(n_23),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_31),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_61),
.B(n_54),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_0),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_36),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_47),
.B1(n_36),
.B2(n_37),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_95),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_87),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_63),
.B(n_51),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_94),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_24),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_73),
.C(n_23),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_66),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_70),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_102),
.B1(n_105),
.B2(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_101),
.C(n_107),
.Y(n_110)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_71),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_91),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_85),
.B1(n_82),
.B2(n_88),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_113),
.A2(n_104),
.B1(n_101),
.B2(n_98),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_94),
.C(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_92),
.C(n_88),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_80),
.C(n_12),
.Y(n_117)
);

BUFx12_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_111),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_103),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_123),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_125),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_23),
.C(n_21),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_124),
.C(n_38),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_21),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_118),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_129),
.C(n_130),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_21),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.C(n_11),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_9),
.Y(n_130)
);

AOI21x1_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_1),
.B(n_2),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_13),
.B(n_12),
.C(n_16),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_134),
.B(n_137),
.Y(n_138)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_131),
.C(n_16),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_1),
.CI(n_2),
.CON(n_143),
.SN(n_143)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_7),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_1),
.B(n_4),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_35),
.B1(n_2),
.B2(n_4),
.Y(n_142)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_143),
.A3(n_144),
.B1(n_5),
.B2(n_6),
.C1(n_18),
.C2(n_139),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_143),
.C(n_5),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_18),
.Y(n_147)
);


endmodule