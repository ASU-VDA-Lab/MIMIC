module real_jpeg_16686_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_249;
wire n_288;
wire n_78;
wire n_83;
wire n_166;
wire n_221;
wire n_176;
wire n_286;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_222;
wire n_19;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

AND2x2_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_0),
.B(n_32),
.Y(n_31)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_0),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_0),
.B(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_0),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_0),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_0),
.B(n_110),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_1),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_1),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_2),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_2),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_3),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_3),
.B(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_3),
.B(n_162),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_4),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_5),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_5),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_6),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_6),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_6),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_6),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_6),
.B(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_7),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_7),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_8),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_9),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_9),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_9),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_10),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_11),
.B(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_13),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g271 ( 
.A(n_13),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22x1_ASAP7_75t_SL g51 ( 
.A1(n_14),
.A2(n_15),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_14),
.B(n_179),
.Y(n_178)
);

AOI31xp33_ASAP7_75t_L g41 ( 
.A1(n_15),
.A2(n_42),
.A3(n_45),
.B(n_51),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_15),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_15),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_15),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_15),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_15),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_15),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_189),
.B1(n_287),
.B2(n_288),
.Y(n_17)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_18),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_R g18 ( 
.A(n_19),
.B(n_187),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_141),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_20),
.B(n_141),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_118),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_21),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_40),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_22),
.B(n_41),
.C(n_58),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.C(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_23),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_24),
.B(n_28),
.Y(n_202)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_24),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_24),
.A2(n_249),
.B1(n_250),
.B2(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_27),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_27),
.Y(n_210)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_31),
.A2(n_36),
.B1(n_37),
.B2(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_31),
.Y(n_199)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_58),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_49),
.Y(n_160)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_51),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_51),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_59),
.B(n_63),
.C(n_68),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_67),
.B(n_219),
.C(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g232 ( 
.A(n_68),
.B(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_70),
.Y(n_260)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_74),
.B(n_118),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_92),
.C(n_106),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_75),
.B(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_76),
.B(n_80),
.C(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_85),
.B1(n_86),
.B2(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_80),
.A2(n_91),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_80),
.B(n_254),
.C(n_258),
.Y(n_278)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_93),
.B(n_107),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_101),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_94),
.A2(n_101),
.B1(n_154),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2x1_ASAP7_75t_L g226 ( 
.A(n_98),
.B(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_101),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_113),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_138),
.Y(n_118)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_120),
.B(n_131),
.C(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_131),
.B1(n_136),
.B2(n_137),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_127),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_140),
.C(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_167),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_151),
.Y(n_155)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_166),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_183),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_189),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_282),
.B(n_286),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_229),
.B(n_281),
.Y(n_191)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_215),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_193),
.B(n_215),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_212),
.B2(n_213),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_196),
.B(n_201),
.C(n_212),
.Y(n_283)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.C(n_207),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_203),
.Y(n_217)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.C(n_225),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_216),
.B(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_226),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_221),
.Y(n_233)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21x1_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_245),
.B(n_280),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_231),
.B(n_243),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_241),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_235),
.B1(n_241),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_236),
.B(n_239),
.Y(n_255)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_268),
.Y(n_267)
);

AOI21x1_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_274),
.B(n_279),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_261),
.B(n_273),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_253),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_267),
.B(n_272),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_265),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2x1_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_278),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);


endmodule