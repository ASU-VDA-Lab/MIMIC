module fake_ibex_526_n_968 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_968);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_968;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_510;
wire n_193;
wire n_418;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_832;
wire n_798;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_899;
wire n_843;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_4),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_105),
.B(n_129),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_87),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_82),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_3),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_59),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_39),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_49),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_15),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_34),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_92),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_98),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_9),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_4),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_97),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_122),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_164),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_89),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_48),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_140),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_78),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_85),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_28),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_101),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_75),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_20),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_124),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_123),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_5),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_146),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_111),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_168),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_43),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_93),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_22),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_13),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_94),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_115),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_65),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_116),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_46),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_41),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_110),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_91),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_95),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_132),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_62),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_80),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_36),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_107),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_158),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_152),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_90),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_176),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_154),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_2),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_86),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_21),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_174),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_55),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_106),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_131),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_96),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_117),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_77),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_57),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_34),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_178),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_149),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_37),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_120),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_14),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_177),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_121),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_113),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_40),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_161),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_150),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_42),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_26),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_0),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_16),
.B(n_74),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_76),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_56),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_32),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_66),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_41),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_13),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_29),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_153),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_23),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_83),
.Y(n_302)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_197),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_202),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_202),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_180),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_202),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_280),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_205),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_240),
.B(n_3),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_278),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_200),
.Y(n_315)
);

AOI22x1_ASAP7_75t_SL g316 ( 
.A1(n_180),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_235),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_191),
.A2(n_88),
.B(n_175),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_287),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g322 ( 
.A(n_206),
.B(n_44),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_191),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_253),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_195),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

BUFx8_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_195),
.B(n_11),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_196),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_285),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_198),
.Y(n_333)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_206),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_246),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_260),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_234),
.B(n_12),
.Y(n_338)
);

BUFx8_ASAP7_75t_L g339 ( 
.A(n_260),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g341 ( 
.A(n_247),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_294),
.Y(n_342)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

CKINVDCx6p67_ASAP7_75t_R g344 ( 
.A(n_226),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_196),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_14),
.Y(n_346)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_294),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_247),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_179),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

BUFx8_ASAP7_75t_SL g351 ( 
.A(n_235),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_196),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_199),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_291),
.Y(n_354)
);

AND2x4_ASAP7_75t_L g355 ( 
.A(n_203),
.B(n_18),
.Y(n_355)
);

OAI22x1_ASAP7_75t_SL g356 ( 
.A1(n_291),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_219),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_268),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_185),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g360 ( 
.A(n_187),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_221),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_229),
.Y(n_362)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_196),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_255),
.B(n_19),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_184),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_289),
.B(n_23),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_236),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_186),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_297),
.B(n_24),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_298),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_299),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_301),
.B(n_24),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_226),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_311),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_346),
.B(n_188),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_330),
.Y(n_379)
);

AOI21x1_ASAP7_75t_L g380 ( 
.A1(n_320),
.A2(n_190),
.B(n_189),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_330),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_346),
.B(n_192),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_332),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_319),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g386 ( 
.A(n_308),
.B(n_225),
.C(n_213),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_344),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_L g388 ( 
.A(n_322),
.B(n_182),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_310),
.B(n_193),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_355),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_354),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_364),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_304),
.B(n_236),
.Y(n_396)
);

NAND2xp33_ASAP7_75t_L g397 ( 
.A(n_322),
.B(n_187),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_364),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_321),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_312),
.B(n_194),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

BUFx6f_ASAP7_75t_SL g403 ( 
.A(n_364),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_373),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_L g408 ( 
.A(n_322),
.B(n_216),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_344),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_309),
.B(n_204),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

NAND3x1_ASAP7_75t_L g413 ( 
.A(n_314),
.B(n_292),
.C(n_210),
.Y(n_413)
);

INVxp67_ASAP7_75t_R g414 ( 
.A(n_336),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_373),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_209),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_340),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_342),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_304),
.B(n_283),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_359),
.B(n_217),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_L g421 ( 
.A1(n_315),
.A2(n_233),
.B1(n_261),
.B2(n_265),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_305),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_L g424 ( 
.A(n_322),
.B(n_183),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_307),
.B(n_222),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_349),
.B(n_228),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_318),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_342),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_341),
.Y(n_430)
);

NOR2x1p5_ASAP7_75t_L g431 ( 
.A(n_303),
.B(n_315),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_323),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_324),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_324),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_359),
.B(n_231),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_232),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_329),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_369),
.B(n_237),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_303),
.A2(n_261),
.B1(n_233),
.B2(n_281),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_326),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_352),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_326),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_352),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_335),
.B(n_288),
.Y(n_448)
);

INVx6_ASAP7_75t_L g449 ( 
.A(n_329),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_358),
.B(n_288),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_360),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_366),
.B(n_238),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_337),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_368),
.Y(n_455)
);

NAND3xp33_ASAP7_75t_L g456 ( 
.A(n_339),
.B(n_262),
.C(n_236),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_339),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_360),
.B(n_279),
.Y(n_458)
);

AO22x2_ASAP7_75t_L g459 ( 
.A1(n_316),
.A2(n_276),
.B1(n_242),
.B2(n_244),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_354),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_353),
.B(n_245),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_369),
.B(n_248),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_368),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_357),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_322),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_334),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_334),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_370),
.A2(n_254),
.B(n_250),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_430),
.B(n_374),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_374),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_395),
.B(n_338),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

OR2x6_ASAP7_75t_L g478 ( 
.A(n_431),
.B(n_306),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_435),
.A2(n_372),
.B1(n_371),
.B2(n_365),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g480 ( 
.A1(n_380),
.A2(n_362),
.B(n_313),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_317),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_327),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_441),
.B(n_201),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_396),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_393),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_419),
.B(n_207),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_457),
.B(n_208),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_403),
.A2(n_348),
.B1(n_356),
.B2(n_257),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_211),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_212),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_468),
.B(n_214),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_416),
.B(n_215),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_416),
.B(n_218),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_421),
.B(n_351),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_SL g496 ( 
.A(n_449),
.B(n_220),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_440),
.B(n_286),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_223),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_384),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_381),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_452),
.B(n_224),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_381),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_399),
.A2(n_405),
.B1(n_415),
.B2(n_404),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_403),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_452),
.B(n_227),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_467),
.B(n_230),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_378),
.A2(n_271),
.B(n_259),
.C(n_263),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_393),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_386),
.B(n_239),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_390),
.Y(n_510)
);

INVx8_ASAP7_75t_L g511 ( 
.A(n_451),
.Y(n_511)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_390),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_392),
.B(n_267),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_422),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_458),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_471),
.B(n_379),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_382),
.B(n_243),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_471),
.B(n_273),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_462),
.A2(n_443),
.B1(n_410),
.B2(n_387),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_375),
.B(n_411),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_397),
.B(n_275),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_459),
.A2(n_351),
.B1(n_262),
.B2(n_236),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx2_ASAP7_75t_SL g525 ( 
.A(n_375),
.Y(n_525)
);

BUFx6f_ASAP7_75t_SL g526 ( 
.A(n_375),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_453),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_413),
.A2(n_391),
.B1(n_401),
.B2(n_411),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_377),
.B(n_249),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_448),
.B(n_251),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_383),
.A2(n_284),
.B1(n_300),
.B2(n_345),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_391),
.A2(n_262),
.B1(n_252),
.B2(n_272),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_426),
.B(n_256),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_444),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_426),
.B(n_258),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_401),
.B(n_264),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_463),
.B(n_266),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_463),
.B(n_269),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_462),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_456),
.B(n_270),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_425),
.B(n_282),
.Y(n_543)
);

BUFx12f_ASAP7_75t_SL g544 ( 
.A(n_459),
.Y(n_544)
);

O2A1O1Ixp33_ASAP7_75t_L g545 ( 
.A1(n_420),
.A2(n_439),
.B(n_442),
.C(n_464),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_446),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_425),
.B(n_296),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_420),
.B(n_331),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_439),
.B(n_331),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_469),
.Y(n_550)
);

OAI221xp5_ASAP7_75t_L g551 ( 
.A1(n_388),
.A2(n_363),
.B1(n_181),
.B2(n_347),
.C(n_28),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_470),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_424),
.B(n_347),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_433),
.B(n_25),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_L g555 ( 
.A1(n_517),
.A2(n_503),
.B(n_519),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_528),
.B(n_25),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_477),
.B(n_26),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_522),
.A2(n_465),
.B1(n_461),
.B2(n_455),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_472),
.B(n_27),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_510),
.B(n_433),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_499),
.B(n_27),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_498),
.B(n_455),
.C(n_454),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_517),
.A2(n_454),
.B1(n_447),
.B2(n_409),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_516),
.Y(n_564)
);

A2O1A1Ixp33_ASAP7_75t_L g565 ( 
.A1(n_482),
.A2(n_447),
.B(n_407),
.C(n_406),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_521),
.B(n_29),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_475),
.B(n_30),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_525),
.B(n_30),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_504),
.B(n_31),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_479),
.B(n_32),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_497),
.B(n_33),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_495),
.B(n_33),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_553),
.A2(n_513),
.B(n_518),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_479),
.B(n_35),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_512),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_511),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_515),
.B(n_35),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_524),
.A2(n_412),
.B1(n_394),
.B2(n_429),
.Y(n_578)
);

AOI21xp33_ASAP7_75t_L g579 ( 
.A1(n_505),
.A2(n_38),
.B(n_45),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_540),
.B(n_47),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_514),
.Y(n_581)
);

O2A1O1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_507),
.A2(n_429),
.B(n_427),
.C(n_423),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_531),
.B(n_50),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_473),
.Y(n_584)
);

OAI321xp33_ASAP7_75t_L g585 ( 
.A1(n_551),
.A2(n_412),
.A3(n_394),
.B1(n_427),
.B2(n_423),
.C(n_418),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_512),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_526),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_481),
.B(n_51),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_486),
.B(n_376),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_480),
.A2(n_402),
.B(n_398),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_500),
.Y(n_591)
);

OAI21xp33_ASAP7_75t_L g592 ( 
.A1(n_538),
.A2(n_418),
.B(n_400),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_533),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_539),
.B(n_538),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_539),
.B(n_52),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_501),
.B(n_53),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_480),
.A2(n_545),
.B(n_502),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_546),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_484),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_481),
.B(n_58),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_536),
.A2(n_417),
.B(n_385),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_543),
.B(n_60),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_488),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_547),
.B(n_61),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_493),
.B(n_494),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_490),
.B(n_63),
.Y(n_609)
);

OAI21xp33_ASAP7_75t_L g610 ( 
.A1(n_532),
.A2(n_535),
.B(n_537),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_529),
.A2(n_445),
.B(n_438),
.C(n_68),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_491),
.A2(n_492),
.B(n_530),
.Y(n_613)
);

AND2x2_ASAP7_75t_SL g614 ( 
.A(n_544),
.B(n_64),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_523),
.B(n_67),
.Y(n_615)
);

AO21x1_ASAP7_75t_L g616 ( 
.A1(n_554),
.A2(n_71),
.B(n_72),
.Y(n_616)
);

BUFx8_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_511),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_522),
.B(n_73),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_483),
.B(n_487),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_508),
.B(n_81),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_534),
.B(n_438),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_509),
.B(n_99),
.Y(n_624)
);

NOR3xp33_ASAP7_75t_L g625 ( 
.A(n_520),
.B(n_100),
.C(n_102),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_522),
.Y(n_626)
);

O2A1O1Ixp33_ASAP7_75t_SL g627 ( 
.A1(n_542),
.A2(n_548),
.B(n_549),
.C(n_552),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_614),
.B(n_489),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_594),
.B(n_478),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_576),
.B(n_496),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_618),
.B(n_478),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_559),
.B(n_506),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_607),
.A2(n_541),
.B(n_108),
.C(n_109),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_564),
.B(n_103),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_617),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_598),
.A2(n_112),
.B(n_114),
.Y(n_636)
);

INVx5_ASAP7_75t_L g637 ( 
.A(n_586),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_600),
.Y(n_638)
);

OAI21xp33_ASAP7_75t_L g639 ( 
.A1(n_610),
.A2(n_118),
.B(n_119),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_555),
.A2(n_596),
.B1(n_567),
.B2(n_626),
.Y(n_640)
);

AOI221x1_ASAP7_75t_L g641 ( 
.A1(n_610),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.C(n_133),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_573),
.A2(n_134),
.B(n_135),
.Y(n_642)
);

AO31x2_ASAP7_75t_L g643 ( 
.A1(n_616),
.A2(n_137),
.A3(n_138),
.B(n_139),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_602),
.A2(n_148),
.B(n_151),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_586),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_596),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_563),
.A2(n_165),
.B(n_167),
.Y(n_647)
);

OAI22xp33_ASAP7_75t_L g648 ( 
.A1(n_572),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_605),
.B(n_620),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_617),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_563),
.A2(n_613),
.B(n_565),
.Y(n_651)
);

A2O1A1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_571),
.A2(n_582),
.B(n_566),
.C(n_577),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_626),
.A2(n_580),
.B1(n_599),
.B2(n_593),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_569),
.B(n_557),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_626),
.A2(n_599),
.B1(n_593),
.B2(n_561),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_569),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_620),
.B(n_591),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_593),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_SL g659 ( 
.A1(n_619),
.A2(n_597),
.B(n_624),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_588),
.A2(n_601),
.B1(n_625),
.B2(n_615),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_627),
.A2(n_592),
.B(n_606),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_584),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_604),
.A2(n_609),
.B(n_623),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_585),
.A2(n_581),
.B(n_562),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_611),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_568),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_575),
.B(n_600),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_621),
.B(n_608),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_578),
.A2(n_558),
.B(n_622),
.Y(n_669)
);

AOI221x1_ASAP7_75t_L g670 ( 
.A1(n_603),
.A2(n_610),
.B1(n_555),
.B2(n_579),
.C(n_532),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_603),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_560),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_560),
.A2(n_614),
.B1(n_528),
.B2(n_555),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_587),
.B(n_474),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_594),
.B(n_528),
.Y(n_675)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_594),
.A2(n_607),
.B(n_610),
.C(n_613),
.Y(n_676)
);

OAI21xp33_ASAP7_75t_L g677 ( 
.A1(n_594),
.A2(n_610),
.B(n_607),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_617),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_594),
.B(n_528),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_620),
.B(n_575),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_614),
.B(n_441),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_594),
.A2(n_408),
.B(n_397),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_564),
.B(n_414),
.Y(n_683)
);

AOI21xp5_ASAP7_75t_L g684 ( 
.A1(n_594),
.A2(n_408),
.B(n_397),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_594),
.B(n_528),
.Y(n_685)
);

BUFx2_ASAP7_75t_L g686 ( 
.A(n_617),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_594),
.B(n_528),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_594),
.B(n_528),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_620),
.B(n_575),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_564),
.B(n_474),
.Y(n_690)
);

AOI211x1_ASAP7_75t_L g691 ( 
.A1(n_556),
.A2(n_574),
.B(n_570),
.C(n_594),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_594),
.B(n_528),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_626),
.B(n_522),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_564),
.B(n_474),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_594),
.B(n_528),
.Y(n_695)
);

BUFx2_ASAP7_75t_L g696 ( 
.A(n_617),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_561),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_617),
.Y(n_698)
);

NAND3x1_ASAP7_75t_L g699 ( 
.A(n_625),
.B(n_489),
.C(n_314),
.Y(n_699)
);

AO31x2_ASAP7_75t_L g700 ( 
.A1(n_616),
.A2(n_612),
.A3(n_565),
.B(n_519),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_594),
.B(n_528),
.Y(n_701)
);

AOI31xp67_ASAP7_75t_L g702 ( 
.A1(n_563),
.A2(n_595),
.A3(n_589),
.B(n_583),
.Y(n_702)
);

OA21x2_ASAP7_75t_L g703 ( 
.A1(n_598),
.A2(n_610),
.B(n_590),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_561),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_614),
.B(n_441),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_594),
.B(n_528),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_614),
.B(n_441),
.Y(n_707)
);

OAI22x1_ASAP7_75t_L g708 ( 
.A1(n_569),
.A2(n_374),
.B1(n_443),
.B2(n_495),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_594),
.B(n_528),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_561),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_561),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_594),
.A2(n_408),
.B(n_397),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_594),
.B(n_528),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_620),
.B(n_575),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_675),
.B(n_679),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_628),
.A2(n_629),
.B1(n_692),
.B2(n_687),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_637),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_650),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_648),
.B(n_646),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_630),
.B(n_656),
.Y(n_720)
);

OA21x2_ASAP7_75t_L g721 ( 
.A1(n_639),
.A2(n_670),
.B(n_641),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_685),
.A2(n_701),
.B1(n_688),
.B2(n_695),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_662),
.Y(n_723)
);

AOI21x1_ASAP7_75t_L g724 ( 
.A1(n_661),
.A2(n_640),
.B(n_663),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_706),
.A2(n_709),
.B1(n_713),
.B2(n_694),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_649),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_673),
.A2(n_656),
.B1(n_660),
.B2(n_691),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_654),
.B(n_690),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_676),
.A2(n_682),
.B(n_684),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_683),
.Y(n_730)
);

AOI221xp5_ASAP7_75t_L g731 ( 
.A1(n_708),
.A2(n_674),
.B1(n_677),
.B2(n_657),
.C(n_711),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_712),
.A2(n_652),
.B(n_677),
.Y(n_732)
);

OAI21xp33_ASAP7_75t_SL g733 ( 
.A1(n_673),
.A2(n_647),
.B(n_636),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_658),
.Y(n_734)
);

OA21x2_ASAP7_75t_L g735 ( 
.A1(n_639),
.A2(n_651),
.B(n_636),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_646),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_697),
.B(n_704),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_664),
.A2(n_647),
.B(n_710),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_633),
.A2(n_632),
.B(n_664),
.C(n_634),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_666),
.B(n_637),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

AOI22x1_ASAP7_75t_SL g742 ( 
.A1(n_635),
.A2(n_698),
.B1(n_678),
.B2(n_686),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_SL g743 ( 
.A(n_696),
.B(n_637),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_645),
.Y(n_744)
);

BUFx12f_ASAP7_75t_L g745 ( 
.A(n_631),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_714),
.Y(n_746)
);

AOI21xp33_ASAP7_75t_L g747 ( 
.A1(n_681),
.A2(n_707),
.B(n_705),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_689),
.B(n_714),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_631),
.B(n_668),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_638),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_645),
.B(n_631),
.Y(n_751)
);

BUFx8_ASAP7_75t_L g752 ( 
.A(n_672),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_630),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_667),
.Y(n_754)
);

INVx6_ASAP7_75t_L g755 ( 
.A(n_699),
.Y(n_755)
);

INVx6_ASAP7_75t_L g756 ( 
.A(n_671),
.Y(n_756)
);

OR2x6_ASAP7_75t_L g757 ( 
.A(n_653),
.B(n_669),
.Y(n_757)
);

INVxp33_ASAP7_75t_SL g758 ( 
.A(n_655),
.Y(n_758)
);

OAI21xp5_ASAP7_75t_L g759 ( 
.A1(n_703),
.A2(n_702),
.B(n_644),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_703),
.A2(n_693),
.B(n_700),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_643),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_700),
.B(n_643),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_650),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_635),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_665),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_659),
.A2(n_676),
.B(n_663),
.Y(n_766)
);

AOI22x1_ASAP7_75t_L g767 ( 
.A1(n_642),
.A2(n_532),
.B1(n_651),
.B2(n_682),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_682),
.A2(n_712),
.B(n_684),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_665),
.Y(n_769)
);

INVx6_ASAP7_75t_SL g770 ( 
.A(n_631),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_614),
.B1(n_656),
.B2(n_675),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_676),
.A2(n_684),
.B(n_682),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_635),
.Y(n_773)
);

CKINVDCx11_ASAP7_75t_R g774 ( 
.A(n_650),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_635),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_662),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_670),
.B(n_691),
.C(n_676),
.Y(n_777)
);

CKINVDCx8_ASAP7_75t_R g778 ( 
.A(n_635),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_635),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_662),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_637),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_670),
.B(n_691),
.C(n_676),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_665),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_675),
.B(n_679),
.Y(n_784)
);

CKINVDCx11_ASAP7_75t_R g785 ( 
.A(n_650),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_646),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_R g787 ( 
.A1(n_680),
.A2(n_569),
.B(n_348),
.Y(n_787)
);

OR2x6_ASAP7_75t_L g788 ( 
.A(n_650),
.B(n_686),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_665),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_662),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_717),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_725),
.B(n_722),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_787),
.A2(n_771),
.B1(n_716),
.B2(n_755),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_751),
.B(n_736),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_717),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_755),
.B(n_728),
.Y(n_797)
);

AO21x2_ASAP7_75t_L g798 ( 
.A1(n_759),
.A2(n_729),
.B(n_772),
.Y(n_798)
);

INVx6_ASAP7_75t_L g799 ( 
.A(n_752),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_715),
.B(n_784),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_765),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_731),
.A2(n_758),
.B1(n_737),
.B2(n_727),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_723),
.B(n_776),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_769),
.Y(n_804)
);

NOR2x1_ASAP7_75t_SL g805 ( 
.A(n_781),
.B(n_791),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_745),
.A2(n_770),
.B1(n_749),
.B2(n_763),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_780),
.B(n_790),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_783),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_718),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_770),
.A2(n_730),
.B1(n_748),
.B2(n_746),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_789),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_777),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_746),
.B(n_748),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_757),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_754),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_726),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_781),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_777),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_782),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_743),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_773),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_751),
.B(n_736),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_750),
.B(n_738),
.Y(n_823)
);

INVx2_ASAP7_75t_SL g824 ( 
.A(n_791),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_791),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_782),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_741),
.B(n_753),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_786),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_761),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_740),
.B(n_788),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_732),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_724),
.Y(n_832)
);

AO21x1_ASAP7_75t_SL g833 ( 
.A1(n_760),
.A2(n_768),
.B(n_719),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_740),
.B(n_747),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_720),
.A2(n_733),
.B1(n_767),
.B2(n_752),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_772),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_762),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_760),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_744),
.B(n_734),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_744),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_734),
.B(n_739),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_757),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_756),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_757),
.Y(n_844)
);

NOR2x1p5_ASAP7_75t_L g845 ( 
.A(n_764),
.B(n_779),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_735),
.A2(n_733),
.B1(n_779),
.B2(n_764),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_829),
.Y(n_847)
);

OR2x6_ASAP7_75t_SL g848 ( 
.A(n_846),
.B(n_774),
.Y(n_848)
);

NAND2x1p5_ASAP7_75t_L g849 ( 
.A(n_828),
.B(n_721),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_796),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_833),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_796),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_823),
.B(n_766),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_808),
.B(n_785),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_793),
.B(n_742),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_808),
.B(n_775),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_812),
.B(n_775),
.Y(n_857)
);

AND2x4_ASAP7_75t_SL g858 ( 
.A(n_795),
.B(n_778),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_809),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_812),
.B(n_818),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_832),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_794),
.A2(n_802),
.B1(n_797),
.B2(n_800),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_836),
.B(n_818),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_819),
.B(n_826),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_819),
.B(n_826),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_837),
.B(n_842),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_803),
.B(n_807),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_838),
.B(n_798),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_807),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_798),
.B(n_831),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_801),
.B(n_804),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_811),
.B(n_841),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_839),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_847),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_851),
.B(n_866),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_861),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_867),
.B(n_815),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_872),
.B(n_853),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_855),
.B(n_821),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_872),
.B(n_837),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_867),
.B(n_816),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_862),
.A2(n_799),
.B1(n_814),
.B2(n_835),
.Y(n_882)
);

BUFx2_ASAP7_75t_SL g883 ( 
.A(n_852),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_866),
.B(n_844),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_SL g885 ( 
.A1(n_858),
.A2(n_820),
.B(n_806),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_849),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_873),
.B(n_842),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_853),
.B(n_833),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_859),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_848),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_886),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_884),
.B(n_866),
.Y(n_892)
);

INVx3_ASAP7_75t_SL g893 ( 
.A(n_875),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_878),
.B(n_869),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_874),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_878),
.B(n_889),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_880),
.B(n_860),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_887),
.B(n_863),
.Y(n_898)
);

OR2x2_ASAP7_75t_L g899 ( 
.A(n_877),
.B(n_868),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_883),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_881),
.B(n_871),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_880),
.B(n_860),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_888),
.B(n_864),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_876),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_897),
.B(n_864),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_897),
.B(n_888),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_900),
.Y(n_907)
);

AND2x4_ASAP7_75t_SL g908 ( 
.A(n_892),
.B(n_875),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_904),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_896),
.B(n_870),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_896),
.B(n_870),
.Y(n_911)
);

OAI31xp33_ASAP7_75t_L g912 ( 
.A1(n_891),
.A2(n_890),
.A3(n_885),
.B(n_858),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_895),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_902),
.B(n_865),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_899),
.B(n_865),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_903),
.B(n_884),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_910),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_910),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_906),
.B(n_916),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_911),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_911),
.Y(n_921)
);

OAI33xp33_ASAP7_75t_L g922 ( 
.A1(n_915),
.A2(n_894),
.A3(n_899),
.B1(n_901),
.B2(n_855),
.B3(n_898),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_907),
.A2(n_890),
.B1(n_893),
.B2(n_848),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_913),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_909),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_907),
.B(n_879),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_913),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_924),
.Y(n_928)
);

NAND2xp33_ASAP7_75t_SL g929 ( 
.A(n_923),
.B(n_893),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_919),
.B(n_906),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_917),
.B(n_905),
.Y(n_931)
);

OAI221xp5_ASAP7_75t_L g932 ( 
.A1(n_929),
.A2(n_912),
.B1(n_926),
.B2(n_882),
.C(n_921),
.Y(n_932)
);

NOR3xp33_ASAP7_75t_L g933 ( 
.A(n_929),
.B(n_922),
.C(n_926),
.Y(n_933)
);

OAI211xp5_ASAP7_75t_SL g934 ( 
.A1(n_931),
.A2(n_912),
.B(n_920),
.C(n_918),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_934),
.B(n_928),
.Y(n_935)
);

OR2x2_ASAP7_75t_L g936 ( 
.A(n_932),
.B(n_914),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_935),
.B(n_933),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_936),
.B(n_845),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_938),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_937),
.B(n_821),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_940),
.Y(n_941)
);

NOR2x1_ASAP7_75t_L g942 ( 
.A(n_939),
.B(n_854),
.Y(n_942)
);

OAI22x1_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_942),
.B1(n_854),
.B2(n_857),
.Y(n_943)
);

XNOR2xp5_ASAP7_75t_L g944 ( 
.A(n_941),
.B(n_858),
.Y(n_944)
);

OAI211xp5_ASAP7_75t_SL g945 ( 
.A1(n_941),
.A2(n_830),
.B(n_810),
.C(n_799),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_944),
.Y(n_946)
);

XOR2x1_ASAP7_75t_L g947 ( 
.A(n_943),
.B(n_799),
.Y(n_947)
);

BUFx4f_ASAP7_75t_SL g948 ( 
.A(n_945),
.Y(n_948)
);

INVxp67_ASAP7_75t_SL g949 ( 
.A(n_944),
.Y(n_949)
);

OR3x1_ASAP7_75t_L g950 ( 
.A(n_945),
.B(n_799),
.C(n_813),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_950),
.A2(n_930),
.B1(n_857),
.B2(n_925),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_948),
.A2(n_856),
.B1(n_927),
.B2(n_925),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_949),
.B(n_946),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_947),
.A2(n_856),
.A3(n_843),
.B1(n_834),
.B2(n_817),
.C(n_825),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_946),
.Y(n_955)
);

AOI21xp33_ASAP7_75t_L g956 ( 
.A1(n_949),
.A2(n_843),
.B(n_817),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_949),
.A2(n_827),
.B(n_824),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_953),
.Y(n_958)
);

OAI21xp5_ASAP7_75t_L g959 ( 
.A1(n_955),
.A2(n_825),
.B(n_824),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_956),
.A2(n_850),
.B(n_792),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_957),
.A2(n_840),
.B1(n_908),
.B2(n_828),
.C(n_822),
.Y(n_961)
);

XNOR2xp5_ASAP7_75t_L g962 ( 
.A(n_958),
.B(n_951),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_959),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_960),
.A2(n_954),
.B(n_952),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_962),
.A2(n_961),
.B(n_805),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_962),
.A2(n_850),
.B(n_792),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_965),
.B(n_963),
.Y(n_967)
);

AOI21xp33_ASAP7_75t_SL g968 ( 
.A1(n_967),
.A2(n_966),
.B(n_964),
.Y(n_968)
);


endmodule