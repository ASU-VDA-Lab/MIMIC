module fake_jpeg_3517_n_489 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_489);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_489;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx3_ASAP7_75t_SL g43 ( 
.A(n_11),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_55),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_58),
.Y(n_149)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_61),
.Y(n_125)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_67),
.B(n_93),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_12),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_70),
.B(n_78),
.Y(n_132)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_73),
.Y(n_156)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_11),
.Y(n_78)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_10),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_96),
.Y(n_105)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_15),
.Y(n_81)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_90),
.Y(n_100)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_97),
.Y(n_126)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_43),
.B(n_45),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_10),
.Y(n_96)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_32),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_17),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_83),
.B1(n_94),
.B2(n_56),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_102),
.A2(n_107),
.B1(n_127),
.B2(n_142),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_65),
.B1(n_90),
.B2(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_108),
.A2(n_119),
.B1(n_143),
.B2(n_87),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_66),
.A2(n_38),
.B1(n_35),
.B2(n_17),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_42),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_141),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_126),
.B(n_43),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_76),
.B1(n_98),
.B2(n_57),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_20),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_72),
.A2(n_17),
.B1(n_24),
.B2(n_40),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_86),
.A2(n_38),
.B1(n_17),
.B2(n_24),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_79),
.A2(n_24),
.B1(n_40),
.B2(n_29),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_142),
.B1(n_39),
.B2(n_24),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_120),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_157),
.B(n_164),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_108),
.A2(n_29),
.B1(n_45),
.B2(n_30),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_159),
.A2(n_185),
.B1(n_198),
.B2(n_157),
.Y(n_206)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_160),
.Y(n_214)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_129),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_47),
.B1(n_92),
.B2(n_68),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

BUFx2_ASAP7_75t_SL g168 ( 
.A(n_138),
.Y(n_168)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_182),
.B1(n_151),
.B2(n_149),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_170),
.B(n_184),
.Y(n_219)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_171),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_93),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_174),
.B(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_110),
.B(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_187),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_181),
.B(n_189),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_53),
.B1(n_77),
.B2(n_38),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_183),
.A2(n_201),
.B(n_43),
.Y(n_225)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g186 ( 
.A(n_114),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_99),
.B(n_39),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_69),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_103),
.B(n_27),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_191),
.Y(n_222)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_130),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

AO22x1_ASAP7_75t_SL g193 ( 
.A1(n_113),
.A2(n_68),
.B1(n_43),
.B2(n_60),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_116),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_196),
.B(n_199),
.Y(n_213)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_100),
.A2(n_31),
.B1(n_22),
.B2(n_18),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_128),
.B(n_43),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_101),
.B(n_43),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_150),
.C(n_134),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_203),
.B(n_221),
.C(n_193),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_161),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_208),
.A2(n_220),
.B1(n_224),
.B2(n_226),
.Y(n_257)
);

MAJx3_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_43),
.C(n_138),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_209),
.A2(n_235),
.B(n_232),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_111),
.B1(n_139),
.B2(n_137),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_104),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_183),
.A2(n_111),
.B1(n_139),
.B2(n_137),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_225),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_112),
.B1(n_151),
.B2(n_149),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_158),
.A2(n_140),
.B1(n_121),
.B2(n_145),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_186),
.B1(n_166),
.B2(n_164),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_207),
.B(n_189),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_250),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_158),
.B1(n_169),
.B2(n_193),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_239),
.A2(n_244),
.B1(n_262),
.B2(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_242),
.A2(n_218),
.B1(n_186),
.B2(n_216),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_202),
.A2(n_190),
.B(n_146),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_245),
.A2(n_255),
.B(n_265),
.Y(n_280)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_246),
.Y(n_292)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_210),
.Y(n_247)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_247),
.Y(n_276)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_175),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_256),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_252),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_258),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_209),
.B(n_219),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_221),
.B(n_184),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_260),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_199),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_261),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_219),
.A2(n_112),
.B1(n_117),
.B2(n_109),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_196),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_249),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_219),
.A2(n_171),
.B(n_166),
.Y(n_264)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_203),
.C(n_209),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_268),
.C(n_271),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_265),
.C(n_258),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_259),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_209),
.C(n_232),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_233),
.C(n_231),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_181),
.C(n_191),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_281),
.B1(n_289),
.B2(n_290),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_279),
.A2(n_284),
.B(n_222),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_220),
.B1(n_206),
.B2(n_226),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_283),
.A2(n_293),
.B1(n_284),
.B2(n_289),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_222),
.B(n_214),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_239),
.A2(n_216),
.B1(n_214),
.B2(n_218),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_217),
.B1(n_176),
.B2(n_173),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_257),
.A2(n_217),
.B1(n_167),
.B2(n_117),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_229),
.B1(n_233),
.B2(n_231),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_248),
.B1(n_247),
.B2(n_240),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_263),
.B1(n_244),
.B2(n_245),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_312),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_297),
.B(n_304),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_298),
.B(n_273),
.Y(n_339)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_237),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_303),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_251),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_302),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_254),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_269),
.B(n_260),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_256),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_307),
.A2(n_310),
.B1(n_320),
.B2(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_270),
.B(n_264),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_322),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_281),
.A2(n_245),
.B1(n_264),
.B2(n_242),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_262),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_314),
.C(n_315),
.Y(n_336)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_286),
.B(n_234),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_313),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_241),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_222),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_317),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_180),
.C(n_192),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_280),
.A2(n_215),
.B(n_229),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_321),
.B(n_316),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_282),
.A2(n_250),
.B1(n_261),
.B2(n_217),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_279),
.B(n_278),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_211),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_282),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_277),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_294),
.A2(n_261),
.B1(n_250),
.B2(n_246),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_320),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_344),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_347),
.B(n_326),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_331),
.Y(n_358)
);

XOR2x2_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_314),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_334),
.A2(n_347),
.B(n_315),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_317),
.A2(n_277),
.B1(n_284),
.B2(n_273),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_335),
.A2(n_292),
.B1(n_228),
.B2(n_204),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_295),
.A2(n_284),
.B1(n_283),
.B2(n_293),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_337),
.A2(n_353),
.B1(n_306),
.B2(n_312),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_350),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_301),
.B(n_274),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_341),
.B(n_310),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_287),
.Y(n_342)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_342),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_324),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_287),
.B(n_276),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_319),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_349),
.B(n_352),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_302),
.B(n_276),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_308),
.C(n_309),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_299),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_305),
.Y(n_353)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_355),
.A2(n_344),
.B1(n_327),
.B2(n_333),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_308),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_365),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_359),
.A2(n_326),
.B(n_332),
.Y(n_383)
);

AOI21xp33_ASAP7_75t_L g398 ( 
.A1(n_360),
.A2(n_325),
.B(n_338),
.Y(n_398)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_354),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_371),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_364),
.B(n_373),
.C(n_351),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_311),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_322),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_374),
.Y(n_390)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_377),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_291),
.B(n_292),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_291),
.C(n_228),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_211),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_375),
.A2(n_381),
.B1(n_352),
.B2(n_346),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_336),
.B(n_215),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_348),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_379),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_234),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_163),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_380),
.B(n_346),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_343),
.A2(n_292),
.B1(n_204),
.B2(n_160),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_362),
.Y(n_382)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_395),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_376),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_388),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_331),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_387),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g388 ( 
.A(n_370),
.B(n_359),
.CI(n_335),
.CON(n_388),
.SN(n_388)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_0),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_332),
.B(n_349),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_399),
.B1(n_345),
.B2(n_379),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_361),
.B(n_353),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_400),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_138),
.Y(n_421)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_194),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_371),
.A2(n_337),
.B1(n_332),
.B2(n_333),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_402),
.A2(n_403),
.B1(n_404),
.B2(n_162),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_374),
.A2(n_340),
.B1(n_329),
.B2(n_345),
.Y(n_404)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_364),
.C(n_356),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_407),
.B(n_415),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_392),
.A2(n_373),
.B1(n_380),
.B2(n_366),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_408),
.A2(n_421),
.B1(n_9),
.B2(n_8),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_409),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_377),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_410),
.B(n_412),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_366),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_365),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g429 ( 
.A(n_413),
.B(n_384),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_378),
.C(n_367),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_385),
.B(n_178),
.C(n_197),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_416),
.B(n_417),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_394),
.B(n_133),
.C(n_145),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_177),
.C(n_140),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_422),
.C(n_390),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_419),
.A2(n_399),
.B1(n_388),
.B2(n_395),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_109),
.C(n_1),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_423),
.B(n_9),
.Y(n_435)
);

OAI321xp33_ASAP7_75t_L g425 ( 
.A1(n_405),
.A2(n_387),
.A3(n_393),
.B1(n_391),
.B2(n_383),
.C(n_402),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_440),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_433),
.Y(n_450)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_428),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_429),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_411),
.A2(n_388),
.B1(n_384),
.B2(n_9),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_438),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_407),
.B(n_0),
.C(n_1),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_434),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_1),
.C(n_2),
.Y(n_434)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_435),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_9),
.Y(n_436)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_8),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_423),
.B(n_1),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_7),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_442),
.B(n_1),
.Y(n_451)
);

BUFx24_ASAP7_75t_SL g446 ( 
.A(n_437),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_446),
.B(n_438),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_414),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_430),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_414),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_451),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_428),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_452),
.B(n_453),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_441),
.B(n_432),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_431),
.B(n_421),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_454),
.B(n_434),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_444),
.A2(n_432),
.B(n_439),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_459),
.A2(n_464),
.B(n_466),
.Y(n_469)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_460),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_465),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_445),
.A2(n_416),
.B(n_417),
.Y(n_463)
);

AO21x1_ASAP7_75t_L g473 ( 
.A1(n_463),
.A2(n_467),
.B(n_457),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_418),
.B(n_436),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_SL g466 ( 
.A1(n_443),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_452),
.A2(n_2),
.B(n_3),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_457),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_468),
.A2(n_448),
.B(n_3),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_455),
.Y(n_471)
);

AO21x1_ASAP7_75t_L g478 ( 
.A1(n_471),
.A2(n_473),
.B(n_476),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_450),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_474),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_466),
.B(n_456),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_2),
.C(n_3),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_6),
.C(n_7),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_4),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_480),
.B(n_481),
.C(n_5),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_4),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_482),
.B(n_483),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_469),
.C(n_6),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_478),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_477),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_487),
.B(n_486),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_488),
.A2(n_6),
.B(n_487),
.Y(n_489)
);


endmodule