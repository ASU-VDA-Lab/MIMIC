module fake_ariane_350_n_82 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_82);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_82;

wire n_56;
wire n_60;
wire n_64;
wire n_38;
wire n_47;
wire n_75;
wire n_67;
wire n_34;
wire n_69;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_20;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_36;
wire n_72;
wire n_44;
wire n_30;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_23;
wire n_61;
wire n_22;
wire n_43;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_4),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_11),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_6),
.B(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_19),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_20),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_26),
.Y(n_41)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_24),
.B(n_22),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_39),
.B(n_32),
.C(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_32),
.B1(n_30),
.B2(n_26),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_26),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

OA21x2_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_25),
.B(n_21),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_21),
.B(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_46),
.Y(n_51)
);

AOI21x1_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_31),
.B(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_45),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_26),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_50),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_23),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_23),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_23),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_50),
.B(n_53),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_48),
.B(n_53),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_59),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

XOR2x2_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_48),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_48),
.B(n_59),
.Y(n_69)
);

OAI211xp5_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_57),
.B1(n_47),
.B2(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_57),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_58),
.B(n_49),
.Y(n_73)
);

AND4x1_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_23),
.C(n_60),
.D(n_64),
.Y(n_74)
);

NOR4xp25_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_60),
.C(n_49),
.D(n_52),
.Y(n_75)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_31),
.C(n_52),
.Y(n_76)
);

NAND4xp75_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_71),
.C(n_72),
.D(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

AOI22x1_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_31),
.B1(n_75),
.B2(n_69),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_72),
.B1(n_52),
.B2(n_31),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_77),
.B(n_31),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_79),
.Y(n_82)
);


endmodule