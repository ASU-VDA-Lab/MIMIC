module fake_jpeg_25900_n_218 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_218);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_28),
.A2(n_30),
.B1(n_17),
.B2(n_21),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_18),
.B(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_19),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_22),
.B1(n_11),
.B2(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_22),
.B1(n_11),
.B2(n_12),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_22),
.B1(n_11),
.B2(n_17),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_30),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_49),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_25),
.B(n_21),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_62),
.B(n_16),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_41),
.Y(n_63)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_28),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_65),
.B(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_31),
.C(n_41),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_71),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_31),
.C(n_41),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_31),
.C(n_41),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_78),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_38),
.C(n_37),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_43),
.B(n_1),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_83),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_33),
.B1(n_41),
.B2(n_29),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_59),
.B1(n_55),
.B2(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_43),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_52),
.B1(n_51),
.B2(n_62),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_94),
.B1(n_96),
.B2(n_105),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.B(n_29),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_89),
.B(n_103),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_33),
.B1(n_58),
.B2(n_57),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_15),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_91),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_99),
.B1(n_74),
.B2(n_77),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_33),
.B1(n_60),
.B2(n_48),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_66),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_32),
.B1(n_43),
.B2(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_19),
.B1(n_15),
.B2(n_23),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_108),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_107),
.B(n_65),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_20),
.B1(n_13),
.B2(n_32),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_76),
.B(n_13),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_111),
.A2(n_0),
.B(n_1),
.Y(n_153)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

OA21x2_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_76),
.B(n_63),
.Y(n_115)
);

NOR2xp67_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_86),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_121),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_89),
.B1(n_105),
.B2(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_68),
.C(n_82),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_129),
.C(n_94),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_68),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_128),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_72),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_66),
.C(n_64),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_72),
.Y(n_130)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_137),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_147),
.B1(n_149),
.B2(n_116),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_127),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_107),
.B(n_89),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_138),
.Y(n_161)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_98),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_85),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_153),
.C(n_125),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_112),
.A2(n_99),
.B1(n_95),
.B2(n_72),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_123),
.B(n_118),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_132),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_77),
.B(n_66),
.C(n_43),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_154),
.B1(n_120),
.B2(n_122),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_43),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_43),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_133),
.C(n_154),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_117),
.B1(n_119),
.B2(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_162),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_110),
.C(n_119),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_163),
.C(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_114),
.B1(n_118),
.B2(n_109),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_113),
.C(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_144),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_130),
.B1(n_113),
.B2(n_77),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_137),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_145),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_144),
.Y(n_173)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_159),
.B(n_142),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_177),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_133),
.C(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_159),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_139),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_176),
.A2(n_165),
.B1(n_161),
.B2(n_168),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_185),
.B1(n_163),
.B2(n_152),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_156),
.B1(n_168),
.B2(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_170),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_178),
.A2(n_166),
.B(n_153),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_151),
.B(n_160),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_199),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_191),
.C(n_9),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_182),
.C(n_190),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_194),
.B(n_198),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_195),
.A2(n_191),
.B(n_188),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_197),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_132),
.B(n_10),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_9),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_203),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_2),
.C(n_3),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_0),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_206),
.B(n_208),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_209),
.B(n_3),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_205),
.B(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_3),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_210),
.A2(n_204),
.B(n_4),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_211),
.A2(n_4),
.B(n_5),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_213),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.C(n_8),
.Y(n_216)
);

OAI221xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_8),
.Y(n_218)
);


endmodule