module fake_jpeg_5716_n_114 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_4),
.B(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_24),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_14),
.A2(n_0),
.B1(n_9),
.B2(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_18),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_5),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_11),
.Y(n_30)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_12),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_18),
.B(n_10),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_7),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_21),
.B1(n_24),
.B2(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_42),
.B(n_49),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_14),
.B1(n_28),
.B2(n_13),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_46),
.B1(n_49),
.B2(n_45),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_33),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_25),
.C(n_24),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_25),
.C(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_50),
.Y(n_53)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_61),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_34),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_47),
.B(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_50),
.C(n_46),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_31),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_45),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g74 ( 
.A1(n_62),
.A2(n_72),
.B(n_61),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_31),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_46),
.C(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_10),
.Y(n_76)
);

NOR4xp25_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_58),
.C(n_54),
.D(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_71),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_36),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_25),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_66),
.C(n_21),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_51),
.B1(n_53),
.B2(n_58),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_39),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_6),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_6),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_38),
.B1(n_22),
.B2(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_39),
.C(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_38),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_90),
.B(n_91),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_39),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_90),
.A2(n_77),
.B1(n_19),
.B2(n_10),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_94),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_89),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_98),
.A2(n_20),
.B(n_19),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_8),
.B(n_1),
.C(n_2),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_96),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_3),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_98),
.B(n_92),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_102),
.C(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_0),
.A3(n_9),
.B1(n_20),
.B2(n_93),
.C1(n_99),
.C2(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_109),
.C(n_9),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_0),
.B(n_111),
.Y(n_114)
);


endmodule