module real_aes_819_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_0), .B(n_237), .Y(n_260) );
OAI22xp5_ASAP7_75t_SL g195 ( .A1(n_1), .A2(n_46), .B1(n_196), .B2(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_1), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_2), .A2(n_232), .B(n_296), .Y(n_295) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_3), .A2(n_55), .B1(n_94), .B2(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_4), .B(n_248), .Y(n_276) );
INVx1_ASAP7_75t_L g215 ( .A(n_5), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_6), .B(n_248), .Y(n_305) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_7), .A2(n_21), .B1(n_94), .B2(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g348 ( .A(n_8), .B(n_246), .Y(n_348) );
INVx2_ASAP7_75t_L g229 ( .A(n_9), .Y(n_229) );
AOI221x1_ASAP7_75t_L g231 ( .A1(n_10), .A2(n_18), .B1(n_232), .B2(n_237), .C(n_244), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g344 ( .A(n_11), .B(n_237), .Y(n_344) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_12), .A2(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_13), .B(n_227), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_14), .A2(n_61), .B1(n_178), .B2(n_181), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_15), .B(n_248), .Y(n_330) );
AO21x1_ASAP7_75t_L g270 ( .A1(n_16), .A2(n_237), .B(n_271), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_17), .A2(n_40), .B1(n_169), .B2(n_172), .Y(n_168) );
NAND2x1_ASAP7_75t_L g258 ( .A(n_19), .B(n_248), .Y(n_258) );
NAND2x1_ASAP7_75t_L g304 ( .A(n_20), .B(n_246), .Y(n_304) );
INVx1_ASAP7_75t_L g550 ( .A(n_20), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g207 ( .A1(n_21), .A2(n_55), .B1(n_60), .B2(n_208), .C(n_210), .Y(n_207) );
OR2x2_ASAP7_75t_L g230 ( .A(n_22), .B(n_68), .Y(n_230) );
OA21x2_ASAP7_75t_L g264 ( .A1(n_22), .A2(n_68), .B(n_229), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_23), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_24), .B(n_246), .Y(n_298) );
INVx3_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_26), .B(n_248), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_27), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_28), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_29), .B(n_246), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g80 ( .A1(n_30), .A2(n_81), .B1(n_185), .B2(n_186), .Y(n_80) );
INVx1_ASAP7_75t_L g186 ( .A(n_30), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_31), .A2(n_232), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g95 ( .A(n_32), .Y(n_95) );
INVx1_ASAP7_75t_L g217 ( .A(n_33), .Y(n_217) );
AND2x2_ASAP7_75t_L g233 ( .A(n_33), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g243 ( .A(n_33), .B(n_215), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_34), .B(n_237), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_35), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_36), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_37), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_38), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_39), .B(n_246), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_41), .A2(n_232), .B(n_303), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_41), .A2(n_81), .B1(n_185), .B2(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_41), .Y(n_535) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_42), .A2(n_60), .B1(n_94), .B2(n_98), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_43), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_44), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_45), .B(n_246), .Y(n_259) );
INVx1_ASAP7_75t_L g197 ( .A(n_46), .Y(n_197) );
INVx1_ASAP7_75t_L g236 ( .A(n_47), .Y(n_236) );
INVx1_ASAP7_75t_L g240 ( .A(n_47), .Y(n_240) );
INVx1_ASAP7_75t_L g96 ( .A(n_48), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_49), .B(n_248), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_50), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_189) );
INVx1_ASAP7_75t_L g191 ( .A(n_50), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_50), .A2(n_232), .B(n_257), .Y(n_256) );
AO21x1_ASAP7_75t_L g273 ( .A1(n_51), .A2(n_232), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_52), .B(n_237), .Y(n_294) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_53), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_54), .B(n_237), .Y(n_306) );
INVxp33_ASAP7_75t_L g212 ( .A(n_55), .Y(n_212) );
INVx1_ASAP7_75t_L g201 ( .A(n_56), .Y(n_201) );
AND2x2_ASAP7_75t_L g287 ( .A(n_57), .B(n_228), .Y(n_287) );
INVx1_ASAP7_75t_L g234 ( .A(n_58), .Y(n_234) );
INVx1_ASAP7_75t_L g242 ( .A(n_58), .Y(n_242) );
AND2x2_ASAP7_75t_L g308 ( .A(n_59), .B(n_262), .Y(n_308) );
INVxp67_ASAP7_75t_L g211 ( .A(n_60), .Y(n_211) );
AND2x2_ASAP7_75t_L g292 ( .A(n_62), .B(n_262), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_63), .B(n_237), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_64), .Y(n_152) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_65), .A2(n_81), .B1(n_185), .B2(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_65), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_66), .B(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g271 ( .A(n_67), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g265 ( .A(n_69), .B(n_262), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_70), .B(n_246), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_71), .B(n_248), .Y(n_285) );
INVx1_ASAP7_75t_L g190 ( .A(n_72), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_72), .A2(n_232), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_73), .B(n_246), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_74), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_74), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_75), .B(n_248), .Y(n_297) );
BUFx2_ASAP7_75t_SL g209 ( .A(n_76), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_77), .A2(n_232), .B(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_204), .B1(n_218), .B2(n_526), .C(n_533), .Y(n_78) );
XOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_187), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_81), .Y(n_185) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND4xp75_ASAP7_75t_L g82 ( .A(n_83), .B(n_121), .C(n_147), .D(n_167), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
OAI221xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_86), .B1(n_106), .B2(n_113), .C(n_114), .Y(n_84) );
INVx3_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
BUFx6f_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx3_ASAP7_75t_SL g88 ( .A(n_89), .Y(n_88) );
INVx6_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_99), .Y(n_90) );
AND2x4_ASAP7_75t_L g174 ( .A(n_91), .B(n_175), .Y(n_174) );
AND2x4_ASAP7_75t_L g183 ( .A(n_91), .B(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g91 ( .A(n_92), .B(n_97), .Y(n_91) );
AND2x2_ASAP7_75t_L g111 ( .A(n_92), .B(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_92), .Y(n_120) );
INVx2_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
OAI22x1_ASAP7_75t_L g92 ( .A1(n_93), .A2(n_94), .B1(n_95), .B2(n_96), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g98 ( .A(n_94), .Y(n_98) );
INVx2_ASAP7_75t_L g102 ( .A(n_94), .Y(n_102) );
INVx1_ASAP7_75t_L g105 ( .A(n_94), .Y(n_105) );
INVx2_ASAP7_75t_L g112 ( .A(n_97), .Y(n_112) );
AND2x2_ASAP7_75t_L g130 ( .A(n_97), .B(n_131), .Y(n_130) );
BUFx2_ASAP7_75t_L g134 ( .A(n_97), .Y(n_134) );
AND2x2_ASAP7_75t_L g142 ( .A(n_99), .B(n_130), .Y(n_142) );
AND2x4_ASAP7_75t_L g151 ( .A(n_99), .B(n_111), .Y(n_151) );
AND2x4_ASAP7_75t_L g162 ( .A(n_99), .B(n_146), .Y(n_162) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_103), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
AND2x4_ASAP7_75t_L g110 ( .A(n_101), .B(n_103), .Y(n_110) );
AND2x2_ASAP7_75t_L g119 ( .A(n_101), .B(n_104), .Y(n_119) );
INVx1_ASAP7_75t_L g129 ( .A(n_101), .Y(n_129) );
INVxp67_ASAP7_75t_L g184 ( .A(n_103), .Y(n_184) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g128 ( .A(n_104), .B(n_129), .Y(n_128) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x4_ASAP7_75t_L g166 ( .A(n_110), .B(n_146), .Y(n_166) );
AND2x4_ASAP7_75t_L g180 ( .A(n_110), .B(n_130), .Y(n_180) );
AND2x2_ASAP7_75t_L g171 ( .A(n_111), .B(n_128), .Y(n_171) );
AND2x4_ASAP7_75t_L g146 ( .A(n_112), .B(n_131), .Y(n_146) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx12f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x4_ASAP7_75t_L g133 ( .A(n_119), .B(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g155 ( .A(n_119), .B(n_146), .Y(n_155) );
NOR2x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_136), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_132), .B2(n_135), .Y(n_122) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_130), .Y(n_127) );
AND2x4_ASAP7_75t_L g145 ( .A(n_128), .B(n_146), .Y(n_145) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
INVx5_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_138), .B1(n_143), .B2(n_144), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx8_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2x1_ASAP7_75t_L g147 ( .A(n_148), .B(n_156), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B1(n_152), .B2(n_153), .Y(n_148) );
INVx6_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx2_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B1(n_163), .B2(n_164), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
INVx8_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_177), .Y(n_167) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx6_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B1(n_193), .B2(n_203), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g192 ( .A(n_190), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_193), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B1(n_198), .B2(n_199), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_195), .Y(n_194) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_206), .Y(n_205) );
AND3x1_ASAP7_75t_SL g206 ( .A(n_207), .B(n_213), .C(n_216), .Y(n_206) );
INVxp67_ASAP7_75t_L g539 ( .A(n_207), .Y(n_539) );
CKINVDCx8_ASAP7_75t_R g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_213), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g546 ( .A1(n_213), .A2(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g530 ( .A(n_214), .B(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_SL g544 ( .A(n_214), .B(n_216), .Y(n_544) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g235 ( .A(n_215), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_216), .B(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND4xp75_ASAP7_75t_L g220 ( .A(n_221), .B(n_436), .C(n_476), .D(n_505), .Y(n_220) );
NOR2x1_ASAP7_75t_L g221 ( .A(n_222), .B(n_398), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_355), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_288), .B(n_309), .Y(n_223) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_225), .B(n_251), .Y(n_224) );
AND2x4_ASAP7_75t_L g354 ( .A(n_225), .B(n_314), .Y(n_354) );
INVx1_ASAP7_75t_SL g407 ( .A(n_225), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_225), .A2(n_443), .B(n_446), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_SL g446 ( .A1(n_225), .A2(n_447), .B(n_448), .C(n_449), .Y(n_446) );
NAND2x1_ASAP7_75t_L g487 ( .A(n_225), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_225), .B(n_448), .Y(n_509) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g312 ( .A(n_226), .Y(n_312) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_226), .Y(n_386) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_231), .B(n_250), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_227), .A2(n_294), .B(n_295), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_227), .Y(n_307) );
OA21x2_ASAP7_75t_L g396 ( .A1(n_227), .A2(n_231), .B(n_250), .Y(n_396) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_SL g228 ( .A(n_229), .B(n_230), .Y(n_228) );
AND2x4_ASAP7_75t_L g272 ( .A(n_229), .B(n_230), .Y(n_272) );
AND2x6_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
BUFx3_ASAP7_75t_L g532 ( .A(n_233), .Y(n_532) );
AND2x6_ASAP7_75t_L g246 ( .A(n_234), .B(n_239), .Y(n_246) );
AND2x4_ASAP7_75t_L g248 ( .A(n_236), .B(n_241), .Y(n_248) );
INVx2_ASAP7_75t_L g531 ( .A(n_236), .Y(n_531) );
AND2x4_ASAP7_75t_L g237 ( .A(n_238), .B(n_243), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_241), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx5_ASAP7_75t_L g249 ( .A(n_243), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_247), .B(n_249), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_249), .A2(n_258), .B(n_259), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_249), .A2(n_275), .B(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_249), .A2(n_284), .B(n_285), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_249), .A2(n_297), .B(n_298), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_249), .A2(n_304), .B(n_305), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_249), .A2(n_330), .B(n_331), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_249), .A2(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_266), .Y(n_251) );
AND2x2_ASAP7_75t_L g378 ( .A(n_252), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g459 ( .A(n_252), .B(n_314), .Y(n_459) );
INVx1_ASAP7_75t_L g519 ( .A(n_252), .Y(n_519) );
BUFx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g363 ( .A(n_253), .B(n_279), .Y(n_363) );
AND2x2_ASAP7_75t_L g488 ( .A(n_253), .B(n_280), .Y(n_488) );
AND2x2_ASAP7_75t_L g493 ( .A(n_253), .B(n_453), .Y(n_493) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVxp67_ASAP7_75t_L g369 ( .A(n_254), .Y(n_369) );
BUFx3_ASAP7_75t_L g402 ( .A(n_254), .Y(n_402) );
AND2x2_ASAP7_75t_L g448 ( .A(n_254), .B(n_280), .Y(n_448) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_261), .B(n_265), .Y(n_254) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_255), .A2(n_261), .B(n_265), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_260), .Y(n_255) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_261), .A2(n_281), .B(n_287), .Y(n_280) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_261), .A2(n_281), .B(n_287), .Y(n_315) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
AND2x2_ASAP7_75t_L g433 ( .A(n_266), .B(n_311), .Y(n_433) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_279), .Y(n_266) );
AND2x4_ASAP7_75t_L g314 ( .A(n_267), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g425 ( .A(n_267), .B(n_409), .Y(n_425) );
AND2x2_ASAP7_75t_SL g468 ( .A(n_267), .B(n_396), .Y(n_468) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx2_ASAP7_75t_L g404 ( .A(n_268), .Y(n_404) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g365 ( .A(n_269), .Y(n_365) );
OAI21x1_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_273), .B(n_277), .Y(n_269) );
INVx1_ASAP7_75t_L g278 ( .A(n_271), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_272), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g326 ( .A(n_272), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_272), .A2(n_344), .B(n_345), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_279), .B(n_365), .Y(n_368) );
AND2x2_ASAP7_75t_L g453 ( .A(n_279), .B(n_396), .Y(n_453) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g450 ( .A(n_280), .B(n_312), .Y(n_450) );
AND2x2_ASAP7_75t_L g470 ( .A(n_280), .B(n_396), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_286), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_288), .B(n_359), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_288), .A2(n_482), .B1(n_483), .B2(n_484), .C(n_486), .Y(n_481) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI332xp33_ASAP7_75t_L g515 ( .A1(n_289), .A2(n_375), .A3(n_382), .B1(n_441), .B2(n_516), .B3(n_517), .C1(n_518), .C2(n_520), .Y(n_515) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_290), .B(n_299), .Y(n_289) );
AND2x2_ASAP7_75t_L g320 ( .A(n_290), .B(n_300), .Y(n_320) );
AND2x2_ASAP7_75t_L g337 ( .A(n_290), .B(n_338), .Y(n_337) );
INVx4_ASAP7_75t_L g350 ( .A(n_290), .Y(n_350) );
AND2x2_ASAP7_75t_SL g410 ( .A(n_290), .B(n_351), .Y(n_410) );
INVx5_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2x1_ASAP7_75t_SL g372 ( .A(n_291), .B(n_338), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_291), .B(n_299), .Y(n_376) );
AND2x2_ASAP7_75t_L g383 ( .A(n_291), .B(n_300), .Y(n_383) );
BUFx2_ASAP7_75t_L g418 ( .A(n_291), .Y(n_418) );
AND2x2_ASAP7_75t_L g473 ( .A(n_291), .B(n_341), .Y(n_473) );
OR2x6_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
OR2x2_ASAP7_75t_L g340 ( .A(n_299), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g351 ( .A(n_299), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g391 ( .A(n_299), .Y(n_391) );
AND2x2_ASAP7_75t_L g461 ( .A(n_299), .B(n_360), .Y(n_461) );
AND2x2_ASAP7_75t_L g474 ( .A(n_299), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_299), .B(n_475), .Y(n_492) );
INVx4_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_307), .B(n_308), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_306), .Y(n_301) );
OAI32xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_316), .A3(n_321), .B1(n_335), .B2(n_353), .Y(n_309) );
INVx2_ASAP7_75t_L g419 ( .A(n_310), .Y(n_419) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
INVx1_ASAP7_75t_L g430 ( .A(n_311), .Y(n_430) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g364 ( .A(n_312), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g497 ( .A(n_312), .B(n_402), .Y(n_497) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g409 ( .A(n_315), .Y(n_409) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx2_ASAP7_75t_L g397 ( .A(n_318), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_318), .B(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_SL g408 ( .A(n_319), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g485 ( .A(n_319), .Y(n_485) );
AND2x2_ASAP7_75t_L g503 ( .A(n_319), .B(n_365), .Y(n_503) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp67_ASAP7_75t_SL g447 ( .A(n_322), .B(n_376), .Y(n_447) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_323), .B(n_358), .Y(n_445) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g521 ( .A(n_324), .B(n_391), .Y(n_521) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
INVx2_ASAP7_75t_L g393 ( .A(n_325), .Y(n_393) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B(n_333), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_326), .B(n_334), .Y(n_333) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_326), .A2(n_327), .B(n_333), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_332), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_349), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_336), .B(n_395), .Y(n_480) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AND3x2_ASAP7_75t_L g435 ( .A(n_337), .B(n_382), .C(n_391), .Y(n_435) );
AND2x2_ASAP7_75t_L g359 ( .A(n_338), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_338), .B(n_341), .Y(n_416) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g370 ( .A(n_340), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
INVx1_ASAP7_75t_L g375 ( .A(n_341), .Y(n_375) );
BUFx3_ASAP7_75t_L g382 ( .A(n_341), .Y(n_382) );
AND2x2_ASAP7_75t_L g392 ( .A(n_341), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x4_ASAP7_75t_L g401 ( .A(n_350), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_350), .B(n_360), .Y(n_444) );
AND2x2_ASAP7_75t_L g400 ( .A(n_351), .B(n_375), .Y(n_400) );
INVx2_ASAP7_75t_L g427 ( .A(n_351), .Y(n_427) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .B(n_366), .C(n_387), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_356), .A2(n_483), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_359), .B(n_418), .Y(n_417) );
AOI211xp5_ASAP7_75t_SL g437 ( .A1(n_359), .A2(n_438), .B(n_442), .C(n_451), .Y(n_437) );
AND2x2_ASAP7_75t_L g423 ( .A(n_360), .B(n_383), .Y(n_423) );
OR2x2_ASAP7_75t_L g426 ( .A(n_360), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_363), .B(n_468), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_364), .B(n_409), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_364), .A2(n_390), .B1(n_470), .B2(n_473), .C(n_479), .Y(n_478) );
AND2x4_ASAP7_75t_L g395 ( .A(n_365), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g441 ( .A(n_365), .B(n_396), .Y(n_441) );
OAI221xp5_ASAP7_75t_SL g366 ( .A1(n_367), .A2(n_370), .B1(n_373), .B2(n_377), .C(n_380), .Y(n_366) );
AND2x2_ASAP7_75t_L g512 ( .A(n_367), .B(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g379 ( .A(n_368), .Y(n_379) );
INVx1_ASAP7_75t_L g465 ( .A(n_369), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_370), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g384 ( .A(n_372), .B(n_375), .Y(n_384) );
AND2x2_ASAP7_75t_L g460 ( .A(n_372), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g385 ( .A(n_379), .B(n_386), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_384), .B(n_385), .Y(n_380) );
INVx1_ASAP7_75t_L g504 ( .A(n_381), .Y(n_504) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g483 ( .A(n_382), .B(n_410), .Y(n_483) );
AND2x2_ASAP7_75t_SL g456 ( .A(n_383), .B(n_392), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_394), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g424 ( .A1(n_388), .A2(n_422), .B1(n_425), .B2(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g494 ( .A(n_388), .Y(n_494) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_L g414 ( .A(n_391), .Y(n_414) );
INVx1_ASAP7_75t_L g475 ( .A(n_393), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_395), .B(n_397), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_395), .B(n_465), .Y(n_516) );
AND2x2_ASAP7_75t_L g484 ( .A(n_396), .B(n_485), .Y(n_484) );
OAI211xp5_ASAP7_75t_L g477 ( .A1(n_397), .A2(n_478), .B(n_481), .C(n_489), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_420), .Y(n_398) );
AOI322xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .A3(n_403), .B1(n_405), .B2(n_410), .C1(n_411), .C2(n_419), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_401), .Y(n_517) );
AND2x2_ASAP7_75t_L g467 ( .A(n_402), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g501 ( .A(n_402), .Y(n_501) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_SL g452 ( .A(n_404), .B(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_404), .B(n_450), .Y(n_458) );
AND2x2_ASAP7_75t_L g482 ( .A(n_404), .B(n_448), .Y(n_482) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g454 ( .A(n_408), .Y(n_454) );
NAND2xp33_ASAP7_75t_SL g411 ( .A(n_412), .B(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_SL g457 ( .A1(n_413), .A2(n_458), .B1(n_459), .B2(n_460), .C(n_462), .Y(n_457) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g524 ( .A(n_416), .Y(n_524) );
AOI211xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B(n_424), .C(n_428), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g499 ( .A(n_423), .Y(n_499) );
INVx1_ASAP7_75t_L g431 ( .A(n_425), .Y(n_431) );
OR2x2_ASAP7_75t_L g518 ( .A(n_425), .B(n_519), .Y(n_518) );
INVx2_ASAP7_75t_SL g514 ( .A(n_426), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_432), .B(n_434), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_430), .B(n_448), .Y(n_525) );
INVx1_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_457), .Y(n_436) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_440), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
OR2x2_ASAP7_75t_L g491 ( .A(n_444), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI21xp33_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_454), .B(n_455), .Y(n_451) );
INVx2_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
AOI31xp33_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .A3(n_469), .B(n_471), .Y(n_462) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_468), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B1(n_494), .B2(n_495), .C(n_498), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_502), .B2(n_504), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_515), .C(n_522), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_507), .B(n_510), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_SL g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_531), .Y(n_547) );
INVx1_ASAP7_75t_L g549 ( .A(n_532), .Y(n_549) );
OAI222xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_536), .B1(n_540), .B2(n_542), .C1(n_545), .C2(n_550), .Y(n_533) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
endmodule