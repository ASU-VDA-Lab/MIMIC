module fake_jpeg_23032_n_300 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_19),
.B1(n_18),
.B2(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_54),
.B1(n_36),
.B2(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_26),
.Y(n_78)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_52),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_42),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_56),
.A2(n_23),
.B1(n_31),
.B2(n_25),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_61),
.B(n_71),
.Y(n_94)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_55),
.B1(n_50),
.B2(n_28),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_30),
.B1(n_25),
.B2(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_39),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_68),
.Y(n_101)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_72),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_83),
.B1(n_89),
.B2(n_28),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_24),
.B1(n_36),
.B2(n_37),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_74),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_16),
.B1(n_41),
.B2(n_38),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_33),
.B(n_27),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_58),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_84),
.C(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_42),
.B1(n_35),
.B2(n_16),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_16),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_26),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_16),
.B1(n_20),
.B2(n_32),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_51),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_35),
.B1(n_37),
.B2(n_33),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_47),
.B1(n_27),
.B2(n_17),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_105),
.B1(n_112),
.B2(n_109),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_104),
.Y(n_125)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_0),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_114),
.B(n_65),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_64),
.B(n_55),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_84),
.C(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_75),
.B1(n_70),
.B2(n_68),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_63),
.B1(n_74),
.B2(n_67),
.Y(n_124)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.Y(n_137)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_121),
.B(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_122),
.B(n_127),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_129),
.C(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_137),
.B1(n_133),
.B2(n_144),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_79),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_69),
.B1(n_88),
.B2(n_84),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_128),
.A2(n_136),
.B1(n_143),
.B2(n_146),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_84),
.C(n_91),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_78),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_142),
.B(n_1),
.Y(n_180)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_140),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_89),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_87),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_147),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_29),
.B(n_28),
.C(n_33),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_94),
.B1(n_96),
.B2(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_60),
.C(n_80),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_90),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_94),
.A2(n_33),
.B1(n_27),
.B2(n_17),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_111),
.A3(n_110),
.B1(n_98),
.B2(n_105),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_1),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_147),
.B(n_143),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_160),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_95),
.C(n_117),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_153),
.B(n_157),
.C(n_179),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_106),
.B1(n_100),
.B2(n_95),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_159),
.B1(n_175),
.B2(n_177),
.Y(n_197)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_180),
.B(n_12),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_106),
.C(n_92),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_110),
.C(n_27),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_163),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_92),
.B1(n_115),
.B2(n_104),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_118),
.B(n_2),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_11),
.C(n_15),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_130),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_1),
.CI(n_2),
.CON(n_169),
.SN(n_169)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_172),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_118),
.B(n_2),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_125),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_174),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_128),
.A2(n_119),
.B1(n_90),
.B2(n_102),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_97),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_133),
.A2(n_102),
.B1(n_80),
.B2(n_10),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_97),
.B1(n_3),
.B2(n_4),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_97),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_161),
.B(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_185),
.B(n_191),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_207),
.B1(n_163),
.B2(n_152),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_3),
.Y(n_189)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_3),
.Y(n_193)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_180),
.B(n_175),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_194),
.A2(n_195),
.B(n_201),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_3),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_154),
.B1(n_169),
.B2(n_172),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_4),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

HAxp5_ASAP7_75t_SL g201 ( 
.A(n_162),
.B(n_4),
.CON(n_201),
.SN(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_150),
.B(n_4),
.C(n_5),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_167),
.C(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_203),
.A2(n_206),
.B(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_151),
.A2(n_11),
.B1(n_12),
.B2(n_7),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_SL g237 ( 
.A(n_209),
.B(n_211),
.C(n_212),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_168),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_215),
.A2(n_217),
.B1(n_225),
.B2(n_207),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_203),
.A2(n_179),
.B1(n_176),
.B2(n_153),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_150),
.C(n_157),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_170),
.C(n_158),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_205),
.B(n_169),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_173),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_224),
.B(n_205),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_192),
.A2(n_170),
.B1(n_6),
.B2(n_7),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_227),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_234),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_224),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_194),
.B(n_204),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_244),
.B(n_247),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_236),
.B(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_229),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_246),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_204),
.B(n_184),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_197),
.B1(n_192),
.B2(n_206),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_210),
.Y(n_257)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_184),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_220),
.C(n_214),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_249),
.C(n_233),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_211),
.C(n_218),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_235),
.A2(n_210),
.B1(n_199),
.B2(n_216),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_228),
.B1(n_199),
.B2(n_219),
.Y(n_271)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_258),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_261),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g258 ( 
.A(n_237),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_183),
.B(n_195),
.C(n_187),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_259),
.A2(n_195),
.B1(n_244),
.B2(n_242),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_262),
.A2(n_266),
.B(n_198),
.Y(n_277)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_264),
.A2(n_273),
.B(n_223),
.Y(n_282)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_265),
.B(n_267),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_246),
.B(n_243),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_182),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.C(n_249),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_242),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_213),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_237),
.C(n_239),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_252),
.B1(n_260),
.B2(n_226),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_201),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_275),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_271),
.B(n_261),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_277),
.A2(n_282),
.B(n_262),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_278),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_230),
.C(n_202),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_281),
.C(n_209),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_230),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g283 ( 
.A1(n_274),
.A2(n_272),
.B(n_273),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_284),
.B(n_287),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_189),
.Y(n_292)
);

AO21x1_ASAP7_75t_L g290 ( 
.A1(n_288),
.A2(n_289),
.B(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_282),
.B(n_190),
.Y(n_289)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_290),
.Y(n_294)
);

NOR4xp25_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.C(n_7),
.D(n_8),
.Y(n_295)
);

OAI31xp33_ASAP7_75t_SL g293 ( 
.A1(n_285),
.A2(n_193),
.A3(n_11),
.B(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_295),
.B(n_8),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_291),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_297),
.A2(n_294),
.B1(n_286),
.B2(n_9),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_9),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_9),
.Y(n_300)
);


endmodule