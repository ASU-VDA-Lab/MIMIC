module real_jpeg_3306_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_1),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_1),
.A2(n_36),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_3),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_33),
.B1(n_50),
.B2(n_51),
.Y(n_151)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_24),
.C(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_9),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_9),
.B(n_23),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_9),
.B(n_51),
.C(n_63),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_9),
.B(n_57),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_9),
.B(n_71),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_68),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_12),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_54),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_118),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_81),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_60),
.C(n_73),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_20),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_39),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_40),
.C(n_48),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_22),
.A2(n_29),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_35),
.Y(n_167)
);

AO22x1_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_23)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_25),
.A2(n_26),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_26),
.B(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_31),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_30),
.A2(n_44),
.A3(n_88),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_76),
.Y(n_75)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_31),
.B(n_45),
.Y(n_110)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_43),
.B(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_44),
.A2(n_45),
.B1(n_87),
.B2(n_88),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_56),
.B(n_78),
.Y(n_77)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_51),
.B(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_55),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_55),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_55),
.A2(n_56),
.B1(n_124),
.B2(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_56),
.B(n_80),
.Y(n_126)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_57),
.A2(n_79),
.B(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_60),
.B(n_73),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_69),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_61),
.B(n_72),
.Y(n_103)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_101),
.B(n_103),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_65),
.A2(n_103),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_65),
.A2(n_67),
.B1(n_132),
.B2(n_140),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_70),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_74),
.A2(n_75),
.B1(n_77),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_77),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_105),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_96),
.B2(n_104),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_91),
.Y(n_92)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_91),
.A2(n_126),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_98),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_116),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_172),
.B(n_176),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_161),
.B(n_171),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_142),
.B(n_160),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_135),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_135),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_133),
.B2(n_134),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_130),
.C(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_137),
.B1(n_139),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_154),
.B(n_159),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_149),
.B(n_153),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_147),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_150),
.B(n_152),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_157),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_162),
.B(n_163),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_175),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_175),
.Y(n_176)
);


endmodule