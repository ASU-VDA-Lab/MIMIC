module fake_jpeg_17591_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_4),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_21),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_10),
.A2(n_15),
.B1(n_12),
.B2(n_16),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_20),
.A2(n_24),
.B1(n_13),
.B2(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_6),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_6),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_25),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_24),
.A2(n_15),
.B1(n_13),
.B2(n_16),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_26),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_7),
.B1(n_19),
.B2(n_34),
.Y(n_39)
);

NOR2x1_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_17),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_32),
.B1(n_26),
.B2(n_31),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_19),
.A2(n_7),
.B1(n_9),
.B2(n_25),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_40),
.B(n_41),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_36),
.C(n_40),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_52),
.C(n_48),
.Y(n_54)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_33),
.B1(n_44),
.B2(n_43),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_39),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_49),
.B(n_43),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_34),
.B(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_56),
.C(n_54),
.Y(n_57)
);

AO21x1_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_28),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_33),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_33),
.Y(n_60)
);


endmodule