module real_jpeg_24763_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_22),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_38),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_78),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_1),
.A2(n_35),
.B1(n_142),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_44),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_5),
.A2(n_26),
.B1(n_32),
.B2(n_72),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_72),
.Y(n_142)
);

INVx8_ASAP7_75t_SL g87 ( 
.A(n_6),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_26),
.B1(n_32),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_26),
.B1(n_32),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_53),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_13),
.Y(n_92)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_13),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_107),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_106),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_73),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_18),
.B(n_73),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_51),
.C(n_63),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_19),
.A2(n_20),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_21),
.B(n_34),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.A3(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_22),
.A2(n_23),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_32),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_26),
.A2(n_30),
.B(n_58),
.C(n_117),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_30),
.B(n_59),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_30),
.B(n_48),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_42),
.B(n_45),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_35),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_35),
.A2(n_132),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_36),
.B(n_49),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_36),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_38),
.B1(n_56),
.B2(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_37),
.B(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_43),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_51),
.A2(n_63),
.B1(n_64),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_51),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_52),
.A2(n_54),
.B1(n_60),
.B2(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_54),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_59),
.A2(n_100),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_96),
.B2(n_97),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_93),
.B(n_95),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_105),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_153),
.B(n_159),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_128),
.B(n_152),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_110),
.B(n_118),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_123),
.C(n_124),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_125),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_138),
.B(n_151),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_130),
.B(n_136),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_145),
.B(n_150),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);


endmodule