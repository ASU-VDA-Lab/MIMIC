module fake_jpeg_11081_n_185 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_15),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_35),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_22),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_84),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_0),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_0),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_87),
.Y(n_92)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_67),
.B1(n_70),
.B2(n_59),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_67),
.Y(n_105)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_77),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_63),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_100),
.B(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_65),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_114),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_69),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_121),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_73),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_92),
.B(n_54),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_127),
.Y(n_145)
);

OR2x6_ASAP7_75t_SL g127 ( 
.A(n_107),
.B(n_60),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_70),
.B1(n_66),
.B2(n_71),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_20),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_118),
.A2(n_66),
.B1(n_77),
.B2(n_68),
.Y(n_131)
);

NAND2x1_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_1),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_51),
.C(n_39),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_13),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_143),
.B1(n_10),
.B2(n_12),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_17),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_29),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_9),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_28),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_149),
.Y(n_163)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_34),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_148),
.B(n_134),
.C(n_129),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_9),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_126),
.B(n_128),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_14),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_49),
.A3(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_158),
.C(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_157),
.B1(n_27),
.B2(n_45),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_125),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_160),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_46),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_144),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_172),
.B1(n_153),
.B2(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_167),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_179),
.A2(n_163),
.B1(n_176),
.B2(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_177),
.C(n_163),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_168),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_145),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_169),
.B(n_173),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_168),
.Y(n_185)
);


endmodule