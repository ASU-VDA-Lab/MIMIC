module real_jpeg_7363_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_1),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_1),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_3),
.B(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_3),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_3),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_3),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_3),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_3),
.B(n_141),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_4),
.B(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_4),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_4),
.B(n_294),
.Y(n_293)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_5),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_6),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_6),
.B(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_6),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_6),
.B(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_8),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_8),
.B(n_165),
.Y(n_164)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_10),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_11),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_12),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_12),
.B(n_60),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_12),
.B(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_12),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_12),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_12),
.B(n_238),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_13),
.B(n_87),
.Y(n_214)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_15),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_15),
.B(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_193),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_191),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_149),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_19),
.B(n_149),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_94),
.C(n_131),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_20),
.B(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_55),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_21),
.B(n_56),
.C(n_73),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.C(n_46),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_22),
.B(n_217),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_22),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_27),
.CI(n_31),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_23),
.B(n_27),
.C(n_31),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g230 ( 
.A(n_26),
.Y(n_230)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_30),
.Y(n_277)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_35),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_36),
.A2(n_46),
.B1(n_47),
.B2(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_36),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.C(n_45),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_37),
.A2(n_45),
.B1(n_170),
.B2(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_37),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_39),
.Y(n_37)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_59),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g157 ( 
.A(n_38),
.B(n_158),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_38),
.B(n_172),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_40),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_41),
.B(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_44),
.Y(n_139)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_44),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_44),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_45),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_45),
.Y(n_170)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_215)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_73),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_58),
.B(n_65),
.C(n_70),
.Y(n_182)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_65),
.A2(n_72),
.B1(n_115),
.B2(n_116),
.Y(n_255)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_72),
.B(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_82),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_74),
.B(n_83),
.C(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_81),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_81),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_87),
.Y(n_296)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_88),
.Y(n_273)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_88),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_91),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_91),
.B(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_91),
.B(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_94),
.B(n_131),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_110),
.C(n_112),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_95),
.A2(n_110),
.B1(n_111),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_109),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_102),
.C(n_105),
.Y(n_133)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_100),
.Y(n_235)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_100),
.Y(n_254)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_112),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.C(n_126),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_113),
.A2(n_114),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_127),
.Y(n_324)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_125),
.Y(n_248)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_133),
.B(n_134),
.C(n_148),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_144),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_140),
.C(n_144),
.Y(n_154)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_177),
.B1(n_189),
.B2(n_190),
.Y(n_151)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_167),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_166),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_169),
.B1(n_174),
.B2(n_175),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_171),
.A2(n_173),
.B1(n_245),
.B2(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_173),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_219),
.B(n_332),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_196),
.B(n_198),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_216),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_199),
.A2(n_200),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_203),
.B(n_216),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.C(n_215),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_204),
.B(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_207),
.B(n_215),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_214),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_214),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_326),
.B(n_331),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_311),
.B(n_325),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_268),
.B(n_310),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_256),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_223),
.B(n_256),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_243),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_239),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_225),
.B(n_239),
.C(n_243),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.C(n_236),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_258)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_244),
.B(n_320),
.C(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.C(n_267),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_259),
.A2(n_267),
.B1(n_302),
.B2(n_308),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_304),
.B(n_309),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_289),
.B(n_303),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_278),
.B(n_288),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_286),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_286),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B(n_285),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_291),
.B1(n_297),
.B2(n_298),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_299),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_299),
.Y(n_303)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_293),
.B(n_297),
.Y(n_305)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B(n_302),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_313),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_319),
.C(n_322),
.Y(n_327)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule