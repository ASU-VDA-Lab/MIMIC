module fake_jpeg_17336_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_40),
.B(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_30),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g60 ( 
.A(n_47),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_54),
.B1(n_48),
.B2(n_32),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_64),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_42),
.C(n_33),
.Y(n_63)
);

XNOR2x1_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_39),
.B1(n_43),
.B2(n_38),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_73),
.B(n_78),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_72),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_27),
.B1(n_30),
.B2(n_18),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_57),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx5_ASAP7_75t_SL g104 ( 
.A(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_27),
.B1(n_37),
.B2(n_36),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_29),
.Y(n_114)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_88),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_25),
.B1(n_17),
.B2(n_66),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_35),
.B1(n_42),
.B2(n_52),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_104),
.B1(n_70),
.B2(n_65),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_9),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_18),
.B(n_28),
.C(n_17),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_60),
.A2(n_32),
.B1(n_27),
.B2(n_30),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_32),
.B1(n_104),
.B2(n_67),
.Y(n_124)
);

CKINVDCx12_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_63),
.B(n_21),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_28),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_124),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_69),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_23),
.C(n_16),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_62),
.B1(n_65),
.B2(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_122),
.B(n_128),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_96),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_72),
.B(n_78),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_119),
.B(n_133),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_18),
.B1(n_25),
.B2(n_21),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_102),
.B1(n_95),
.B2(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_79),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_131),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_79),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_90),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_104),
.B1(n_100),
.B2(n_93),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_119),
.B1(n_137),
.B2(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_105),
.A3(n_97),
.B1(n_103),
.B2(n_98),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_147),
.A2(n_148),
.B(n_151),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_117),
.B(n_139),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_123),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_90),
.B(n_108),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_31),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_91),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_161),
.Y(n_192)
);

AOI32xp33_ASAP7_75t_L g159 ( 
.A1(n_118),
.A2(n_103),
.A3(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_31),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_127),
.A2(n_112),
.B1(n_103),
.B2(n_101),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_116),
.B1(n_20),
.B2(n_115),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_107),
.B(n_16),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_0),
.B(n_2),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_116),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_126),
.B(n_23),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_166),
.B1(n_52),
.B2(n_74),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_136),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_42),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_74),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_170),
.B(n_83),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_157),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_174),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_134),
.C(n_128),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_185),
.C(n_188),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_179),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_181),
.B(n_197),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_141),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_193),
.B1(n_162),
.B2(n_161),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_187),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_115),
.C(n_80),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_167),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_199),
.B1(n_169),
.B2(n_166),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_144),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_196),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_145),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_153),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_200),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_145),
.B(n_165),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_31),
.C(n_24),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_140),
.C(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_183),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_208),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_188),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_159),
.B(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_174),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_218),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_165),
.B(n_151),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_230),
.B(n_195),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_225),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_226),
.C(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_229),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_147),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_178),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_155),
.C(n_149),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_164),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_172),
.A2(n_152),
.B(n_10),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_239),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_237),
.Y(n_255)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_218),
.Y(n_260)
);

OAI321xp33_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_173),
.A3(n_172),
.B1(n_197),
.B2(n_182),
.C(n_199),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_202),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_221),
.C(n_228),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_243),
.B(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_213),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_194),
.B(n_186),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_250),
.A2(n_220),
.B(n_214),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_223),
.B1(n_210),
.B2(n_212),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_238),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_257),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_251),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_226),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_266),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_204),
.C(n_230),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_233),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_263),
.A2(n_245),
.B1(n_243),
.B2(n_207),
.Y(n_273)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_205),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_268),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_207),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_252),
.A2(n_239),
.B1(n_231),
.B2(n_242),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_177),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_273),
.B(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_284),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_252),
.A2(n_247),
.B1(n_240),
.B2(n_250),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_269),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_255),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_177),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_255),
.C(n_261),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_288),
.C(n_292),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_258),
.C(n_266),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_272),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_225),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_294),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_248),
.C(n_234),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_215),
.C(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_271),
.B(n_186),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_279),
.B1(n_236),
.B2(n_277),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_274),
.C(n_281),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_24),
.C(n_16),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_301),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_293),
.A2(n_180),
.B1(n_190),
.B2(n_177),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_3),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_9),
.B(n_14),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_312),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_313),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_8),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_306),
.C(n_12),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_7),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_7),
.Y(n_313)
);

OAI21x1_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_308),
.B(n_314),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_303),
.B1(n_299),
.B2(n_309),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_309),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_315),
.A3(n_316),
.B1(n_300),
.B2(n_6),
.C1(n_10),
.C2(n_11),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_5),
.B(n_6),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_11),
.B(n_14),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_14),
.C(n_3),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_4),
.B(n_322),
.Y(n_327)
);


endmodule