module fake_jpeg_24076_n_324 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_25),
.B1(n_21),
.B2(n_19),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_25),
.B1(n_19),
.B2(n_17),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_25),
.B1(n_21),
.B2(n_19),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_20),
.C(n_14),
.Y(n_62)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_29),
.B(n_14),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_10),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_74),
.B1(n_49),
.B2(n_58),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_66),
.B1(n_72),
.B2(n_44),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_20),
.B1(n_13),
.B2(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_70),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_20),
.B1(n_23),
.B2(n_17),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_77),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_84),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_94),
.B1(n_64),
.B2(n_68),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_89),
.Y(n_101)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_61),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_98),
.B(n_71),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_112),
.B1(n_83),
.B2(n_86),
.Y(n_128)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_107),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_44),
.B1(n_52),
.B2(n_43),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_100),
.B1(n_95),
.B2(n_91),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_94),
.B1(n_85),
.B2(n_79),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_28),
.C(n_61),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_119),
.C(n_82),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_28),
.B(n_71),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_33),
.B(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_89),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_73),
.B1(n_40),
.B2(n_57),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_100),
.B1(n_95),
.B2(n_93),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_40),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_59),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_29),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_88),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_127),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_131),
.B1(n_133),
.B2(n_120),
.Y(n_159)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_134),
.B1(n_145),
.B2(n_118),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_92),
.B1(n_43),
.B2(n_100),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_132),
.A2(n_148),
.B(n_101),
.Y(n_162)
);

AOI22x1_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_65),
.B1(n_95),
.B2(n_99),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_88),
.B1(n_43),
.B2(n_52),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_91),
.B(n_88),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_129),
.B(n_130),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_141),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_112),
.C(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_117),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_52),
.B1(n_33),
.B2(n_18),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_170),
.B1(n_134),
.B2(n_125),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_105),
.B1(n_115),
.B2(n_113),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_152),
.A2(n_158),
.B1(n_167),
.B2(n_175),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_119),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_160),
.C(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_115),
.B1(n_120),
.B2(n_107),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g200 ( 
.A1(n_159),
.A2(n_174),
.B1(n_27),
.B2(n_26),
.Y(n_200)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_171),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_162),
.A2(n_176),
.B(n_142),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_122),
.C(n_121),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_168),
.C(n_129),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_122),
.B1(n_111),
.B2(n_110),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_110),
.C(n_18),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_141),
.A2(n_126),
.B1(n_144),
.B2(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_131),
.A2(n_27),
.B1(n_26),
.B2(n_24),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_177),
.A2(n_149),
.B1(n_174),
.B2(n_170),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_176),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_192),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_190),
.C(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_183),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_153),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_187),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_151),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_135),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_195),
.B(n_165),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_142),
.C(n_27),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_201),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_169),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_194),
.B(n_165),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_8),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_202),
.B(n_166),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_174),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_7),
.B(n_1),
.Y(n_202)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_206),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_208),
.A2(n_213),
.B1(n_218),
.B2(n_6),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_182),
.B1(n_201),
.B2(n_196),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_197),
.B1(n_203),
.B2(n_214),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_217),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_158),
.Y(n_214)
);

OR2x6_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_207),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_202),
.Y(n_217)
);

OA21x2_ASAP7_75t_SL g221 ( 
.A1(n_189),
.A2(n_152),
.B(n_154),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_221),
.A2(n_222),
.B(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_175),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_197),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_181),
.C(n_190),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_239),
.C(n_243),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_235),
.B(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_234),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_195),
.Y(n_230)
);

XNOR2x1_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_214),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_191),
.B1(n_178),
.B2(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_223),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_178),
.B1(n_186),
.B2(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_236),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_186),
.C(n_195),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_200),
.B(n_174),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_225),
.A2(n_200),
.B(n_1),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_24),
.C(n_0),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_219),
.B1(n_205),
.B2(n_209),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_12),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_218),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_207),
.C(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_220),
.C(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_215),
.Y(n_250)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_257),
.C(n_243),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_253),
.B(n_246),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_227),
.B1(n_232),
.B2(n_242),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_209),
.C(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_265),
.B(n_7),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_230),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_262),
.B(n_263),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_238),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_7),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_238),
.B(n_264),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_272),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_239),
.B(n_245),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_219),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_278),
.C(n_247),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_6),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_277),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_7),
.B(n_1),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_247),
.A2(n_8),
.B(n_2),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_281),
.Y(n_290)
);

OA21x2_ASAP7_75t_L g281 ( 
.A1(n_253),
.A2(n_9),
.B(n_3),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_248),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_282),
.B(n_286),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_280),
.B(n_260),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_258),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_293),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_251),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_256),
.B1(n_269),
.B2(n_271),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_298),
.B1(n_305),
.B2(n_4),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_289),
.C(n_267),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_299),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_267),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_4),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_287),
.A2(n_281),
.B1(n_262),
.B2(n_277),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g299 ( 
.A(n_284),
.B(n_281),
.C(n_285),
.Y(n_299)
);

NOR2xp67_ASAP7_75t_SL g302 ( 
.A(n_292),
.B(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_12),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_288),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_309),
.B(n_310),
.Y(n_316)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_296),
.B(n_303),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_4),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_301),
.B1(n_300),
.B2(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_5),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_297),
.B(n_312),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_315),
.Y(n_319)
);

OAI322xp33_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_314),
.A3(n_5),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_5),
.B(n_10),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_12),
.CI(n_0),
.CON(n_323),
.SN(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_0),
.B(n_290),
.Y(n_324)
);


endmodule