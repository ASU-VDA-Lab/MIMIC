module fake_jpeg_15565_n_357 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_357);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_357;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_49),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_10),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_56),
.Y(n_67)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_49),
.B(n_26),
.CON(n_68),
.SN(n_68)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_73),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_26),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_71),
.A2(n_34),
.B1(n_20),
.B2(n_26),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_19),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_72),
.B(n_79),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_20),
.B1(n_51),
.B2(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_84),
.B1(n_100),
.B2(n_103),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_51),
.B1(n_54),
.B2(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_111),
.B1(n_36),
.B2(n_21),
.Y(n_136)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_45),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_107),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_51),
.B1(n_47),
.B2(n_46),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_104),
.B1(n_66),
.B2(n_53),
.Y(n_125)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_101),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_74),
.A2(n_38),
.B1(n_34),
.B2(n_46),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_38),
.B1(n_26),
.B2(n_44),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_44),
.B1(n_38),
.B2(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_52),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_52),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_53),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_57),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_112),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_33),
.B1(n_29),
.B2(n_37),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_37),
.Y(n_112)
);

FAx1_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_68),
.CI(n_80),
.CON(n_114),
.SN(n_114)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_120),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_72),
.B1(n_24),
.B2(n_32),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_118),
.B1(n_130),
.B2(n_133),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_41),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_122),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_55),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_69),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_64),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_131),
.C(n_63),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_87),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_137),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_28),
.B1(n_21),
.B2(n_36),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_48),
.C(n_79),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_76),
.B1(n_42),
.B2(n_56),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_140),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_76),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_41),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_86),
.Y(n_155)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_144),
.B(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_85),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_149),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_128),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_94),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_157),
.B1(n_162),
.B2(n_167),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_96),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_157),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_110),
.Y(n_157)
);

XOR2x2_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_56),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_138),
.B(n_132),
.Y(n_192)
);

INVx6_ASAP7_75t_SL g159 ( 
.A(n_121),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_162),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_59),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_110),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_28),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_36),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_59),
.Y(n_165)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_60),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g197 ( 
.A(n_168),
.Y(n_197)
);

CKINVDCx10_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_169),
.Y(n_193)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_164),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_122),
.B1(n_171),
.B2(n_125),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_180),
.B1(n_181),
.B2(n_194),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_126),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_176),
.A2(n_166),
.B1(n_145),
.B2(n_146),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_135),
.B1(n_118),
.B2(n_122),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_177),
.A2(n_178),
.B1(n_30),
.B2(n_23),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_158),
.A2(n_113),
.B1(n_115),
.B2(n_114),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_130),
.B1(n_29),
.B2(n_140),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_131),
.B1(n_133),
.B2(n_138),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_182),
.B(n_163),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_185),
.C(n_155),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_141),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_153),
.A2(n_21),
.B(n_139),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_188),
.A2(n_195),
.B1(n_89),
.B2(n_90),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_151),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_148),
.A2(n_153),
.B1(n_165),
.B2(n_154),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_117),
.B(n_128),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_154),
.A2(n_117),
.B1(n_93),
.B2(n_86),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_202),
.B1(n_145),
.B2(n_161),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_151),
.A2(n_93),
.B1(n_89),
.B2(n_127),
.Y(n_202)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

AO21x2_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_169),
.B(n_144),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_229),
.B1(n_193),
.B2(n_187),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_206),
.B(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_185),
.C(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_218),
.B(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_147),
.C(n_149),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_214),
.Y(n_234)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_215),
.B(n_217),
.Y(n_239)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_156),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_172),
.B(n_150),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_172),
.B(n_159),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_39),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_168),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_226),
.B(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_231),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_168),
.B1(n_60),
.B2(n_2),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_175),
.B(n_188),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_39),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_201),
.B1(n_202),
.B2(n_174),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_233),
.A2(n_236),
.B1(n_244),
.B2(n_255),
.Y(n_280)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_175),
.B(n_183),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_176),
.B(n_183),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_232),
.B1(n_225),
.B2(n_216),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_30),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_221),
.B(n_191),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g255 ( 
.A(n_205),
.B(n_198),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_205),
.A2(n_187),
.B1(n_181),
.B2(n_177),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_257),
.A2(n_227),
.B1(n_224),
.B2(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_173),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_210),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_261),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_206),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_213),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_263),
.C(n_269),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_248),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_240),
.B1(n_259),
.B2(n_236),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_218),
.B1(n_219),
.B2(n_207),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_272),
.B1(n_246),
.B2(n_237),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_SL g268 ( 
.A(n_235),
.B(n_178),
.C(n_211),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_268),
.A2(n_238),
.B(n_239),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_223),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_230),
.C(n_231),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_105),
.C(n_204),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_105),
.C(n_25),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_238),
.B(n_14),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_281),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_277),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_250),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_237),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_265),
.Y(n_289)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_242),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_245),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_255),
.B1(n_253),
.B2(n_247),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_287),
.B1(n_295),
.B2(n_273),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_262),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_260),
.C(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_271),
.A2(n_243),
.B1(n_249),
.B2(n_245),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_292),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_236),
.B1(n_249),
.B2(n_242),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_296),
.A2(n_14),
.B(n_17),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_297),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_263),
.B(n_246),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_267),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_309),
.C(n_310),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_284),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_304),
.B(n_22),
.Y(n_324)
);

OAI321xp33_ASAP7_75t_L g305 ( 
.A1(n_288),
.A2(n_286),
.A3(n_283),
.B1(n_289),
.B2(n_287),
.C(n_295),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_305),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_307),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_274),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_25),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_290),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_313),
.B(n_1),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_30),
.C(n_23),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_316),
.C(n_290),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_30),
.C(n_23),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_298),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_306),
.B1(n_329),
.B2(n_301),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_320),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_25),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_27),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_22),
.C(n_12),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_327),
.C(n_308),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_326),
.B(n_302),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_325),
.A2(n_328),
.B1(n_321),
.B2(n_13),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_309),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_22),
.C(n_12),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_335),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_331),
.A2(n_336),
.B(n_5),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_316),
.C(n_301),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_334),
.C(n_338),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_27),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_329),
.A2(n_6),
.B1(n_16),
.B2(n_3),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_6),
.C(n_16),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_322),
.C(n_5),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_340),
.A2(n_345),
.B(n_4),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_343),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_5),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_338),
.Y(n_348)
);

AOI31xp67_ASAP7_75t_L g345 ( 
.A1(n_336),
.A2(n_3),
.A3(n_4),
.B(n_13),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_348),
.C(n_349),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_332),
.C(n_331),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_341),
.C(n_15),
.Y(n_351)
);

AOI322xp5_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_1),
.A3(n_2),
.B1(n_15),
.B2(n_27),
.C1(n_345),
.C2(n_328),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_352),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_353),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_354),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_355),
.B(n_350),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_356),
.B(n_15),
.Y(n_357)
);


endmodule