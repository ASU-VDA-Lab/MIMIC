module fake_netlist_5_1670_n_1494 (n_137, n_294, n_318, n_380, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_385, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1494);

input n_137;
input n_294;
input n_318;
input n_380;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_385;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1494;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_329),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_160),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_39),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g392 ( 
.A(n_267),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_268),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_205),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_212),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_328),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_315),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_213),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_173),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_171),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_35),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_41),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_92),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_385),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_224),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_196),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_134),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_114),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_144),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_214),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_197),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_111),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_15),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_310),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_67),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_53),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_184),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_159),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_372),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_166),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_68),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_185),
.B(n_190),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_38),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_8),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_294),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_209),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_51),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_79),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_358),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_356),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_136),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_163),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_164),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_20),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_235),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_44),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_128),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_180),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_170),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_65),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_168),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_343),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_251),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_322),
.Y(n_451)
);

BUFx2_ASAP7_75t_SL g452 ( 
.A(n_296),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_331),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_146),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_269),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_98),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_157),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_193),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_241),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_260),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_257),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_186),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_225),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_248),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_342),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_161),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_378),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g468 ( 
.A(n_105),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g469 ( 
.A(n_348),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_66),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_280),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_114),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_202),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_352),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_69),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_347),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_48),
.Y(n_477)
);

NOR2xp67_ASAP7_75t_L g478 ( 
.A(n_221),
.B(n_216),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_218),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_25),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_43),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_240),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_314),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_273),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_25),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_183),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_78),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_201),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_232),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_379),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_277),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_325),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_167),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_226),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_222),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_204),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_361),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_252),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_247),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_261),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_198),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_191),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_68),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_26),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_266),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_341),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_52),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_48),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_206),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_337),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_106),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_22),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_319),
.Y(n_513)
);

HB1xp67_ASAP7_75t_SL g514 ( 
.A(n_5),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_344),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_119),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_249),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_227),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_263),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_386),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_366),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_165),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_375),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_73),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_367),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_194),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_300),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_308),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_211),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_339),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_135),
.Y(n_531)
);

INVxp67_ASAP7_75t_L g532 ( 
.A(n_293),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_318),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_13),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_162),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_250),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_169),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_139),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_23),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_309),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_11),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_297),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_387),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_130),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_228),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_137),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_311),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_220),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_63),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_320),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_324),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_256),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_80),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_103),
.Y(n_554)
);

INVxp67_ASAP7_75t_SL g555 ( 
.A(n_242),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_67),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_1),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_152),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_272),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_254),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_153),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_182),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_357),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_155),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_334),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_229),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_69),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_405),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_390),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_460),
.B(n_0),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_391),
.A2(n_125),
.B(n_124),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_433),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_445),
.Y(n_573)
);

INVxp33_ASAP7_75t_SL g574 ( 
.A(n_390),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_428),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_428),
.B(n_2),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_407),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_417),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_435),
.B(n_3),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_402),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_549),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_445),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_411),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_403),
.B(n_3),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_403),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_404),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_420),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_514),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_588)
);

BUFx12f_ASAP7_75t_L g589 ( 
.A(n_407),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_487),
.A2(n_8),
.B1(n_4),
.B2(n_7),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_445),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_422),
.B(n_439),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_446),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_422),
.B(n_7),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_417),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_455),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_439),
.B(n_9),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_455),
.B(n_126),
.Y(n_600)
);

OA21x2_ASAP7_75t_L g601 ( 
.A1(n_391),
.A2(n_9),
.B(n_10),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_455),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_476),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_435),
.B(n_10),
.Y(n_604)
);

BUFx3_ASAP7_75t_L g605 ( 
.A(n_490),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_466),
.B(n_11),
.Y(n_606)
);

OA21x2_ASAP7_75t_L g607 ( 
.A1(n_414),
.A2(n_12),
.B(n_13),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_442),
.A2(n_15),
.B1(n_12),
.B2(n_14),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_429),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_460),
.B(n_14),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_476),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_476),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_429),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_470),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_504),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_416),
.Y(n_616)
);

CKINVDCx6p67_ASAP7_75t_R g617 ( 
.A(n_389),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_507),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_470),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_541),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_554),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_503),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_624)
);

AO22x1_ASAP7_75t_L g625 ( 
.A1(n_524),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_466),
.B(n_19),
.Y(n_626)
);

OA21x2_ASAP7_75t_L g627 ( 
.A1(n_414),
.A2(n_495),
.B(n_436),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_528),
.B(n_21),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_475),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_419),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_475),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_499),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_499),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_436),
.A2(n_22),
.B(n_24),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_425),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_495),
.A2(n_24),
.B(n_26),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_553),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_499),
.B(n_127),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_530),
.B(n_27),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_434),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_567),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_499),
.Y(n_642)
);

BUFx8_ASAP7_75t_L g643 ( 
.A(n_512),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_490),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_545),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_545),
.B(n_28),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_573),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_544),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_448),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_629),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_585),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_629),
.Y(n_652)
);

BUFx4f_ASAP7_75t_L g653 ( 
.A(n_627),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_600),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_570),
.B(n_610),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_600),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_586),
.B(n_544),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_600),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_573),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_628),
.B(n_396),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_573),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_SL g663 ( 
.A1(n_579),
.A2(n_508),
.B1(n_477),
.B2(n_481),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_582),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_617),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_582),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_587),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_639),
.B(n_584),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_593),
.B(n_536),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_581),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_582),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_635),
.B(n_640),
.Y(n_673)
);

BUFx8_ASAP7_75t_SL g674 ( 
.A(n_581),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_505),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_584),
.B(n_548),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_582),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_570),
.B(n_493),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_615),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_592),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_616),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_592),
.Y(n_683)
);

INVx6_ASAP7_75t_L g684 ( 
.A(n_643),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_592),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_616),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_618),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_597),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_597),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_621),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_605),
.B(n_505),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_597),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_605),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_597),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_574),
.A2(n_502),
.B1(n_492),
.B2(n_393),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_569),
.B(n_572),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_599),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_644),
.B(n_543),
.Y(n_698)
);

XOR2xp5_ASAP7_75t_L g699 ( 
.A(n_630),
.B(n_492),
.Y(n_699)
);

INVx4_ASAP7_75t_L g700 ( 
.A(n_600),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_574),
.A2(n_502),
.B1(n_395),
.B2(n_462),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_655),
.B(n_630),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_699),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_655),
.B(n_579),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_678),
.A2(n_627),
.B1(n_607),
.B2(n_601),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_673),
.B(n_577),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_667),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_653),
.B(n_427),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_651),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_656),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_656),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_661),
.A2(n_610),
.B1(n_424),
.B2(n_525),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_669),
.B(n_590),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_656),
.Y(n_714)
);

BUFx12f_ASAP7_75t_L g715 ( 
.A(n_684),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_677),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_660),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_651),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_668),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_674),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_653),
.B(n_478),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_649),
.B(n_604),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_660),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_654),
.B(n_543),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_669),
.B(n_603),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_677),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_654),
.B(n_550),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_693),
.B(n_595),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_661),
.B(n_604),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_670),
.B(n_603),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_648),
.A2(n_607),
.B1(n_634),
.B2(n_601),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_654),
.B(n_700),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_689),
.B(n_632),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_689),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_696),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_697),
.B(n_633),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_697),
.B(n_646),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_676),
.B(n_606),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_693),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_697),
.B(n_646),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_676),
.B(n_650),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_658),
.B(n_645),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_647),
.B(n_595),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_682),
.A2(n_517),
.B1(n_626),
.B2(n_606),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_647),
.B(n_694),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_700),
.B(n_550),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_662),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_698),
.A2(n_576),
.B(n_626),
.C(n_608),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_660),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_664),
.B(n_598),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_664),
.B(n_575),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_672),
.B(n_575),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_SL g753 ( 
.A(n_665),
.B(n_588),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_679),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_672),
.B(n_599),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_680),
.B(n_599),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_681),
.B(n_602),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_681),
.B(n_602),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_652),
.B(n_675),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_648),
.A2(n_568),
.B1(n_576),
.B2(n_440),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_683),
.B(n_602),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_691),
.B(n_663),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_687),
.A2(n_623),
.B(n_641),
.C(n_622),
.Y(n_763)
);

O2A1O1Ixp5_ASAP7_75t_L g764 ( 
.A1(n_685),
.A2(n_609),
.B(n_631),
.C(n_596),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_657),
.B(n_394),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_685),
.B(n_602),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_690),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_686),
.Y(n_768)
);

O2A1O1Ixp5_ASAP7_75t_L g769 ( 
.A1(n_688),
.A2(n_609),
.B(n_631),
.C(n_596),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_686),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_704),
.B(n_671),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_704),
.B(n_688),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_706),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_702),
.B(n_695),
.Y(n_774)
);

CKINVDCx11_ASAP7_75t_R g775 ( 
.A(n_715),
.Y(n_775)
);

O2A1O1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_729),
.A2(n_738),
.B(n_748),
.C(n_722),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_708),
.A2(n_659),
.B(n_657),
.Y(n_777)
);

O2A1O1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_729),
.A2(n_738),
.B(n_702),
.C(n_762),
.Y(n_778)
);

NOR2x1_ASAP7_75t_L g779 ( 
.A(n_718),
.B(n_648),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_708),
.A2(n_659),
.B(n_657),
.Y(n_780)
);

O2A1O1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_762),
.A2(n_588),
.B(n_418),
.C(n_432),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_721),
.A2(n_659),
.B(n_692),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_721),
.A2(n_636),
.B1(n_634),
.B2(n_600),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_741),
.A2(n_701),
.B1(n_469),
.B2(n_555),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_739),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_705),
.A2(n_571),
.B(n_659),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_728),
.B(n_392),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_724),
.A2(n_447),
.B(n_532),
.C(n_431),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_712),
.B(n_589),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_747),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_759),
.B(n_684),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_728),
.B(n_479),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_735),
.B(n_744),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_732),
.A2(n_694),
.B(n_692),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_L g795 ( 
.A(n_760),
.B(n_591),
.C(n_624),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_732),
.A2(n_725),
.B(n_737),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_768),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_707),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_742),
.B(n_735),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_709),
.B(n_486),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_770),
.B(n_591),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_705),
.B(n_399),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_731),
.A2(n_565),
.B1(n_409),
.B2(n_412),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_730),
.B(n_388),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_717),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_719),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_731),
.B(n_413),
.Y(n_807)
);

AOI22x1_ASAP7_75t_SL g808 ( 
.A1(n_720),
.A2(n_511),
.B1(n_516),
.B2(n_485),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_740),
.A2(n_666),
.B(n_660),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_724),
.A2(n_636),
.B(n_638),
.Y(n_810)
);

A2O1A1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_743),
.A2(n_426),
.B(n_430),
.C(n_421),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_750),
.A2(n_666),
.B(n_612),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_754),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_727),
.A2(n_746),
.B(n_713),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_767),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_727),
.A2(n_438),
.B1(n_441),
.B2(n_437),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_753),
.B(n_580),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_746),
.A2(n_769),
.B(n_764),
.C(n_763),
.Y(n_818)
);

INVx3_ASAP7_75t_SL g819 ( 
.A(n_765),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_703),
.B(n_674),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_717),
.Y(n_821)
);

OA22x2_ASAP7_75t_L g822 ( 
.A1(n_751),
.A2(n_637),
.B1(n_468),
.B2(n_472),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_752),
.B(n_449),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_SL g824 ( 
.A(n_733),
.B(n_548),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_710),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_745),
.A2(n_451),
.B(n_454),
.C(n_450),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_723),
.B(n_456),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_711),
.B(n_594),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_736),
.A2(n_620),
.B(n_611),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_755),
.A2(n_620),
.B(n_611),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_717),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_714),
.A2(n_458),
.B1(n_461),
.B2(n_457),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_716),
.A2(n_464),
.B1(n_465),
.B2(n_463),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_756),
.A2(n_620),
.B(n_611),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_723),
.B(n_467),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_726),
.Y(n_836)
);

AOI21x1_ASAP7_75t_L g837 ( 
.A1(n_757),
.A2(n_474),
.B(n_471),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_749),
.B(n_483),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_758),
.A2(n_642),
.B(n_620),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_749),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_734),
.B(n_484),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_761),
.B(n_480),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_766),
.A2(n_491),
.B1(n_494),
.B2(n_489),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_717),
.A2(n_498),
.B1(n_500),
.B2(n_497),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_747),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_704),
.A2(n_398),
.B1(n_400),
.B2(n_397),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_704),
.B(n_506),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_SL g848 ( 
.A1(n_703),
.A2(n_556),
.B1(n_557),
.B2(n_539),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_708),
.A2(n_642),
.B(n_515),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_704),
.B(n_513),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_708),
.A2(n_642),
.B(n_520),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_718),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_708),
.A2(n_642),
.B(n_521),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_704),
.A2(n_406),
.B1(n_408),
.B2(n_401),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_708),
.A2(n_523),
.B(n_518),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_747),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_704),
.B(n_410),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_527),
.B(n_526),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_704),
.B(n_415),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_747),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_704),
.B(n_423),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_704),
.B(n_531),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_723),
.Y(n_863)
);

HB1xp67_ASAP7_75t_L g864 ( 
.A(n_735),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_708),
.A2(n_535),
.B(n_533),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_708),
.A2(n_540),
.B(n_538),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_704),
.A2(n_552),
.B(n_561),
.C(n_559),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_707),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_704),
.B(n_443),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_704),
.B(n_564),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_704),
.B(n_566),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_718),
.Y(n_872)
);

O2A1O1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_704),
.A2(n_578),
.B(n_614),
.C(n_613),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_708),
.A2(n_453),
.B(n_444),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_706),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_747),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_704),
.A2(n_578),
.B(n_619),
.C(n_614),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_704),
.B(n_459),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_704),
.B(n_638),
.Y(n_879)
);

INVx4_ASAP7_75t_SL g880 ( 
.A(n_819),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_778),
.A2(n_619),
.B(n_452),
.C(n_473),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_828),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_775),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_828),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_776),
.A2(n_488),
.B(n_496),
.C(n_482),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_771),
.B(n_501),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_785),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_786),
.A2(n_510),
.B(n_509),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_799),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_861),
.B(n_519),
.Y(n_890)
);

AO31x2_ASAP7_75t_L g891 ( 
.A1(n_803),
.A2(n_638),
.A3(n_31),
.B(n_29),
.Y(n_891)
);

AO21x2_ASAP7_75t_L g892 ( 
.A1(n_802),
.A2(n_807),
.B(n_814),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_782),
.A2(n_772),
.B(n_809),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_783),
.A2(n_529),
.B(n_522),
.Y(n_894)
);

AO21x2_ASAP7_75t_L g895 ( 
.A1(n_810),
.A2(n_131),
.B(n_129),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_864),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_869),
.A2(n_563),
.B1(n_542),
.B2(n_546),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_878),
.A2(n_547),
.B(n_551),
.C(n_537),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_774),
.A2(n_560),
.B1(n_562),
.B2(n_558),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_773),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_875),
.B(n_30),
.Y(n_901)
);

OAI22x1_ASAP7_75t_L g902 ( 
.A1(n_789),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_818),
.A2(n_133),
.B(n_132),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_805),
.A2(n_140),
.B(n_138),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_817),
.B(n_32),
.Y(n_905)
);

BUFx2_ASAP7_75t_R g906 ( 
.A(n_793),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_801),
.Y(n_907)
);

BUFx2_ASAP7_75t_R g908 ( 
.A(n_857),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_797),
.Y(n_909)
);

AO31x2_ASAP7_75t_L g910 ( 
.A1(n_847),
.A2(n_35),
.A3(n_33),
.B(n_34),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_831),
.A2(n_142),
.B(n_141),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_785),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_852),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_791),
.B(n_33),
.Y(n_914)
);

AO31x2_ASAP7_75t_L g915 ( 
.A1(n_850),
.A2(n_37),
.A3(n_34),
.B(n_36),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_852),
.Y(n_916)
);

BUFx12f_ASAP7_75t_L g917 ( 
.A(n_852),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_798),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_779),
.B(n_143),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_815),
.Y(n_920)
);

AOI221x1_ASAP7_75t_L g921 ( 
.A1(n_862),
.A2(n_148),
.B1(n_149),
.B2(n_147),
.C(n_145),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_870),
.B(n_37),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_777),
.A2(n_151),
.B(n_150),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_871),
.B(n_38),
.Y(n_924)
);

INVxp67_ASAP7_75t_SL g925 ( 
.A(n_821),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_872),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_868),
.Y(n_927)
);

O2A1O1Ixp5_ASAP7_75t_SL g928 ( 
.A1(n_844),
.A2(n_42),
.B(n_39),
.C(n_40),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_784),
.A2(n_44),
.B(n_40),
.C(n_42),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_780),
.A2(n_156),
.B(n_154),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_SL g931 ( 
.A1(n_811),
.A2(n_867),
.B(n_826),
.C(n_816),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_842),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_872),
.B(n_158),
.Y(n_933)
);

AO31x2_ASAP7_75t_L g934 ( 
.A1(n_855),
.A2(n_47),
.A3(n_45),
.B(n_46),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_813),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_872),
.Y(n_936)
);

BUFx2_ASAP7_75t_SL g937 ( 
.A(n_806),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_801),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_820),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_822),
.Y(n_940)
);

AO31x2_ASAP7_75t_L g941 ( 
.A1(n_858),
.A2(n_50),
.A3(n_47),
.B(n_49),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_781),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_827),
.B(n_787),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_846),
.A2(n_174),
.B1(n_175),
.B2(n_172),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_792),
.B(n_53),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_825),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_824),
.B(n_176),
.Y(n_947)
);

AO31x2_ASAP7_75t_L g948 ( 
.A1(n_865),
.A2(n_56),
.A3(n_54),
.B(n_55),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_804),
.A2(n_178),
.B(n_177),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_854),
.B(n_54),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_840),
.A2(n_181),
.B(n_179),
.Y(n_951)
);

INVx5_ASAP7_75t_L g952 ( 
.A(n_863),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_808),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_848),
.Y(n_954)
);

NOR2x1_ASAP7_75t_SL g955 ( 
.A(n_823),
.B(n_187),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_866),
.B(n_56),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_790),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_836),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_835),
.A2(n_189),
.B(n_188),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_800),
.B(n_57),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_845),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_838),
.A2(n_195),
.B(n_192),
.Y(n_962)
);

AO31x2_ASAP7_75t_L g963 ( 
.A1(n_849),
.A2(n_851),
.A3(n_853),
.B(n_843),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_856),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_874),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_SL g966 ( 
.A1(n_788),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_860),
.B(n_61),
.Y(n_967)
);

INVx5_ASAP7_75t_L g968 ( 
.A(n_876),
.Y(n_968)
);

AO31x2_ASAP7_75t_L g969 ( 
.A1(n_832),
.A2(n_63),
.A3(n_61),
.B(n_62),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_812),
.A2(n_200),
.B(n_199),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_873),
.B(n_62),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_877),
.B(n_64),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_841),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_829),
.B(n_64),
.Y(n_974)
);

AOI221x1_ASAP7_75t_L g975 ( 
.A1(n_833),
.A2(n_276),
.B1(n_384),
.B2(n_383),
.C(n_381),
.Y(n_975)
);

AO31x2_ASAP7_75t_L g976 ( 
.A1(n_830),
.A2(n_70),
.A3(n_65),
.B(n_66),
.Y(n_976)
);

AO31x2_ASAP7_75t_L g977 ( 
.A1(n_834),
.A2(n_72),
.A3(n_70),
.B(n_71),
.Y(n_977)
);

OA21x2_ASAP7_75t_L g978 ( 
.A1(n_839),
.A2(n_207),
.B(n_203),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_837),
.Y(n_979)
);

AOI21x1_ASAP7_75t_SL g980 ( 
.A1(n_879),
.A2(n_71),
.B(n_72),
.Y(n_980)
);

OR2x2_ASAP7_75t_L g981 ( 
.A(n_864),
.B(n_73),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_796),
.A2(n_210),
.B(n_208),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_859),
.A2(n_217),
.B1(n_219),
.B2(n_215),
.Y(n_983)
);

AOI221xp5_ASAP7_75t_SL g984 ( 
.A1(n_778),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.C(n_77),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_778),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_859),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_785),
.B(n_223),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_785),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_828),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_799),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_785),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_778),
.A2(n_81),
.B(n_82),
.C(n_83),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_785),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_859),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_778),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_785),
.B(n_230),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_796),
.A2(n_233),
.B(n_231),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_859),
.A2(n_290),
.B1(n_380),
.B2(n_377),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_778),
.A2(n_87),
.B(n_88),
.C(n_89),
.Y(n_999)
);

OAI221xp5_ASAP7_75t_L g1000 ( 
.A1(n_778),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.C(n_90),
.Y(n_1000)
);

OA21x2_ASAP7_75t_L g1001 ( 
.A1(n_786),
.A2(n_236),
.B(n_234),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_796),
.A2(n_238),
.B(n_237),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_828),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_828),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_864),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_796),
.A2(n_243),
.B(n_239),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_796),
.A2(n_245),
.B(n_244),
.Y(n_1007)
);

AND2x6_ASAP7_75t_L g1008 ( 
.A(n_879),
.B(n_246),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_796),
.A2(n_255),
.B(n_253),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_828),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_859),
.B(n_91),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_828),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_775),
.Y(n_1013)
);

AO31x2_ASAP7_75t_L g1014 ( 
.A1(n_803),
.A2(n_93),
.A3(n_94),
.B(n_95),
.Y(n_1014)
);

AO31x2_ASAP7_75t_L g1015 ( 
.A1(n_803),
.A2(n_93),
.A3(n_94),
.B(n_95),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_828),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_796),
.A2(n_259),
.B(n_258),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_859),
.B(n_96),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_828),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_778),
.A2(n_96),
.B(n_97),
.C(n_99),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_785),
.Y(n_1021)
);

NAND3x1_ASAP7_75t_L g1022 ( 
.A(n_795),
.B(n_100),
.C(n_101),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_785),
.B(n_262),
.Y(n_1023)
);

AO32x2_ASAP7_75t_L g1024 ( 
.A1(n_803),
.A2(n_100),
.A3(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_796),
.A2(n_265),
.B(n_264),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_785),
.Y(n_1026)
);

AO21x2_ASAP7_75t_L g1027 ( 
.A1(n_786),
.A2(n_306),
.B(n_374),
.Y(n_1027)
);

NAND2x1_ASAP7_75t_L g1028 ( 
.A(n_991),
.B(n_270),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_943),
.B(n_104),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_905),
.B(n_105),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_1011),
.A2(n_312),
.B1(n_371),
.B2(n_370),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_920),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1005),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_1018),
.A2(n_305),
.B(n_369),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_892),
.A2(n_304),
.B(n_368),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_914),
.B(n_106),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_896),
.B(n_107),
.Y(n_1037)
);

OA21x2_ASAP7_75t_L g1038 ( 
.A1(n_903),
.A2(n_303),
.B(n_365),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_952),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_909),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_889),
.B(n_107),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_927),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_913),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_890),
.A2(n_302),
.B1(n_364),
.B2(n_363),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_973),
.B(n_108),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_888),
.A2(n_301),
.B(n_362),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_922),
.B(n_108),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_924),
.B(n_109),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_990),
.B(n_109),
.Y(n_1049)
);

BUFx2_ASAP7_75t_L g1050 ( 
.A(n_916),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_957),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_900),
.B(n_110),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_887),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_925),
.A2(n_299),
.B(n_360),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1001),
.A2(n_298),
.B(n_359),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_935),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_1027),
.A2(n_295),
.B(n_355),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_940),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_947),
.B(n_112),
.C(n_113),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_961),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_886),
.B(n_113),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_981),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_952),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_932),
.B(n_115),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_883),
.Y(n_1065)
);

OR2x6_ASAP7_75t_L g1066 ( 
.A(n_917),
.B(n_115),
.Y(n_1066)
);

OAI211xp5_ASAP7_75t_L g1067 ( 
.A1(n_986),
.A2(n_116),
.B(n_117),
.C(n_118),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_907),
.Y(n_1068)
);

OA21x2_ASAP7_75t_L g1069 ( 
.A1(n_921),
.A2(n_313),
.B(n_353),
.Y(n_1069)
);

BUFx4_ASAP7_75t_SL g1070 ( 
.A(n_1013),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_882),
.Y(n_1071)
);

AO21x2_ASAP7_75t_L g1072 ( 
.A1(n_982),
.A2(n_292),
.B(n_350),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_880),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_1003),
.Y(n_1074)
);

AO31x2_ASAP7_75t_L g1075 ( 
.A1(n_975),
.A2(n_116),
.A3(n_117),
.B(n_118),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_885),
.A2(n_316),
.B(n_349),
.Y(n_1076)
);

INVx5_ASAP7_75t_L g1077 ( 
.A(n_887),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_988),
.B(n_291),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_912),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_965),
.A2(n_317),
.B1(n_346),
.B2(n_345),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_884),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_938),
.B(n_119),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_937),
.B(n_120),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_901),
.B(n_120),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_967),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_964),
.B(n_121),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_939),
.B(n_121),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_989),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_964),
.B(n_945),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_946),
.B(n_122),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_946),
.B(n_122),
.Y(n_1091)
);

BUFx8_ASAP7_75t_L g1092 ( 
.A(n_912),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_880),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_926),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_926),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_958),
.B(n_123),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1004),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_936),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_881),
.A2(n_321),
.B(n_271),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_936),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_906),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1010),
.B(n_123),
.Y(n_1102)
);

AO21x2_ASAP7_75t_L g1103 ( 
.A1(n_997),
.A2(n_274),
.B(n_275),
.Y(n_1103)
);

INVx6_ASAP7_75t_L g1104 ( 
.A(n_993),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1012),
.B(n_278),
.Y(n_1105)
);

AO21x2_ASAP7_75t_L g1106 ( 
.A1(n_1002),
.A2(n_279),
.B(n_281),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1016),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_993),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1019),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_974),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1006),
.A2(n_282),
.B(n_283),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_958),
.B(n_284),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_968),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_968),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_1026),
.Y(n_1115)
);

CKINVDCx6p67_ASAP7_75t_R g1116 ( 
.A(n_1026),
.Y(n_1116)
);

AO21x2_ASAP7_75t_L g1117 ( 
.A1(n_1007),
.A2(n_285),
.B(n_286),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1009),
.A2(n_287),
.B(n_288),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_SL g1119 ( 
.A(n_960),
.B(n_899),
.C(n_942),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1021),
.B(n_289),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_897),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_933),
.B(n_330),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1017),
.A2(n_333),
.B(n_335),
.Y(n_1123)
);

AO21x2_ASAP7_75t_L g1124 ( 
.A1(n_1025),
.A2(n_338),
.B(n_340),
.Y(n_1124)
);

OAI21xp33_ASAP7_75t_SL g1125 ( 
.A1(n_994),
.A2(n_971),
.B(n_956),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_987),
.B(n_1023),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_996),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_980),
.A2(n_951),
.B(n_904),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_984),
.A2(n_894),
.B(n_985),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_908),
.B(n_954),
.Y(n_1130)
);

NOR2x1_ASAP7_75t_SL g1131 ( 
.A(n_895),
.B(n_972),
.Y(n_1131)
);

BUFx8_ASAP7_75t_L g1132 ( 
.A(n_1024),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_919),
.B(n_898),
.Y(n_1133)
);

AO21x1_ASAP7_75t_L g1134 ( 
.A1(n_995),
.A2(n_999),
.B(n_944),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_992),
.A2(n_1020),
.A3(n_955),
.B(n_929),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_928),
.A2(n_949),
.B(n_911),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_972),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_983),
.A2(n_998),
.B1(n_1022),
.B2(n_1000),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_959),
.A2(n_962),
.B(n_930),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_919),
.B(n_1008),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1008),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_970),
.A2(n_923),
.B(n_891),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_902),
.B(n_978),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_919),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_963),
.A2(n_1008),
.B(n_931),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_910),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_953),
.B(n_1014),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_963),
.A2(n_891),
.B(n_948),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_966),
.A2(n_1015),
.B(n_1014),
.Y(n_1149)
);

HB1xp67_ASAP7_75t_L g1150 ( 
.A(n_934),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_1024),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_934),
.B(n_941),
.Y(n_1152)
);

AO21x2_ASAP7_75t_L g1153 ( 
.A1(n_941),
.A2(n_948),
.B(n_976),
.Y(n_1153)
);

OR2x6_ASAP7_75t_L g1154 ( 
.A(n_969),
.B(n_977),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_915),
.A2(n_893),
.B(n_794),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_L g1156 ( 
.A(n_950),
.B(n_702),
.C(n_778),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_903),
.A2(n_786),
.B(n_979),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_943),
.B(n_704),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_918),
.Y(n_1159)
);

AOI21xp33_ASAP7_75t_L g1160 ( 
.A1(n_1011),
.A2(n_778),
.B(n_859),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_918),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_918),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_887),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_892),
.A2(n_653),
.B(n_732),
.Y(n_1164)
);

OAI21xp33_ASAP7_75t_SL g1165 ( 
.A1(n_903),
.A2(n_783),
.B(n_1018),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1005),
.Y(n_1166)
);

AO21x2_ASAP7_75t_L g1167 ( 
.A1(n_903),
.A2(n_888),
.B(n_721),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_887),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_893),
.A2(n_794),
.B(n_786),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_921),
.A2(n_975),
.A3(n_979),
.B(n_985),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1011),
.A2(n_778),
.B(n_704),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_889),
.B(n_990),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_889),
.B(n_774),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_889),
.B(n_774),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_893),
.A2(n_794),
.B(n_786),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1032),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1032),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1094),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1158),
.B(n_1171),
.Y(n_1179)
);

AO21x2_ASAP7_75t_L g1180 ( 
.A1(n_1160),
.A2(n_1149),
.B(n_1136),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1173),
.B(n_1174),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1033),
.B(n_1166),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1042),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1043),
.B(n_1126),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1159),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1089),
.B(n_1156),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1159),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1092),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1060),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1060),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1064),
.B(n_1062),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1161),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1041),
.B(n_1049),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1145),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1102),
.B(n_1029),
.Y(n_1195)
);

INVxp67_ASAP7_75t_SL g1196 ( 
.A(n_1132),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1162),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1077),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1040),
.B(n_1137),
.Y(n_1199)
);

BUFx8_ASAP7_75t_SL g1200 ( 
.A(n_1065),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1068),
.B(n_1083),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1056),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1056),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1088),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1092),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1045),
.B(n_1081),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1107),
.B(n_1097),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1139),
.A2(n_1167),
.B(n_1099),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1039),
.B(n_1063),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1169),
.A2(n_1175),
.B(n_1164),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1109),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1094),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1109),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1051),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1071),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1079),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1131),
.A2(n_1076),
.B(n_1046),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1074),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1172),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1130),
.B(n_1037),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1150),
.Y(n_1221)
);

AO21x2_ASAP7_75t_L g1222 ( 
.A1(n_1131),
.A2(n_1128),
.B(n_1153),
.Y(n_1222)
);

INVx2_ASAP7_75t_SL g1223 ( 
.A(n_1104),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1087),
.B(n_1052),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1085),
.B(n_1082),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1110),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1110),
.Y(n_1227)
);

OR2x2_ASAP7_75t_L g1228 ( 
.A(n_1047),
.B(n_1048),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1086),
.Y(n_1229)
);

AO21x2_ASAP7_75t_L g1230 ( 
.A1(n_1152),
.A2(n_1057),
.B(n_1034),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1090),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1085),
.B(n_1132),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1091),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1152),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_R g1235 ( 
.A(n_1157),
.B(n_1144),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1039),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1063),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1146),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1096),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1127),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1127),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1030),
.B(n_1095),
.Y(n_1242)
);

OA21x2_ASAP7_75t_L g1243 ( 
.A1(n_1035),
.A2(n_1055),
.B(n_1134),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1151),
.B(n_1125),
.Y(n_1244)
);

OR2x4_ASAP7_75t_L g1245 ( 
.A(n_1147),
.B(n_1119),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1111),
.A2(n_1118),
.B(n_1123),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1165),
.A2(n_1061),
.B(n_1138),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1098),
.Y(n_1248)
);

AND2x4_ASAP7_75t_L g1249 ( 
.A(n_1108),
.B(n_1077),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1151),
.B(n_1036),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1115),
.B(n_1058),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1084),
.B(n_1105),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1112),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_SL g1254 ( 
.A1(n_1038),
.A2(n_1133),
.B(n_1069),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1135),
.B(n_1170),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1113),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1114),
.Y(n_1257)
);

OR2x2_ASAP7_75t_SL g1258 ( 
.A(n_1059),
.B(n_1093),
.Y(n_1258)
);

AO21x2_ASAP7_75t_L g1259 ( 
.A1(n_1140),
.A2(n_1106),
.B(n_1124),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1154),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1104),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1154),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1077),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1163),
.Y(n_1264)
);

AO21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1080),
.A2(n_1075),
.B(n_1067),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1163),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1116),
.Y(n_1267)
);

INVxp67_ASAP7_75t_L g1268 ( 
.A(n_1168),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1028),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1168),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1168),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1129),
.A2(n_1143),
.B(n_1142),
.Y(n_1272)
);

OR2x2_ASAP7_75t_L g1273 ( 
.A(n_1101),
.B(n_1100),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1122),
.Y(n_1274)
);

INVx1_ASAP7_75t_SL g1275 ( 
.A(n_1050),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1053),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1066),
.B(n_1073),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1066),
.B(n_1078),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1141),
.B(n_1129),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1120),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1135),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_SL g1282 ( 
.A1(n_1121),
.A2(n_1031),
.B(n_1044),
.C(n_1141),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1075),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1072),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1103),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1117),
.B(n_1054),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1070),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1173),
.B(n_1174),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1182),
.Y(n_1289)
);

OAI211xp5_ASAP7_75t_L g1290 ( 
.A1(n_1247),
.A2(n_1233),
.B(n_1229),
.C(n_1231),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1189),
.Y(n_1291)
);

INVxp67_ASAP7_75t_SL g1292 ( 
.A(n_1189),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1213),
.B(n_1195),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1179),
.B(n_1203),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1216),
.Y(n_1295)
);

INVxp33_ASAP7_75t_L g1296 ( 
.A(n_1181),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1176),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1190),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1179),
.B(n_1226),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1288),
.B(n_1252),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1177),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1183),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1186),
.B(n_1228),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1225),
.B(n_1232),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1185),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1190),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1187),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1250),
.B(n_1244),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1207),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1227),
.B(n_1250),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1244),
.B(n_1255),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1247),
.B(n_1204),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1202),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1211),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1232),
.B(n_1214),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1192),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1219),
.B(n_1239),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1197),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1206),
.B(n_1224),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1234),
.B(n_1196),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1215),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1218),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1193),
.B(n_1242),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1196),
.B(n_1281),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1221),
.Y(n_1325)
);

OR2x6_ASAP7_75t_L g1326 ( 
.A(n_1260),
.B(n_1262),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1253),
.B(n_1251),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1238),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1248),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1274),
.B(n_1265),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1280),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1279),
.B(n_1180),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1283),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1256),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1267),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1201),
.B(n_1191),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1272),
.B(n_1184),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1267),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1184),
.B(n_1278),
.Y(n_1339)
);

BUFx2_ASAP7_75t_SL g1340 ( 
.A(n_1205),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1257),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1264),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1266),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1184),
.B(n_1220),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1240),
.B(n_1241),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1270),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1236),
.B(n_1237),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1273),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1284),
.B(n_1285),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1178),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1245),
.B(n_1209),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1303),
.B(n_1304),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1293),
.B(n_1245),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1320),
.B(n_1222),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1327),
.A2(n_1217),
.B1(n_1230),
.B2(n_1208),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1325),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1291),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1312),
.B(n_1208),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1298),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1320),
.B(n_1269),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1300),
.B(n_1308),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1312),
.B(n_1194),
.Y(n_1364)
);

CKINVDCx16_ASAP7_75t_R g1365 ( 
.A(n_1336),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1306),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1307),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_1292),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1293),
.B(n_1199),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1333),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1297),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1330),
.B(n_1249),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1315),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1332),
.B(n_1217),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1301),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1302),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1323),
.Y(n_1377)
);

NAND2xp33_ASAP7_75t_L g1378 ( 
.A(n_1331),
.B(n_1286),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1315),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1296),
.B(n_1268),
.Y(n_1380)
);

AND2x4_ASAP7_75t_SL g1381 ( 
.A(n_1350),
.B(n_1249),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1310),
.B(n_1210),
.Y(n_1382)
);

OR2x2_ASAP7_75t_L g1383 ( 
.A(n_1308),
.B(n_1258),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1319),
.B(n_1275),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1337),
.B(n_1294),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1305),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1313),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1314),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1327),
.B(n_1289),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1336),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1296),
.B(n_1276),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1299),
.B(n_1277),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1330),
.B(n_1326),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1344),
.B(n_1268),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1317),
.B(n_1198),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1309),
.B(n_1198),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1290),
.A2(n_1243),
.B1(n_1286),
.B2(n_1246),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1377),
.B(n_1353),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1393),
.B(n_1347),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1385),
.B(n_1348),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1385),
.B(n_1348),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1374),
.B(n_1311),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1370),
.Y(n_1403)
);

HB1xp67_ASAP7_75t_L g1404 ( 
.A(n_1359),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1360),
.B(n_1311),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1367),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1371),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1375),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1374),
.B(n_1351),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1363),
.B(n_1344),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1376),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1354),
.B(n_1324),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1359),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1386),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1373),
.B(n_1324),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1379),
.B(n_1339),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1390),
.B(n_1339),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1387),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1393),
.B(n_1326),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1388),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1366),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1389),
.B(n_1316),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1395),
.B(n_1318),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1398),
.A2(n_1383),
.B1(n_1365),
.B2(n_1355),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1400),
.B(n_1364),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1403),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1403),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1407),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1404),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1406),
.Y(n_1430)
);

AOI21xp33_ASAP7_75t_L g1431 ( 
.A1(n_1422),
.A2(n_1391),
.B(n_1326),
.Y(n_1431)
);

AOI21xp33_ASAP7_75t_L g1432 ( 
.A1(n_1423),
.A2(n_1326),
.B(n_1384),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1401),
.B(n_1356),
.Y(n_1433)
);

INVx2_ASAP7_75t_SL g1434 ( 
.A(n_1413),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1419),
.A2(n_1393),
.B1(n_1410),
.B2(n_1417),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1416),
.B(n_1368),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1408),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1412),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1411),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1402),
.B(n_1361),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1409),
.B(n_1382),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1409),
.B(n_1382),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1414),
.Y(n_1443)
);

OAI211xp5_ASAP7_75t_L g1444 ( 
.A1(n_1431),
.A2(n_1357),
.B(n_1421),
.C(n_1396),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1424),
.A2(n_1369),
.B(n_1392),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1426),
.Y(n_1446)
);

NOR4xp25_ASAP7_75t_SL g1447 ( 
.A(n_1432),
.B(n_1235),
.C(n_1358),
.D(n_1418),
.Y(n_1447)
);

NAND4xp25_ASAP7_75t_L g1448 ( 
.A(n_1436),
.B(n_1380),
.C(n_1328),
.D(n_1394),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1429),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1427),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1426),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1428),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1434),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1437),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1438),
.B(n_1402),
.Y(n_1455)
);

AOI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1439),
.A2(n_1420),
.B(n_1378),
.C(n_1329),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1430),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1430),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1443),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1435),
.A2(n_1399),
.B1(n_1419),
.B2(n_1372),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1440),
.Y(n_1461)
);

AOI222xp33_ASAP7_75t_L g1462 ( 
.A1(n_1445),
.A2(n_1357),
.B1(n_1341),
.B2(n_1334),
.C1(n_1381),
.C2(n_1349),
.Y(n_1462)
);

AOI211xp5_ASAP7_75t_L g1463 ( 
.A1(n_1444),
.A2(n_1378),
.B(n_1434),
.C(n_1419),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1449),
.B(n_1441),
.Y(n_1464)
);

AOI211xp5_ASAP7_75t_L g1465 ( 
.A1(n_1460),
.A2(n_1282),
.B(n_1338),
.C(n_1295),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1461),
.A2(n_1399),
.B1(n_1372),
.B2(n_1362),
.Y(n_1466)
);

OAI21xp33_ASAP7_75t_L g1467 ( 
.A1(n_1448),
.A2(n_1405),
.B(n_1415),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1456),
.A2(n_1338),
.B(n_1361),
.C(n_1295),
.Y(n_1468)
);

AOI21xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1468),
.A2(n_1287),
.B(n_1453),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1467),
.B(n_1200),
.Y(n_1470)
);

AOI322xp5_ASAP7_75t_L g1471 ( 
.A1(n_1464),
.A2(n_1449),
.A3(n_1455),
.B1(n_1442),
.B2(n_1441),
.C1(n_1425),
.C2(n_1433),
.Y(n_1471)
);

NOR4xp25_ASAP7_75t_L g1472 ( 
.A(n_1463),
.B(n_1459),
.C(n_1454),
.D(n_1452),
.Y(n_1472)
);

XNOR2xp5_ASAP7_75t_L g1473 ( 
.A(n_1465),
.B(n_1188),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1472),
.A2(n_1462),
.B(n_1205),
.C(n_1282),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1469),
.A2(n_1466),
.B1(n_1450),
.B2(n_1340),
.C(n_1451),
.Y(n_1475)
);

NAND4xp75_ASAP7_75t_L g1476 ( 
.A(n_1470),
.B(n_1346),
.C(n_1343),
.D(n_1342),
.Y(n_1476)
);

NAND4xp25_ASAP7_75t_L g1477 ( 
.A(n_1471),
.B(n_1397),
.C(n_1349),
.D(n_1372),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_SL g1478 ( 
.A(n_1473),
.Y(n_1478)
);

NAND4xp25_ASAP7_75t_L g1479 ( 
.A(n_1470),
.B(n_1321),
.C(n_1322),
.D(n_1345),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1476),
.B(n_1442),
.Y(n_1480)
);

NOR3xp33_ASAP7_75t_SL g1481 ( 
.A(n_1475),
.B(n_1235),
.C(n_1200),
.Y(n_1481)
);

OAI211xp5_ASAP7_75t_L g1482 ( 
.A1(n_1474),
.A2(n_1447),
.B(n_1254),
.C(n_1457),
.Y(n_1482)
);

OR4x2_ASAP7_75t_L g1483 ( 
.A(n_1481),
.B(n_1478),
.C(n_1477),
.D(n_1479),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1480),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1483),
.A2(n_1335),
.B1(n_1263),
.B2(n_1482),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1485),
.A2(n_1484),
.B1(n_1483),
.B2(n_1399),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1486),
.A2(n_1484),
.B1(n_1223),
.B2(n_1261),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1486),
.Y(n_1488)
);

OAI21xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1487),
.A2(n_1457),
.B(n_1458),
.Y(n_1489)
);

AOI21xp33_ASAP7_75t_L g1490 ( 
.A1(n_1488),
.A2(n_1345),
.B(n_1352),
.Y(n_1490)
);

XOR2xp5_ASAP7_75t_L g1491 ( 
.A(n_1490),
.B(n_1212),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1489),
.B(n_1446),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1492),
.A2(n_1458),
.B(n_1446),
.Y(n_1493)
);

AOI21xp33_ASAP7_75t_L g1494 ( 
.A1(n_1493),
.A2(n_1491),
.B(n_1212),
.Y(n_1494)
);


endmodule