module fake_jpeg_1106_n_197 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_14),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_39),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_6),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx11_ASAP7_75t_SL g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_59),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_60),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_85),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_59),
.B1(n_65),
.B2(n_51),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_84),
.B1(n_60),
.B2(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_67),
.B1(n_65),
.B2(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_55),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_67),
.B1(n_66),
.B2(n_68),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_92),
.A2(n_76),
.B1(n_64),
.B2(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_105),
.Y(n_114)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_100),
.B1(n_103),
.B2(n_109),
.Y(n_117)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_73),
.B(n_79),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_102),
.B(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_89),
.A2(n_64),
.B1(n_71),
.B2(n_68),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_70),
.B1(n_63),
.B2(n_56),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_58),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_0),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_111),
.B(n_80),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_82),
.B1(n_98),
.B2(n_103),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_113),
.A2(n_26),
.B1(n_44),
.B2(n_43),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_112),
.C(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_25),
.C(n_47),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_85),
.A3(n_80),
.B1(n_52),
.B2(n_73),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_73),
.B1(n_62),
.B2(n_61),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_129),
.B(n_6),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_22),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_73),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_113),
.B(n_117),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_52),
.B1(n_1),
.B2(n_3),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_18),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_SL g132 ( 
.A(n_94),
.B(n_52),
.C(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_1),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_134),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_5),
.Y(n_134)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_23),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_141),
.C(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_21),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_17),
.C(n_38),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_19),
.C(n_46),
.Y(n_143)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_114),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_147),
.B(n_148),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_157),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_5),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_156),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_119),
.B(n_127),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_7),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_171),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_164),
.A2(n_165),
.B(n_168),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_138),
.A2(n_28),
.B(n_41),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_143),
.C(n_170),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_155),
.B(n_138),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_146),
.B(n_144),
.C(n_141),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_137),
.B(n_9),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_177),
.C(n_178),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_150),
.B1(n_139),
.B2(n_135),
.C(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_169),
.B1(n_163),
.B2(n_159),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_11),
.B(n_12),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_31),
.C(n_35),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_180),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_184),
.Y(n_188)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_162),
.C(n_168),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_161),
.C(n_172),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_29),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_176),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_189),
.A2(n_190),
.B1(n_33),
.B2(n_48),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_189),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_188),
.B(n_191),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_185),
.C(n_184),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_34),
.Y(n_197)
);


endmodule