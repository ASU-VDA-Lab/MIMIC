module fake_jpeg_14963_n_148 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_148);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_17),
.Y(n_54)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_45),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_25),
.B(n_18),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_19),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_25),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_28),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_16),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_27),
.B1(n_23),
.B2(n_15),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_21),
.B1(n_19),
.B2(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_54),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_57),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_60),
.Y(n_79)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_28),
.B(n_38),
.C(n_24),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_76),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_68),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_26),
.B1(n_17),
.B2(n_21),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_69),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_26),
.B1(n_29),
.B2(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_72),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_10),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_41),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_43),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_55),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_90),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_55),
.B(n_47),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_65),
.C(n_61),
.Y(n_95)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_77),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_42),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_95),
.B(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_89),
.A2(n_75),
.B1(n_62),
.B2(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_100),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_64),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_102),
.C(n_108),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_53),
.B1(n_72),
.B2(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_76),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_60),
.B1(n_77),
.B2(n_63),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_92),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_51),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_51),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_104),
.B(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_83),
.C(n_93),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_119),
.C(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_91),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_86),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_103),
.B1(n_80),
.B2(n_88),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_2),
.B(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_86),
.B1(n_95),
.B2(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_113),
.B(n_119),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_4),
.C(n_5),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_131),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_111),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_132),
.A2(n_122),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_138),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_127),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.C(n_133),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_131),
.B(n_125),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_144),
.B(n_12),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_134),
.A3(n_4),
.B1(n_5),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_144)
);

AOI21x1_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_140),
.B(n_11),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_146),
.Y(n_148)
);


endmodule