module fake_jpeg_5916_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

HB1xp67_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx24_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_14),
.B(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g17 ( 
.A1(n_8),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_12),
.B1(n_13),
.B2(n_10),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_19),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

AO21x1_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_17),
.B(n_14),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_29),
.A2(n_23),
.B1(n_16),
.B2(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_24),
.B(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_18),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_25),
.C(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_31),
.C(n_29),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_27),
.C(n_28),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_22),
.B1(n_13),
.B2(n_27),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_10),
.B(n_11),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_21),
.B(n_11),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_21),
.B1(n_40),
.B2(n_5),
.Y(n_43)
);


endmodule