module real_jpeg_4898_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_249;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_244;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_127;
wire n_53;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_2),
.A2(n_39),
.B1(n_67),
.B2(n_69),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_39),
.B1(n_80),
.B2(n_83),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_39),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_2),
.B(n_69),
.C(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_178),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_2),
.A2(n_185),
.B(n_187),
.C(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_2),
.B(n_199),
.C(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_2),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_2),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_18),
.Y(n_226)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_7),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_7),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_58),
.B1(n_91),
.B2(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_8),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_9),
.A2(n_93),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_10),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_10),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_170),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_168),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_146),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_14),
.B(n_146),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_120),
.C(n_132),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_15),
.B(n_120),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_70),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_16),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_16),
.A2(n_134),
.B1(n_166),
.B2(n_249),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_41),
.Y(n_16)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_17),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_17),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_17),
.B(n_145),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_17),
.A2(n_133),
.B1(n_181),
.B2(n_192),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_17),
.B(n_95),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_28),
.B(n_37),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_29),
.Y(n_28)
);

AO22x1_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_24),
.Y(n_190)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_39),
.A2(n_55),
.B(n_58),
.Y(n_187)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_41),
.A2(n_133),
.B(n_134),
.C(n_144),
.Y(n_132)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_41),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_41),
.A2(n_95),
.B1(n_130),
.B2(n_145),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_41),
.A2(n_145),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

AO21x2_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_54),
.B(n_66),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_54),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_43)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_44),
.Y(n_186)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_54),
.Y(n_178)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_60),
.B2(n_63),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_70),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_95),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_71),
.A2(n_95),
.B1(n_130),
.B2(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_71),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_78),
.B1(n_85),
.B2(n_87),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_87),
.B1(n_122),
.B2(n_126),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_72),
.B(n_76),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_74),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_121),
.B1(n_130),
.B2(n_131),
.Y(n_120)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_95),
.B(n_121),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_95),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_95),
.A2(n_130),
.B1(n_177),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_95),
.A2(n_130),
.B1(n_196),
.B2(n_197),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_95),
.A2(n_130),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_95),
.A2(n_145),
.B(n_183),
.C(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_95),
.B(n_145),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g201 ( 
.A(n_98),
.Y(n_201)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

NAND2x1_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_103),
.A2(n_112),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_103),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B1(n_108),
.B2(n_111),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_104),
.B(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_119),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_116),
.Y(n_200)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_177),
.C(n_179),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_130),
.B(n_222),
.C(n_229),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_132),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_134),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_142),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_179),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_142),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_142),
.A2(n_179),
.B1(n_184),
.B2(n_191),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_142),
.B(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_142),
.A2(n_179),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_142),
.B(n_184),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_142),
.B(n_145),
.C(n_225),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

AND3x1_ASAP7_75t_L g255 ( 
.A(n_144),
.B(n_232),
.C(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_164),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_163),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_244),
.B(n_262),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_234),
.B(n_243),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_220),
.B(n_233),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_193),
.B(n_219),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_179),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_179),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_192),
.Y(n_180)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_205),
.B(n_218),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_202),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_213),
.Y(n_206)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_230),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_230),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_236),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_257),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_254),
.C(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_260),
.Y(n_264)
);


endmodule