module fake_netlist_1_2427_n_1580 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1580);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1580;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_613;
wire n_648;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_659;
wire n_432;
wire n_386;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1518;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_261), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_272), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_78), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_316), .Y(n_352) );
BUFx2_ASAP7_75t_SL g353 ( .A(n_334), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_36), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_16), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_221), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_245), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_183), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_229), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_15), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_247), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_337), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_69), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_309), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_319), .Y(n_366) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_282), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_246), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_133), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_199), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_153), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_206), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_48), .Y(n_373) );
BUFx10_ASAP7_75t_L g374 ( .A(n_160), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_277), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_323), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_190), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_264), .Y(n_378) );
INVxp33_ASAP7_75t_SL g379 ( .A(n_310), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_139), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_222), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_160), .Y(n_382) );
CKINVDCx20_ASAP7_75t_R g383 ( .A(n_149), .Y(n_383) );
CKINVDCx14_ASAP7_75t_R g384 ( .A(n_28), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_211), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_269), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_32), .Y(n_387) );
BUFx3_ASAP7_75t_L g388 ( .A(n_72), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_240), .Y(n_389) );
INVxp33_ASAP7_75t_L g390 ( .A(n_46), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_250), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_82), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_214), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_216), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_96), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_27), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_174), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_65), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_313), .Y(n_400) );
CKINVDCx14_ASAP7_75t_R g401 ( .A(n_31), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_326), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_307), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_275), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_179), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_52), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_332), .Y(n_407) );
INVxp33_ASAP7_75t_L g408 ( .A(n_202), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_136), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_278), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_103), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_254), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_267), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_77), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_283), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_178), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_317), .Y(n_417) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_290), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_268), .Y(n_419) );
INVxp67_ASAP7_75t_SL g420 ( .A(n_50), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_265), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_152), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_61), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_239), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_145), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_180), .Y(n_426) );
BUFx5_ASAP7_75t_L g427 ( .A(n_80), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_195), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_339), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_292), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_208), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_56), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_133), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_166), .B(n_24), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_14), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_340), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_103), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_342), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_324), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_140), .Y(n_440) );
NOR2xp67_ASAP7_75t_L g441 ( .A(n_284), .B(n_297), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_279), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_241), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_223), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_14), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_26), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_286), .Y(n_447) );
BUFx2_ASAP7_75t_L g448 ( .A(n_251), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_87), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_50), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_113), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g452 ( .A(n_263), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_236), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_194), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_122), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_45), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_118), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_8), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_287), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_338), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_234), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_35), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_57), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_293), .B(n_253), .Y(n_464) );
INVxp67_ASAP7_75t_L g465 ( .A(n_196), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_12), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_34), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_242), .B(n_299), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_207), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_141), .Y(n_470) );
CKINVDCx14_ASAP7_75t_R g471 ( .A(n_6), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_101), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_70), .Y(n_473) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_300), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_96), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_25), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_105), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_114), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_285), .Y(n_479) );
CKINVDCx5p33_ASAP7_75t_R g480 ( .A(n_94), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_235), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_244), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_31), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_43), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_298), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_67), .Y(n_486) );
CKINVDCx14_ASAP7_75t_R g487 ( .A(n_71), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_203), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_5), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_29), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_197), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_101), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_32), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_219), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_301), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_306), .Y(n_496) );
INVxp67_ASAP7_75t_SL g497 ( .A(n_64), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_140), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_147), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_170), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_105), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_225), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_227), .Y(n_503) );
BUFx8_ASAP7_75t_SL g504 ( .A(n_34), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_118), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_3), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_172), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_112), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_325), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_188), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_330), .Y(n_511) );
NOR2xp67_ASAP7_75t_L g512 ( .A(n_40), .B(n_335), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_321), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_204), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_173), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_38), .Y(n_516) );
BUFx5_ASAP7_75t_L g517 ( .A(n_1), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_30), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_348), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_64), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_276), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_259), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_143), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_248), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_12), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_84), .Y(n_526) );
INVxp67_ASAP7_75t_SL g527 ( .A(n_60), .Y(n_527) );
INVxp67_ASAP7_75t_SL g528 ( .A(n_75), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_4), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_3), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_198), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_66), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_314), .B(n_121), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_142), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_8), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_419), .Y(n_536) );
INVx2_ASAP7_75t_SL g537 ( .A(n_402), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_448), .B(n_0), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_402), .B(n_0), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_427), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_402), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_427), .Y(n_542) );
AND2x6_ASAP7_75t_L g543 ( .A(n_375), .B(n_177), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_384), .A2(n_4), .B1(n_1), .B2(n_2), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_390), .B(n_2), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_384), .A2(n_7), .B1(n_5), .B2(n_6), .Y(n_546) );
BUFx8_ASAP7_75t_L g547 ( .A(n_427), .Y(n_547) );
NOR2x1_ASAP7_75t_L g548 ( .A(n_363), .B(n_7), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_401), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_427), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_427), .Y(n_551) );
OA21x2_ASAP7_75t_L g552 ( .A1(n_442), .A2(n_182), .B(n_181), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_401), .Y(n_553) );
INVx5_ASAP7_75t_L g554 ( .A(n_375), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_378), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_410), .Y(n_556) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_442), .A2(n_185), .B(n_184), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_427), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_427), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_390), .B(n_9), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_517), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_471), .Y(n_562) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_391), .B(n_186), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
AND2x2_ASAP7_75t_SL g565 ( .A(n_403), .B(n_347), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_373), .B(n_9), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_517), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_410), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_517), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_373), .B(n_10), .Y(n_570) );
XNOR2x1_ASAP7_75t_L g571 ( .A(n_409), .B(n_458), .Y(n_571) );
INVx6_ASAP7_75t_L g572 ( .A(n_517), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_408), .B(n_10), .Y(n_574) );
INVx4_ASAP7_75t_L g575 ( .A(n_363), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
AND2x4_ASAP7_75t_L g577 ( .A(n_382), .B(n_11), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_432), .B(n_11), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_555), .B(n_408), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_542), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_545), .A2(n_487), .B1(n_471), .B2(n_354), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_555), .B(n_487), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_553), .B(n_445), .Y(n_583) );
INVxp67_ASAP7_75t_SL g584 ( .A(n_547), .Y(n_584) );
NOR2x1_ASAP7_75t_L g585 ( .A(n_538), .B(n_387), .Y(n_585) );
BUFx3_ASAP7_75t_L g586 ( .A(n_547), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_563), .A2(n_486), .B1(n_367), .B2(n_376), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_571), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_571), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_553), .B(n_400), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_562), .B(n_409), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_539), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_539), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_562), .B(n_458), .Y(n_595) );
BUFx10_ASAP7_75t_L g596 ( .A(n_539), .Y(n_596) );
INVx4_ASAP7_75t_L g597 ( .A(n_539), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_540), .Y(n_598) );
INVx4_ASAP7_75t_SL g599 ( .A(n_543), .Y(n_599) );
BUFx4f_ASAP7_75t_L g600 ( .A(n_543), .Y(n_600) );
INVx4_ASAP7_75t_L g601 ( .A(n_543), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_574), .B(n_476), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_557), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_536), .B(n_465), .Y(n_604) );
INVx5_ASAP7_75t_L g605 ( .A(n_543), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_537), .B(n_379), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_574), .B(n_476), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_537), .B(n_379), .Y(n_609) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_543), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_540), .Y(n_611) );
INVx4_ASAP7_75t_L g612 ( .A(n_543), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g614 ( .A1(n_544), .A2(n_480), .B1(n_518), .B2(n_506), .Y(n_614) );
INVx4_ASAP7_75t_L g615 ( .A(n_543), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_547), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_551), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_558), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_574), .B(n_480), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_547), .B(n_357), .C(n_350), .Y(n_620) );
INVx4_ASAP7_75t_L g621 ( .A(n_586), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_583), .B(n_571), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_583), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_602), .B(n_578), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_606), .B(n_538), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_579), .B(n_545), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_587), .Y(n_627) );
NOR2xp33_ASAP7_75t_R g628 ( .A(n_586), .B(n_549), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_581), .A2(n_565), .B1(n_563), .B2(n_545), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_597), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_597), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_609), .B(n_560), .Y(n_632) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_586), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_582), .B(n_563), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_608), .B(n_560), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_619), .B(n_560), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_585), .B(n_565), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_597), .A2(n_565), .B1(n_570), .B2(n_566), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_585), .B(n_566), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_597), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_591), .B(n_592), .Y(n_641) );
AO22x1_ASAP7_75t_L g642 ( .A1(n_588), .A2(n_520), .B1(n_518), .B2(n_566), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_616), .B(n_566), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_595), .B(n_575), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_589), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_589), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_593), .B(n_578), .Y(n_647) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_616), .B(n_577), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_593), .B(n_575), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_590), .Y(n_650) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_616), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_594), .B(n_566), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_594), .Y(n_653) );
NAND2x1p5_ASAP7_75t_L g654 ( .A(n_594), .B(n_577), .Y(n_654) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_601), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_584), .B(n_570), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_601), .B(n_570), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_596), .B(n_570), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_614), .A2(n_546), .B1(n_544), .B2(n_577), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_596), .B(n_577), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_596), .Y(n_661) );
BUFx3_ASAP7_75t_L g662 ( .A(n_600), .Y(n_662) );
INVx3_ASAP7_75t_L g663 ( .A(n_603), .Y(n_663) );
INVx4_ASAP7_75t_L g664 ( .A(n_605), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_598), .B(n_577), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_604), .B(n_349), .Y(n_666) );
NAND2xp33_ASAP7_75t_SL g667 ( .A(n_601), .B(n_352), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_599), .B(n_478), .Y(n_668) );
INVx8_ASAP7_75t_L g669 ( .A(n_605), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_599), .B(n_546), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_580), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_600), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_600), .A2(n_610), .B(n_603), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_620), .A2(n_558), .B1(n_564), .B2(n_561), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_580), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_598), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_611), .B(n_349), .Y(n_677) );
BUFx4f_ASAP7_75t_L g678 ( .A(n_603), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_601), .B(n_607), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_599), .B(n_374), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_620), .A2(n_352), .B1(n_376), .B2(n_367), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_613), .B(n_370), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_613), .B(n_370), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_603), .B(n_520), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_610), .A2(n_564), .B1(n_576), .B2(n_541), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_607), .B(n_576), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_617), .Y(n_687) );
AND2x4_ASAP7_75t_L g688 ( .A(n_599), .B(n_548), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_618), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_607), .B(n_405), .Y(n_690) );
BUFx6f_ASAP7_75t_L g691 ( .A(n_607), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_610), .A2(n_541), .B1(n_550), .B2(n_542), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_612), .A2(n_541), .B1(n_550), .B2(n_542), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_612), .Y(n_694) );
AND2x4_ASAP7_75t_SL g695 ( .A(n_612), .B(n_430), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_615), .B(n_482), .Y(n_696) );
A2O1A1Ixp33_ASAP7_75t_L g697 ( .A1(n_605), .A2(n_557), .B(n_559), .C(n_550), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_615), .B(n_482), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_615), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_615), .B(n_559), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_605), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_623), .B(n_383), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_695), .Y(n_703) );
INVx5_ASAP7_75t_L g704 ( .A(n_633), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_645), .Y(n_705) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_621), .B(n_605), .Y(n_706) );
O2A1O1Ixp5_ASAP7_75t_L g707 ( .A1(n_678), .A2(n_474), .B(n_418), .C(n_533), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_678), .A2(n_605), .B(n_557), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_631), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_633), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_646), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_624), .B(n_450), .Y(n_712) );
NOR2x1_ASAP7_75t_L g713 ( .A(n_670), .B(n_430), .Y(n_713) );
AND3x1_ASAP7_75t_L g714 ( .A(n_659), .B(n_548), .C(n_435), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_700), .A2(n_552), .B(n_559), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_621), .B(n_488), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_634), .A2(n_438), .B1(n_444), .B2(n_436), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_634), .A2(n_438), .B1(n_444), .B2(n_436), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_640), .Y(n_719) );
OA22x2_ASAP7_75t_L g720 ( .A1(n_650), .A2(n_435), .B1(n_437), .B2(n_383), .Y(n_720) );
O2A1O1Ixp33_ASAP7_75t_L g721 ( .A1(n_626), .A2(n_434), .B(n_497), .C(n_420), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_700), .A2(n_552), .B(n_567), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_670), .A2(n_572), .B1(n_388), .B2(n_397), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_653), .Y(n_724) );
BUFx8_ASAP7_75t_L g725 ( .A(n_622), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_625), .B(n_396), .Y(n_726) );
AO21x1_ASAP7_75t_L g727 ( .A1(n_637), .A2(n_359), .B(n_358), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_638), .A2(n_513), .B1(n_521), .B2(n_510), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_638), .A2(n_629), .B1(n_695), .B2(n_654), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_625), .B(n_399), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_641), .B(n_504), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_654), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_686), .A2(n_552), .B(n_567), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_635), .B(n_433), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_641), .B(n_568), .C(n_556), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_636), .B(n_440), .Y(n_736) );
INVx1_ASAP7_75t_SL g737 ( .A(n_684), .Y(n_737) );
INVx6_ASAP7_75t_L g738 ( .A(n_639), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_632), .B(n_504), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_647), .A2(n_513), .B1(n_521), .B2(n_510), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_640), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_681), .B(n_437), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_656), .A2(n_522), .B1(n_457), .B2(n_490), .Y(n_743) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_651), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_686), .A2(n_552), .B(n_569), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_630), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_683), .B(n_462), .Y(n_747) );
AOI21x1_ASAP7_75t_L g748 ( .A1(n_657), .A2(n_552), .B(n_573), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_627), .A2(n_522), .B1(n_457), .B2(n_490), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_679), .A2(n_364), .B(n_361), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_688), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_683), .B(n_466), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_679), .A2(n_366), .B(n_365), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g754 ( .A(n_642), .B(n_528), .C(n_527), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_666), .B(n_451), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_657), .A2(n_372), .B(n_368), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_689), .Y(n_757) );
OR2x6_ASAP7_75t_L g758 ( .A(n_648), .B(n_353), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_651), .B(n_488), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_651), .B(n_495), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_666), .B(n_467), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_689), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_L g763 ( .A1(n_652), .A2(n_355), .B(n_360), .C(n_351), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_649), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_676), .A2(n_455), .B(n_526), .C(n_388), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_639), .B(n_495), .Y(n_766) );
INVx4_ASAP7_75t_L g767 ( .A(n_669), .Y(n_767) );
NOR2xp33_ASAP7_75t_R g768 ( .A(n_667), .B(n_451), .Y(n_768) );
OAI22xp5_ASAP7_75t_SL g769 ( .A1(n_648), .A2(n_516), .B1(n_369), .B2(n_380), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_677), .B(n_516), .Y(n_770) );
AO22x2_ASAP7_75t_L g771 ( .A1(n_688), .A2(n_371), .B1(n_398), .B2(n_393), .Y(n_771) );
A2O1A1Ixp33_ASAP7_75t_L g772 ( .A1(n_687), .A2(n_665), .B(n_658), .C(n_660), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_682), .B(n_374), .Y(n_773) );
AND2x4_ASAP7_75t_L g774 ( .A(n_680), .B(n_406), .Y(n_774) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_655), .Y(n_775) );
OR2x2_ASAP7_75t_L g776 ( .A(n_668), .B(n_414), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_628), .B(n_374), .Y(n_777) );
AND2x4_ASAP7_75t_L g778 ( .A(n_661), .B(n_422), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_643), .A2(n_572), .B1(n_526), .B2(n_455), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_644), .B(n_423), .Y(n_780) );
BUFx2_ASAP7_75t_L g781 ( .A(n_628), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_643), .A2(n_572), .B1(n_446), .B2(n_449), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_671), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_675), .B(n_425), .Y(n_784) );
INVx4_ASAP7_75t_L g785 ( .A(n_669), .Y(n_785) );
O2A1O1Ixp33_ASAP7_75t_L g786 ( .A1(n_697), .A2(n_463), .B(n_470), .C(n_456), .Y(n_786) );
NAND2xp33_ASAP7_75t_SL g787 ( .A(n_655), .B(n_362), .Y(n_787) );
O2A1O1Ixp5_ASAP7_75t_L g788 ( .A1(n_673), .A2(n_469), .B(n_511), .C(n_459), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_685), .B(n_472), .Y(n_789) );
A2O1A1Ixp33_ASAP7_75t_L g790 ( .A1(n_674), .A2(n_475), .B(n_477), .C(n_473), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_663), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g792 ( .A1(n_694), .A2(n_381), .B(n_377), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_699), .A2(n_389), .B(n_385), .Y(n_793) );
BUFx12f_ASAP7_75t_L g794 ( .A(n_664), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_690), .B(n_484), .Y(n_795) );
A2O1A1Ixp33_ASAP7_75t_L g796 ( .A1(n_674), .A2(n_492), .B(n_493), .C(n_489), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_692), .A2(n_499), .B(n_500), .C(n_498), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_685), .A2(n_572), .B1(n_543), .B2(n_505), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_664), .Y(n_799) );
INVx3_ASAP7_75t_L g800 ( .A(n_662), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_655), .B(n_386), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_692), .B(n_501), .Y(n_802) );
A2O1A1Ixp33_ASAP7_75t_SL g803 ( .A1(n_693), .A2(n_464), .B(n_469), .C(n_459), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_655), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_696), .A2(n_404), .B(n_395), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_698), .B(n_507), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_662), .B(n_508), .Y(n_807) );
NOR2xp33_ASAP7_75t_R g808 ( .A(n_669), .B(n_392), .Y(n_808) );
O2A1O1Ixp33_ASAP7_75t_L g809 ( .A1(n_672), .A2(n_523), .B(n_525), .C(n_515), .Y(n_809) );
NOR2xp33_ASAP7_75t_SL g810 ( .A(n_672), .B(n_394), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_691), .A2(n_412), .B(n_407), .Y(n_811) );
BUFx2_ASAP7_75t_L g812 ( .A(n_691), .Y(n_812) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_691), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_691), .A2(n_701), .B1(n_530), .B2(n_534), .Y(n_814) );
INVx5_ASAP7_75t_L g815 ( .A(n_633), .Y(n_815) );
A2O1A1Ixp33_ASAP7_75t_L g816 ( .A1(n_634), .A2(n_529), .B(n_535), .C(n_512), .Y(n_816) );
NAND2xp33_ASAP7_75t_SL g817 ( .A(n_638), .B(n_452), .Y(n_817) );
INVx2_ASAP7_75t_L g818 ( .A(n_631), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_678), .A2(n_415), .B(n_413), .Y(n_819) );
BUFx8_ASAP7_75t_L g820 ( .A(n_623), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_645), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_678), .A2(n_417), .B(n_416), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_631), .Y(n_823) );
NAND2x1p5_ASAP7_75t_L g824 ( .A(n_621), .B(n_411), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_678), .A2(n_424), .B(n_421), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_673), .A2(n_514), .B(n_511), .Y(n_826) );
CKINVDCx8_ASAP7_75t_R g827 ( .A(n_670), .Y(n_827) );
INVxp67_ASAP7_75t_L g828 ( .A(n_623), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_634), .A2(n_426), .B1(n_431), .B2(n_429), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_631), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_623), .B(n_356), .Y(n_831) );
NAND3xp33_ASAP7_75t_L g832 ( .A(n_816), .B(n_568), .C(n_556), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_731), .B(n_428), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_784), .Y(n_834) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_755), .B(n_481), .Y(n_835) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_772), .A2(n_443), .B(n_439), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_733), .A2(n_453), .B(n_447), .Y(n_837) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_745), .A2(n_461), .B(n_454), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_778), .Y(n_839) );
A2O1A1Ixp33_ASAP7_75t_L g840 ( .A1(n_786), .A2(n_485), .B(n_491), .C(n_479), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_757), .Y(n_841) );
AOI21xp5_ASAP7_75t_L g842 ( .A1(n_715), .A2(n_496), .B(n_494), .Y(n_842) );
CKINVDCx12_ASAP7_75t_R g843 ( .A(n_769), .Y(n_843) );
O2A1O1Ixp33_ASAP7_75t_SL g844 ( .A1(n_803), .A2(n_503), .B(n_509), .C(n_502), .Y(n_844) );
NOR2xp33_ASAP7_75t_SL g845 ( .A(n_767), .B(n_460), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_778), .Y(n_846) );
NOR2xp33_ASAP7_75t_SL g847 ( .A(n_767), .B(n_554), .Y(n_847) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_740), .A2(n_532), .B1(n_483), .B2(n_554), .Y(n_848) );
INVx3_ASAP7_75t_L g849 ( .A(n_785), .Y(n_849) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_728), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g851 ( .A(n_810), .B(n_531), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_705), .Y(n_852) );
NAND2x1p5_ASAP7_75t_L g853 ( .A(n_785), .B(n_483), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_711), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_732), .B(n_441), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g856 ( .A1(n_722), .A2(n_524), .B(n_519), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_724), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_762), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_820), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_751), .B(n_468), .Y(n_860) );
INVx8_ASAP7_75t_L g861 ( .A(n_758), .Y(n_861) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_820), .Y(n_862) );
OAI21xp5_ASAP7_75t_L g863 ( .A1(n_788), .A2(n_514), .B(n_554), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_740), .A2(n_532), .B1(n_483), .B2(n_554), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_821), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_829), .B(n_532), .Y(n_866) );
BUFx2_ASAP7_75t_L g867 ( .A(n_768), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_708), .A2(n_554), .B(n_556), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g869 ( .A1(n_717), .A2(n_554), .B1(n_568), .B2(n_556), .Y(n_869) );
O2A1O1Ixp33_ASAP7_75t_L g870 ( .A1(n_790), .A2(n_16), .B(n_13), .C(n_15), .Y(n_870) );
OAI222xp33_ASAP7_75t_L g871 ( .A1(n_717), .A2(n_554), .B1(n_17), .B2(n_18), .C1(n_19), .C2(n_20), .Y(n_871) );
O2A1O1Ixp33_ASAP7_75t_SL g872 ( .A1(n_765), .A2(n_797), .B(n_796), .C(n_806), .Y(n_872) );
AO21x2_ASAP7_75t_L g873 ( .A1(n_826), .A2(n_568), .B(n_189), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_L g874 ( .A1(n_795), .A2(n_568), .B(n_18), .C(n_13), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_709), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_829), .B(n_737), .Y(n_876) );
A2O1A1Ixp33_ASAP7_75t_L g877 ( .A1(n_805), .A2(n_568), .B(n_20), .C(n_17), .Y(n_877) );
OAI222xp33_ASAP7_75t_L g878 ( .A1(n_718), .A2(n_19), .B1(n_21), .B2(n_22), .C1(n_23), .C2(n_24), .Y(n_878) );
OAI22x1_ASAP7_75t_L g879 ( .A1(n_718), .A2(n_23), .B1(n_21), .B2(n_22), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g880 ( .A1(n_706), .A2(n_191), .B(n_187), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_748), .A2(n_193), .B(n_192), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_738), .Y(n_882) );
OAI22x1_ASAP7_75t_L g883 ( .A1(n_713), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_738), .Y(n_884) );
AO31x2_ASAP7_75t_L g885 ( .A1(n_727), .A2(n_30), .A3(n_28), .B(n_29), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_702), .B(n_33), .Y(n_886) );
NOR2xp33_ASAP7_75t_L g887 ( .A(n_739), .B(n_770), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_743), .A2(n_36), .B1(n_33), .B2(n_35), .Y(n_888) );
INVxp67_ASAP7_75t_SL g889 ( .A(n_749), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_776), .Y(n_890) );
AOI221xp5_ASAP7_75t_SL g891 ( .A1(n_763), .A2(n_37), .B1(n_38), .B2(n_39), .C(n_40), .Y(n_891) );
AO31x2_ASAP7_75t_L g892 ( .A1(n_729), .A2(n_42), .A3(n_39), .B(n_41), .Y(n_892) );
AO32x2_ASAP7_75t_L g893 ( .A1(n_769), .A2(n_41), .A3(n_42), .B1(n_43), .B2(n_44), .Y(n_893) );
AO31x2_ASAP7_75t_L g894 ( .A1(n_780), .A2(n_47), .A3(n_45), .B(n_46), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_737), .A2(n_51), .B1(n_48), .B2(n_49), .Y(n_895) );
BUFx3_ASAP7_75t_L g896 ( .A(n_794), .Y(n_896) );
NAND2xp5_ASAP7_75t_SL g897 ( .A(n_810), .B(n_828), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_742), .A2(n_52), .B1(n_49), .B2(n_51), .Y(n_898) );
INVx1_ASAP7_75t_SL g899 ( .A(n_781), .Y(n_899) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_758), .Y(n_900) );
O2A1O1Ixp33_ASAP7_75t_L g901 ( .A1(n_721), .A2(n_55), .B(n_53), .C(n_54), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_758), .Y(n_902) );
AO21x2_ASAP7_75t_L g903 ( .A1(n_735), .A2(n_201), .B(n_200), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_774), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_726), .B(n_53), .Y(n_905) );
O2A1O1Ixp33_ASAP7_75t_SL g906 ( .A1(n_759), .A2(n_209), .B(n_210), .C(n_205), .Y(n_906) );
A2O1A1Ixp33_ASAP7_75t_L g907 ( .A1(n_809), .A2(n_56), .B(n_54), .C(n_55), .Y(n_907) );
AO21x1_ASAP7_75t_L g908 ( .A1(n_817), .A2(n_213), .B(n_212), .Y(n_908) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_764), .A2(n_217), .B(n_215), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_723), .A2(n_59), .B1(n_57), .B2(n_58), .Y(n_910) );
AO32x2_ASAP7_75t_L g911 ( .A1(n_782), .A2(n_58), .A3(n_59), .B1(n_60), .B2(n_61), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_719), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_818), .Y(n_913) );
CKINVDCx12_ASAP7_75t_R g914 ( .A(n_777), .Y(n_914) );
BUFx3_ASAP7_75t_L g915 ( .A(n_725), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g916 ( .A1(n_750), .A2(n_220), .B(n_218), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_824), .A2(n_65), .B1(n_62), .B2(n_63), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_823), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g919 ( .A1(n_756), .A2(n_226), .B(n_224), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_730), .B(n_62), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_754), .A2(n_63), .B1(n_66), .B2(n_67), .Y(n_921) );
AOI21xp5_ASAP7_75t_L g922 ( .A1(n_753), .A2(n_230), .B(n_228), .Y(n_922) );
O2A1O1Ixp33_ASAP7_75t_L g923 ( .A1(n_734), .A2(n_68), .B(n_69), .C(n_71), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_774), .A2(n_68), .B1(n_72), .B2(n_73), .Y(n_924) );
O2A1O1Ixp33_ASAP7_75t_SL g925 ( .A1(n_760), .A2(n_346), .B(n_345), .C(n_344), .Y(n_925) );
O2A1O1Ixp33_ASAP7_75t_L g926 ( .A1(n_736), .A2(n_73), .B(n_74), .C(n_75), .Y(n_926) );
AO31x2_ASAP7_75t_L g927 ( .A1(n_819), .A2(n_74), .A3(n_76), .B(n_77), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_824), .A2(n_76), .B1(n_78), .B2(n_79), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_808), .Y(n_929) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_798), .A2(n_232), .B(n_231), .Y(n_930) );
AO21x1_ASAP7_75t_L g931 ( .A1(n_822), .A2(n_237), .B(n_233), .Y(n_931) );
AOI21xp5_ASAP7_75t_L g932 ( .A1(n_783), .A2(n_243), .B(n_238), .Y(n_932) );
O2A1O1Ixp33_ASAP7_75t_L g933 ( .A1(n_747), .A2(n_79), .B(n_80), .C(n_81), .Y(n_933) );
OAI21x1_ASAP7_75t_L g934 ( .A1(n_811), .A2(n_252), .B(n_249), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_792), .A2(n_256), .B(n_255), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_714), .A2(n_81), .B1(n_82), .B2(n_83), .C(n_84), .Y(n_936) );
AO31x2_ASAP7_75t_L g937 ( .A1(n_825), .A2(n_83), .A3(n_85), .B(n_86), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_712), .B(n_85), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_771), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_752), .A2(n_258), .B(n_257), .Y(n_940) );
O2A1O1Ixp33_ASAP7_75t_SL g941 ( .A1(n_791), .A2(n_343), .B(n_341), .C(n_336), .Y(n_941) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_714), .B(n_86), .C(n_87), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_707), .A2(n_88), .B(n_89), .C(n_90), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_771), .Y(n_944) );
A2O1A1Ixp33_ASAP7_75t_L g945 ( .A1(n_773), .A2(n_88), .B(n_89), .C(n_90), .Y(n_945) );
NOR2xp33_ASAP7_75t_SL g946 ( .A(n_704), .B(n_260), .Y(n_946) );
BUFx2_ASAP7_75t_L g947 ( .A(n_703), .Y(n_947) );
A2O1A1Ixp33_ASAP7_75t_L g948 ( .A1(n_807), .A2(n_91), .B(n_92), .C(n_93), .Y(n_948) );
O2A1O1Ixp33_ASAP7_75t_L g949 ( .A1(n_761), .A2(n_91), .B(n_92), .C(n_93), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_746), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_802), .B(n_94), .Y(n_951) );
OAI22xp33_ASAP7_75t_L g952 ( .A1(n_720), .A2(n_95), .B1(n_97), .B2(n_98), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_793), .A2(n_95), .B(n_98), .C(n_99), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_827), .B(n_99), .Y(n_954) );
AO31x2_ASAP7_75t_L g955 ( .A1(n_789), .A2(n_100), .A3(n_102), .B(n_104), .Y(n_955) );
NOR2xp67_ASAP7_75t_R g956 ( .A(n_704), .B(n_102), .Y(n_956) );
AOI221x1_ASAP7_75t_L g957 ( .A1(n_814), .A2(n_831), .B1(n_787), .B2(n_710), .C(n_744), .Y(n_957) );
O2A1O1Ixp33_ASAP7_75t_L g958 ( .A1(n_766), .A2(n_104), .B(n_106), .C(n_107), .Y(n_958) );
OAI21x1_ASAP7_75t_L g959 ( .A1(n_800), .A2(n_333), .B(n_329), .Y(n_959) );
INVx4_ASAP7_75t_L g960 ( .A(n_704), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_741), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g962 ( .A(n_725), .B(n_106), .Y(n_962) );
OAI21x1_ASAP7_75t_L g963 ( .A1(n_800), .A2(n_328), .B(n_327), .Y(n_963) );
O2A1O1Ixp33_ASAP7_75t_SL g964 ( .A1(n_716), .A2(n_322), .B(n_320), .C(n_318), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_830), .Y(n_965) );
AOI21xp5_ASAP7_75t_L g966 ( .A1(n_804), .A2(n_312), .B(n_311), .Y(n_966) );
A2O1A1Ixp33_ASAP7_75t_L g967 ( .A1(n_779), .A2(n_107), .B(n_108), .C(n_109), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_801), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_815), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_799), .Y(n_970) );
O2A1O1Ixp33_ASAP7_75t_SL g971 ( .A1(n_815), .A2(n_308), .B(n_305), .C(n_304), .Y(n_971) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_812), .A2(n_110), .B1(n_111), .B2(n_112), .Y(n_972) );
OAI21xp5_ASAP7_75t_L g973 ( .A1(n_815), .A2(n_303), .B(n_302), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_775), .B(n_111), .Y(n_974) );
INVx2_ASAP7_75t_SL g975 ( .A(n_775), .Y(n_975) );
CKINVDCx5p33_ASAP7_75t_R g976 ( .A(n_775), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_813), .Y(n_977) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_710), .A2(n_296), .B(n_295), .Y(n_978) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_744), .A2(n_294), .B(n_291), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_744), .A2(n_289), .B(n_288), .Y(n_980) );
AO31x2_ASAP7_75t_L g981 ( .A1(n_813), .A2(n_113), .A3(n_114), .B(n_115), .Y(n_981) );
NOR2xp33_ASAP7_75t_SL g982 ( .A(n_813), .B(n_262), .Y(n_982) );
INVx3_ASAP7_75t_SL g983 ( .A(n_758), .Y(n_983) );
BUFx3_ASAP7_75t_L g984 ( .A(n_820), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_702), .B(n_115), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g986 ( .A1(n_731), .A2(n_116), .B1(n_117), .B2(n_119), .C(n_120), .Y(n_986) );
INVx3_ASAP7_75t_L g987 ( .A(n_767), .Y(n_987) );
AND2x4_ASAP7_75t_L g988 ( .A(n_767), .B(n_116), .Y(n_988) );
INVx1_ASAP7_75t_SL g989 ( .A(n_737), .Y(n_989) );
AO31x2_ASAP7_75t_L g990 ( .A1(n_908), .A2(n_117), .A3(n_119), .B(n_120), .Y(n_990) );
INVx2_ASAP7_75t_L g991 ( .A(n_841), .Y(n_991) );
AOI21xp5_ASAP7_75t_L g992 ( .A1(n_837), .A2(n_281), .B(n_280), .Y(n_992) );
INVx3_ASAP7_75t_L g993 ( .A(n_960), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_852), .Y(n_994) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_989), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_854), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_834), .B(n_121), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_857), .Y(n_998) );
A2O1A1Ixp33_ASAP7_75t_L g999 ( .A1(n_887), .A2(n_942), .B(n_901), .C(n_958), .Y(n_999) );
INVx2_ASAP7_75t_L g1000 ( .A(n_858), .Y(n_1000) );
AND2x4_ASAP7_75t_L g1001 ( .A(n_849), .B(n_122), .Y(n_1001) );
AOI21xp5_ASAP7_75t_L g1002 ( .A1(n_838), .A2(n_274), .B(n_273), .Y(n_1002) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_876), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_1003) );
INVx1_ASAP7_75t_SL g1004 ( .A(n_989), .Y(n_1004) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_861), .A2(n_123), .B1(n_124), .B2(n_125), .Y(n_1005) );
AOI222xp33_ASAP7_75t_L g1006 ( .A1(n_889), .A2(n_126), .B1(n_127), .B2(n_128), .C1(n_129), .C2(n_130), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_865), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_939), .A2(n_126), .B1(n_127), .B2(n_128), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_944), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_890), .B(n_862), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_842), .A2(n_271), .B(n_270), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_961), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_850), .B(n_129), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_950), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_904), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_942), .A2(n_130), .B1(n_131), .B2(n_132), .Y(n_1016) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_849), .B(n_131), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_886), .B(n_134), .Y(n_1018) );
AOI22xp5_ASAP7_75t_L g1019 ( .A1(n_859), .A2(n_134), .B1(n_135), .B2(n_136), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_988), .Y(n_1020) );
BUFx12f_ASAP7_75t_L g1021 ( .A(n_984), .Y(n_1021) );
OAI21xp5_ASAP7_75t_L g1022 ( .A1(n_840), .A2(n_135), .B(n_137), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_861), .A2(n_137), .B1(n_138), .B2(n_139), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_896), .B(n_138), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_875), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_839), .B(n_141), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_861), .A2(n_936), .B1(n_867), .B2(n_848), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_846), .B(n_142), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_988), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_985), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_983), .B(n_143), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_905), .B(n_144), .Y(n_1032) );
AO31x2_ASAP7_75t_L g1033 ( .A1(n_931), .A2(n_144), .A3(n_145), .B(n_146), .Y(n_1033) );
OAI21x1_ASAP7_75t_L g1034 ( .A1(n_881), .A2(n_266), .B(n_147), .Y(n_1034) );
AO21x2_ASAP7_75t_L g1035 ( .A1(n_873), .A2(n_148), .B(n_149), .Y(n_1035) );
CKINVDCx11_ASAP7_75t_R g1036 ( .A(n_915), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_879), .Y(n_1037) );
AO31x2_ASAP7_75t_L g1038 ( .A1(n_943), .A2(n_150), .A3(n_151), .B(n_152), .Y(n_1038) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_920), .B(n_150), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_872), .B(n_151), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_835), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_1041) );
AOI221xp5_ASAP7_75t_L g1042 ( .A1(n_952), .A2(n_154), .B1(n_155), .B2(n_156), .C(n_157), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_947), .B(n_156), .Y(n_1043) );
AO21x2_ASAP7_75t_L g1044 ( .A1(n_873), .A2(n_157), .B(n_158), .Y(n_1044) );
INVx1_ASAP7_75t_SL g1045 ( .A(n_976), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_938), .Y(n_1046) );
AO21x2_ASAP7_75t_L g1047 ( .A1(n_863), .A2(n_158), .B(n_159), .Y(n_1047) );
INVxp67_ASAP7_75t_L g1048 ( .A(n_845), .Y(n_1048) );
OAI21x1_ASAP7_75t_L g1049 ( .A1(n_959), .A2(n_159), .B(n_161), .Y(n_1049) );
INVxp67_ASAP7_75t_L g1050 ( .A(n_845), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_955), .Y(n_1051) );
A2O1A1Ixp33_ASAP7_75t_L g1052 ( .A1(n_949), .A2(n_161), .B(n_162), .C(n_163), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_951), .B(n_162), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_864), .A2(n_163), .B1(n_164), .B2(n_165), .Y(n_1054) );
OA21x2_ASAP7_75t_L g1055 ( .A1(n_930), .A2(n_164), .B(n_165), .Y(n_1055) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_960), .Y(n_1056) );
AO31x2_ASAP7_75t_L g1057 ( .A1(n_836), .A2(n_166), .A3(n_167), .B(n_168), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_965), .B(n_167), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g1059 ( .A1(n_900), .A2(n_168), .B1(n_169), .B2(n_170), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_912), .B(n_169), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_913), .B(n_171), .Y(n_1061) );
INVx2_ASAP7_75t_L g1062 ( .A(n_918), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_883), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_954), .B(n_171), .Y(n_1064) );
OAI21x1_ASAP7_75t_L g1065 ( .A1(n_963), .A2(n_172), .B(n_173), .Y(n_1065) );
INVx3_ASAP7_75t_L g1066 ( .A(n_987), .Y(n_1066) );
AOI21xp5_ASAP7_75t_L g1067 ( .A1(n_844), .A2(n_174), .B(n_175), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_970), .B(n_175), .Y(n_1068) );
OA21x2_ASAP7_75t_L g1069 ( .A1(n_832), .A2(n_176), .B(n_891), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_917), .Y(n_1070) );
BUFx2_ASAP7_75t_SL g1071 ( .A(n_929), .Y(n_1071) );
A2O1A1Ixp33_ASAP7_75t_L g1072 ( .A1(n_923), .A2(n_176), .B(n_926), .C(n_933), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_833), .A2(n_902), .B1(n_986), .B2(n_897), .Y(n_1073) );
OAI22xp33_ASAP7_75t_L g1074 ( .A1(n_888), .A2(n_843), .B1(n_869), .B2(n_972), .Y(n_1074) );
AOI21xp33_ASAP7_75t_SL g1075 ( .A1(n_962), .A2(n_928), .B(n_969), .Y(n_1075) );
OAI21xp33_ASAP7_75t_L g1076 ( .A1(n_945), .A2(n_874), .B(n_866), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_927), .Y(n_1077) );
AOI21xp33_ASAP7_75t_L g1078 ( .A1(n_832), .A2(n_891), .B(n_974), .Y(n_1078) );
BUFx2_ASAP7_75t_L g1079 ( .A(n_853), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_882), .B(n_884), .Y(n_1080) );
BUFx12f_ASAP7_75t_L g1081 ( .A(n_855), .Y(n_1081) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_946), .A2(n_895), .B1(n_853), .B2(n_910), .Y(n_1082) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_878), .A2(n_871), .B1(n_898), .B2(n_870), .C(n_860), .Y(n_1083) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_924), .A2(n_907), .B1(n_948), .B2(n_921), .Y(n_1084) );
NAND2x1p5_ASAP7_75t_L g1085 ( .A(n_987), .B(n_975), .Y(n_1085) );
INVx4_ASAP7_75t_L g1086 ( .A(n_977), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_914), .Y(n_1087) );
AO31x2_ASAP7_75t_L g1088 ( .A1(n_877), .A2(n_953), .A3(n_940), .B(n_909), .Y(n_1088) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_899), .Y(n_1089) );
NOR2x1_ASAP7_75t_R g1090 ( .A(n_851), .B(n_855), .Y(n_1090) );
AOI21xp5_ASAP7_75t_L g1091 ( .A1(n_847), .A2(n_941), .B(n_919), .Y(n_1091) );
NAND2xp5_ASAP7_75t_L g1092 ( .A(n_968), .B(n_892), .Y(n_1092) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_967), .A2(n_973), .B1(n_946), .B2(n_935), .C(n_922), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_892), .B(n_885), .Y(n_1094) );
OAI21xp5_ASAP7_75t_L g1095 ( .A1(n_916), .A2(n_934), .B(n_880), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_885), .B(n_860), .Y(n_1096) );
INVx6_ASAP7_75t_SL g1097 ( .A(n_956), .Y(n_1097) );
OA21x2_ASAP7_75t_L g1098 ( .A1(n_932), .A2(n_966), .B(n_979), .Y(n_1098) );
AOI21xp5_ASAP7_75t_L g1099 ( .A1(n_982), .A2(n_964), .B(n_971), .Y(n_1099) );
BUFx3_ASAP7_75t_L g1100 ( .A(n_894), .Y(n_1100) );
NAND2xp5_ASAP7_75t_L g1101 ( .A(n_894), .B(n_937), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_894), .B(n_937), .Y(n_1102) );
NAND2xp5_ASAP7_75t_SL g1103 ( .A(n_982), .B(n_980), .Y(n_1103) );
AO31x2_ASAP7_75t_L g1104 ( .A1(n_978), .A2(n_903), .A3(n_956), .B(n_927), .Y(n_1104) );
CKINVDCx16_ASAP7_75t_R g1105 ( .A(n_893), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_906), .B(n_925), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_893), .B(n_911), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_937), .B(n_981), .Y(n_1108) );
OA21x2_ASAP7_75t_L g1109 ( .A1(n_903), .A2(n_981), .B(n_911), .Y(n_1109) );
OR2x2_ASAP7_75t_L g1110 ( .A(n_989), .B(n_622), .Y(n_1110) );
INVx2_ASAP7_75t_L g1111 ( .A(n_841), .Y(n_1111) );
AOI21xp5_ASAP7_75t_L g1112 ( .A1(n_837), .A2(n_678), .B(n_838), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_834), .B(n_634), .Y(n_1113) );
BUFx3_ASAP7_75t_L g1114 ( .A(n_859), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_989), .B(n_889), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_852), .Y(n_1116) );
OAI21xp5_ASAP7_75t_L g1117 ( .A1(n_837), .A2(n_772), .B(n_786), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_989), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_834), .B(n_634), .Y(n_1119) );
NOR2xp67_ASAP7_75t_L g1120 ( .A(n_862), .B(n_984), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g1121 ( .A(n_989), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_834), .B(n_634), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_989), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_841), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_887), .A2(n_755), .B1(n_627), .B2(n_769), .Y(n_1125) );
NOR2x1_ASAP7_75t_SL g1126 ( .A(n_960), .B(n_758), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g1127 ( .A1(n_887), .A2(n_728), .B1(n_587), .B2(n_740), .Y(n_1127) );
AOI21x1_ASAP7_75t_L g1128 ( .A1(n_868), .A2(n_957), .B(n_708), .Y(n_1128) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_983), .A2(n_740), .B1(n_717), .B2(n_718), .Y(n_1129) );
A2O1A1Ixp33_ASAP7_75t_L g1130 ( .A1(n_887), .A2(n_634), .B(n_942), .C(n_901), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_989), .B(n_622), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_984), .Y(n_1132) );
AO31x2_ASAP7_75t_L g1133 ( .A1(n_908), .A2(n_856), .A3(n_842), .B(n_837), .Y(n_1133) );
CKINVDCx5p33_ASAP7_75t_R g1134 ( .A(n_859), .Y(n_1134) );
NAND2x1_ASAP7_75t_L g1135 ( .A(n_960), .B(n_849), .Y(n_1135) );
INVx6_ASAP7_75t_L g1136 ( .A(n_984), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_841), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_837), .A2(n_678), .B(n_838), .Y(n_1138) );
AOI21xp5_ASAP7_75t_L g1139 ( .A1(n_837), .A2(n_678), .B(n_838), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_834), .B(n_634), .Y(n_1140) );
AO31x2_ASAP7_75t_L g1141 ( .A1(n_908), .A2(n_856), .A3(n_842), .B(n_837), .Y(n_1141) );
OAI22xp33_ASAP7_75t_L g1142 ( .A1(n_983), .A2(n_740), .B1(n_717), .B2(n_718), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_993), .B(n_1079), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1144 ( .A(n_1127), .B(n_1129), .Y(n_1144) );
OA21x2_ASAP7_75t_L g1145 ( .A1(n_1094), .A2(n_1102), .B(n_1101), .Y(n_1145) );
OAI221xp5_ASAP7_75t_L g1146 ( .A1(n_1125), .A2(n_1073), .B1(n_999), .B2(n_1083), .C(n_1130), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1012), .Y(n_1147) );
OA21x2_ASAP7_75t_L g1148 ( .A1(n_1094), .A2(n_1102), .B(n_1101), .Y(n_1148) );
AO21x2_ASAP7_75t_L g1149 ( .A1(n_1078), .A2(n_1128), .B(n_1096), .Y(n_1149) );
AND2x4_ASAP7_75t_L g1150 ( .A(n_993), .B(n_1009), .Y(n_1150) );
AO21x2_ASAP7_75t_L g1151 ( .A1(n_1078), .A2(n_1096), .B(n_1051), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1142), .B(n_1110), .Y(n_1152) );
NOR2xp33_ASAP7_75t_L g1153 ( .A(n_1131), .B(n_1113), .Y(n_1153) );
OR2x6_ASAP7_75t_L g1154 ( .A(n_1001), .B(n_1017), .Y(n_1154) );
INVx1_ASAP7_75t_L g1155 ( .A(n_994), .Y(n_1155) );
HB1xp67_ASAP7_75t_L g1156 ( .A(n_995), .Y(n_1156) );
AO21x2_ASAP7_75t_L g1157 ( .A1(n_1077), .A2(n_1091), .B(n_1092), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1115), .B(n_996), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g1159 ( .A(n_1118), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_998), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1007), .Y(n_1161) );
BUFx3_ASAP7_75t_L g1162 ( .A(n_1056), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_991), .B(n_1000), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1116), .B(n_1113), .Y(n_1164) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1136), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1025), .B(n_1062), .Y(n_1166) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1014), .Y(n_1167) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1015), .Y(n_1168) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1097), .Y(n_1169) );
AND2x4_ASAP7_75t_L g1170 ( .A(n_1020), .B(n_1029), .Y(n_1170) );
OR2x6_ASAP7_75t_L g1171 ( .A(n_1001), .B(n_1017), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_997), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g1173 ( .A1(n_1075), .A2(n_1030), .B1(n_1046), .B2(n_1083), .C(n_1003), .Y(n_1173) );
OAI21xp5_ASAP7_75t_L g1174 ( .A1(n_1072), .A2(n_1084), .B(n_1013), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1004), .B(n_1121), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_1123), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1111), .B(n_1124), .Y(n_1177) );
INVx2_ASAP7_75t_SL g1178 ( .A(n_1136), .Y(n_1178) );
INVx4_ASAP7_75t_L g1179 ( .A(n_1085), .Y(n_1179) );
INVx2_ASAP7_75t_SL g1180 ( .A(n_1135), .Y(n_1180) );
INVx2_ASAP7_75t_L g1181 ( .A(n_1137), .Y(n_1181) );
OAI222xp33_ASAP7_75t_L g1182 ( .A1(n_1003), .A2(n_1063), .B1(n_1037), .B2(n_1019), .C1(n_1005), .C2(n_1050), .Y(n_1182) );
OR2x6_ASAP7_75t_L g1183 ( .A(n_1048), .B(n_1022), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1184 ( .A(n_1004), .B(n_1010), .Y(n_1184) );
AOI221xp5_ASAP7_75t_L g1185 ( .A1(n_1070), .A2(n_1074), .B1(n_1042), .B2(n_1084), .C(n_1054), .Y(n_1185) );
CKINVDCx20_ASAP7_75t_R g1186 ( .A(n_1134), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1119), .B(n_1122), .Y(n_1187) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_1006), .A2(n_1042), .B1(n_1022), .B2(n_1076), .Y(n_1188) );
INVx3_ASAP7_75t_L g1189 ( .A(n_1097), .Y(n_1189) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_1045), .B(n_1043), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_997), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1006), .B(n_1107), .Y(n_1192) );
OAI222xp33_ASAP7_75t_L g1193 ( .A1(n_1082), .A2(n_1105), .B1(n_1059), .B2(n_1054), .C1(n_1027), .C2(n_1016), .Y(n_1193) );
BUFx3_ASAP7_75t_L g1194 ( .A(n_1021), .Y(n_1194) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_1041), .B(n_1052), .C(n_1023), .Y(n_1195) );
HB1xp67_ASAP7_75t_L g1196 ( .A(n_1089), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1119), .B(n_1122), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_1018), .A2(n_1013), .B1(n_1140), .B2(n_1053), .Y(n_1198) );
OAI211xp5_ASAP7_75t_L g1199 ( .A1(n_1008), .A2(n_1064), .B(n_1032), .C(n_1039), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1045), .B(n_1058), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1058), .Y(n_1201) );
OA21x2_ASAP7_75t_L g1202 ( .A1(n_1108), .A2(n_1049), .B(n_1065), .Y(n_1202) );
INVx4_ASAP7_75t_L g1203 ( .A(n_1066), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_1032), .A2(n_1039), .B1(n_1100), .B2(n_1053), .Y(n_1204) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1068), .B(n_1080), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1206 ( .A(n_1068), .B(n_1024), .Y(n_1206) );
OA21x2_ASAP7_75t_L g1207 ( .A1(n_1095), .A2(n_1040), .B(n_1099), .Y(n_1207) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1026), .B(n_1028), .Y(n_1208) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1026), .B(n_1028), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1060), .Y(n_1210) );
AO21x2_ASAP7_75t_L g1211 ( .A1(n_1035), .A2(n_1044), .B(n_1040), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1140), .B(n_1090), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1060), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1057), .B(n_1061), .Y(n_1214) );
AOI21xp5_ASAP7_75t_SL g1215 ( .A1(n_1055), .A2(n_1093), .B(n_1069), .Y(n_1215) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1034), .Y(n_1216) );
INVx4_ASAP7_75t_SL g1217 ( .A(n_1038), .Y(n_1217) );
OAI21xp5_ASAP7_75t_L g1218 ( .A1(n_1117), .A2(n_1067), .B(n_1138), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1061), .Y(n_1219) );
INVx3_ASAP7_75t_L g1220 ( .A(n_1086), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1057), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1038), .B(n_1086), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1069), .B(n_1038), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1126), .Y(n_1224) );
OA21x2_ASAP7_75t_L g1225 ( .A1(n_1095), .A2(n_1117), .B(n_1106), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1109), .B(n_1087), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1031), .Y(n_1227) );
AOI21xp5_ASAP7_75t_L g1228 ( .A1(n_1103), .A2(n_1112), .B(n_1139), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1033), .B(n_990), .Y(n_1229) );
INVx2_ASAP7_75t_SL g1230 ( .A(n_1132), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_1055), .A2(n_1081), .B1(n_1047), .B2(n_1035), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1120), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_990), .B(n_1047), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_990), .B(n_1044), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1114), .B(n_1071), .Y(n_1235) );
CKINVDCx5p33_ASAP7_75t_R g1236 ( .A(n_1036), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1109), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1088), .B(n_1104), .Y(n_1238) );
OR2x2_ASAP7_75t_L g1239 ( .A(n_1088), .B(n_1104), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1088), .B(n_1141), .Y(n_1240) );
OAI21xp5_ASAP7_75t_L g1241 ( .A1(n_992), .A2(n_1002), .B(n_1011), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_1098), .A2(n_740), .B1(n_717), .B2(n_718), .Y(n_1242) );
AND2x4_ASAP7_75t_L g1243 ( .A(n_1133), .B(n_1141), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1133), .B(n_989), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_994), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1246 ( .A1(n_1127), .A2(n_740), .B1(n_717), .B2(n_718), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_991), .B(n_1000), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_991), .B(n_1000), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1127), .B(n_889), .Y(n_1249) );
OA21x2_ASAP7_75t_L g1250 ( .A1(n_1094), .A2(n_1102), .B(n_1101), .Y(n_1250) );
INVx3_ASAP7_75t_L g1251 ( .A(n_1097), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_994), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1012), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1127), .B(n_889), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_991), .B(n_1000), .Y(n_1255) );
BUFx4f_ASAP7_75t_SL g1256 ( .A(n_1021), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1009), .B(n_1004), .Y(n_1257) );
INVx1_ASAP7_75t_L g1258 ( .A(n_994), .Y(n_1258) );
INVx1_ASAP7_75t_L g1259 ( .A(n_994), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1214), .B(n_1229), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1257), .B(n_1226), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1262 ( .A(n_1153), .B(n_1152), .Y(n_1262) );
AND2x4_ASAP7_75t_SL g1263 ( .A(n_1154), .B(n_1171), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1221), .Y(n_1264) );
INVx3_ASAP7_75t_L g1265 ( .A(n_1220), .Y(n_1265) );
HB1xp67_ASAP7_75t_L g1266 ( .A(n_1162), .Y(n_1266) );
BUFx3_ASAP7_75t_L g1267 ( .A(n_1162), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1214), .B(n_1229), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1234), .B(n_1147), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1234), .B(n_1147), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1257), .B(n_1226), .Y(n_1271) );
INVxp67_ASAP7_75t_L g1272 ( .A(n_1184), .Y(n_1272) );
INVxp67_ASAP7_75t_L g1273 ( .A(n_1230), .Y(n_1273) );
HB1xp67_ASAP7_75t_L g1274 ( .A(n_1154), .Y(n_1274) );
BUFx3_ASAP7_75t_L g1275 ( .A(n_1143), .Y(n_1275) );
INVxp33_ASAP7_75t_L g1276 ( .A(n_1196), .Y(n_1276) );
BUFx2_ASAP7_75t_L g1277 ( .A(n_1154), .Y(n_1277) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1237), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_1154), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1145), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1145), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1145), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1253), .B(n_1222), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1253), .B(n_1222), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1148), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1148), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1163), .B(n_1166), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1153), .B(n_1192), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1163), .B(n_1166), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1177), .B(n_1247), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1192), .B(n_1164), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1148), .Y(n_1292) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_1171), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1250), .Y(n_1294) );
INVx1_ASAP7_75t_SL g1295 ( .A(n_1165), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g1296 ( .A(n_1156), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1177), .B(n_1247), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1155), .Y(n_1298) );
AND2x4_ASAP7_75t_L g1299 ( .A(n_1171), .B(n_1220), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1160), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1161), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1167), .Y(n_1302) );
INVx4_ASAP7_75t_L g1303 ( .A(n_1171), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1245), .Y(n_1304) );
HB1xp67_ASAP7_75t_L g1305 ( .A(n_1175), .Y(n_1305) );
INVx3_ASAP7_75t_L g1306 ( .A(n_1203), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1248), .B(n_1255), .Y(n_1307) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1158), .B(n_1159), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1244), .B(n_1176), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1144), .B(n_1200), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1173), .B(n_1252), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g1312 ( .A(n_1198), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_1212), .B(n_1235), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1258), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1223), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1259), .B(n_1185), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1223), .Y(n_1317) );
HB1xp67_ASAP7_75t_L g1318 ( .A(n_1143), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1205), .B(n_1206), .Y(n_1319) );
BUFx2_ASAP7_75t_L g1320 ( .A(n_1143), .Y(n_1320) );
AOI221xp5_ASAP7_75t_L g1321 ( .A1(n_1246), .A2(n_1146), .B1(n_1242), .B2(n_1182), .C(n_1193), .Y(n_1321) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1249), .B(n_1254), .Y(n_1322) );
INVx3_ASAP7_75t_L g1323 ( .A(n_1203), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1217), .Y(n_1324) );
BUFx2_ASAP7_75t_L g1325 ( .A(n_1203), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1233), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1248), .B(n_1255), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1328 ( .A(n_1181), .B(n_1225), .Y(n_1328) );
BUFx2_ASAP7_75t_L g1329 ( .A(n_1183), .Y(n_1329) );
INVx4_ASAP7_75t_L g1330 ( .A(n_1179), .Y(n_1330) );
NOR2xp33_ASAP7_75t_L g1331 ( .A(n_1276), .B(n_1186), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1264), .Y(n_1332) );
NAND2xp5_ASAP7_75t_SL g1333 ( .A(n_1330), .B(n_1224), .Y(n_1333) );
INVx2_ASAP7_75t_SL g1334 ( .A(n_1267), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1287), .B(n_1168), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1260), .B(n_1238), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1287), .B(n_1172), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1264), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1260), .B(n_1238), .Y(n_1339) );
INVx1_ASAP7_75t_SL g1340 ( .A(n_1267), .Y(n_1340) );
INVx4_ASAP7_75t_L g1341 ( .A(n_1330), .Y(n_1341) );
HB1xp67_ASAP7_75t_L g1342 ( .A(n_1266), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1343 ( .A(n_1261), .B(n_1240), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1268), .B(n_1243), .Y(n_1344) );
AND2x4_ASAP7_75t_SL g1345 ( .A(n_1303), .B(n_1179), .Y(n_1345) );
AND2x4_ASAP7_75t_L g1346 ( .A(n_1324), .B(n_1243), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1268), .B(n_1243), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1289), .B(n_1191), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1349 ( .A(n_1261), .B(n_1151), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1283), .B(n_1225), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1283), .B(n_1225), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1289), .B(n_1201), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1290), .B(n_1227), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1290), .B(n_1219), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1355 ( .A(n_1284), .B(n_1149), .Y(n_1355) );
CKINVDCx20_ASAP7_75t_R g1356 ( .A(n_1295), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1325), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_1321), .A2(n_1188), .B1(n_1183), .B2(n_1195), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1297), .B(n_1213), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1297), .B(n_1210), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1284), .B(n_1149), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1271), .B(n_1239), .Y(n_1362) );
NAND2x1p5_ASAP7_75t_L g1363 ( .A(n_1330), .B(n_1179), .Y(n_1363) );
OR2x2_ASAP7_75t_L g1364 ( .A(n_1271), .B(n_1183), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1269), .B(n_1157), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1269), .B(n_1157), .Y(n_1366) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_1325), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1368 ( .A(n_1270), .B(n_1211), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1270), .B(n_1211), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1307), .B(n_1204), .Y(n_1370) );
HB1xp67_ASAP7_75t_L g1371 ( .A(n_1296), .Y(n_1371) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1278), .Y(n_1372) );
BUFx2_ASAP7_75t_SL g1373 ( .A(n_1306), .Y(n_1373) );
AND2x4_ASAP7_75t_SL g1374 ( .A(n_1303), .B(n_1183), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1307), .B(n_1204), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1309), .B(n_1190), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1326), .B(n_1207), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1327), .B(n_1150), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1379 ( .A(n_1309), .B(n_1174), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_1328), .B(n_1207), .Y(n_1380) );
NAND2x1p5_ASAP7_75t_L g1381 ( .A(n_1306), .B(n_1169), .Y(n_1381) );
OAI21xp5_ASAP7_75t_L g1382 ( .A1(n_1312), .A2(n_1188), .B(n_1199), .Y(n_1382) );
AND3x1_ASAP7_75t_L g1383 ( .A(n_1288), .B(n_1189), .C(n_1169), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1384 ( .A(n_1328), .B(n_1207), .Y(n_1384) );
NOR2xp33_ASAP7_75t_L g1385 ( .A(n_1313), .B(n_1186), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1322), .B(n_1209), .Y(n_1386) );
NAND2xp67_ASAP7_75t_L g1387 ( .A(n_1263), .B(n_1216), .Y(n_1387) );
NOR2xp33_ASAP7_75t_R g1388 ( .A(n_1306), .B(n_1256), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1327), .B(n_1202), .Y(n_1389) );
OR2x2_ASAP7_75t_L g1390 ( .A(n_1322), .B(n_1208), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1332), .Y(n_1391) );
NAND2x1_ASAP7_75t_L g1392 ( .A(n_1341), .B(n_1303), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1371), .B(n_1305), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1370), .B(n_1272), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1332), .Y(n_1395) );
OAI31xp33_ASAP7_75t_L g1396 ( .A1(n_1363), .A2(n_1263), .A3(n_1311), .B(n_1277), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1389), .B(n_1315), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1376), .Y(n_1398) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1389), .B(n_1315), .Y(n_1399) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1362), .B(n_1308), .Y(n_1400) );
AND3x2_ASAP7_75t_L g1401 ( .A(n_1385), .B(n_1277), .C(n_1293), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1375), .B(n_1308), .Y(n_1402) );
INVxp67_ASAP7_75t_L g1403 ( .A(n_1342), .Y(n_1403) );
NOR2xp33_ASAP7_75t_L g1404 ( .A(n_1356), .B(n_1165), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1376), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1386), .B(n_1298), .Y(n_1406) );
OR2x2_ASAP7_75t_L g1407 ( .A(n_1362), .B(n_1319), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1408 ( .A(n_1386), .B(n_1300), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1338), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1390), .B(n_1301), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1336), .B(n_1317), .Y(n_1411) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_1357), .Y(n_1412) );
OR2x2_ASAP7_75t_L g1413 ( .A(n_1343), .B(n_1319), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1390), .B(n_1302), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1337), .B(n_1304), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1336), .B(n_1317), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1417 ( .A(n_1343), .B(n_1280), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1348), .B(n_1314), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1339), .B(n_1280), .Y(n_1419) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1352), .B(n_1310), .Y(n_1420) );
OR2x2_ASAP7_75t_L g1421 ( .A(n_1379), .B(n_1281), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1339), .B(n_1281), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1350), .B(n_1351), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1350), .B(n_1282), .Y(n_1424) );
INVx2_ASAP7_75t_L g1425 ( .A(n_1372), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1351), .B(n_1282), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1354), .B(n_1359), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1344), .B(n_1285), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1344), .B(n_1285), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1379), .B(n_1286), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1347), .B(n_1286), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1360), .B(n_1310), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1335), .B(n_1262), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1353), .B(n_1291), .Y(n_1434) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1349), .B(n_1292), .Y(n_1435) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1331), .B(n_1178), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1347), .B(n_1292), .Y(n_1437) );
INVx1_ASAP7_75t_SL g1438 ( .A(n_1340), .Y(n_1438) );
INVx1_ASAP7_75t_SL g1439 ( .A(n_1340), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1355), .B(n_1294), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1423), .B(n_1355), .Y(n_1441) );
OR2x2_ASAP7_75t_L g1442 ( .A(n_1423), .B(n_1349), .Y(n_1442) );
NOR2xp67_ASAP7_75t_L g1443 ( .A(n_1403), .B(n_1341), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1400), .B(n_1368), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1435), .Y(n_1445) );
OAI32xp33_ASAP7_75t_L g1446 ( .A1(n_1438), .A2(n_1341), .A3(n_1363), .B1(n_1367), .B2(n_1381), .Y(n_1446) );
HB1xp67_ASAP7_75t_L g1447 ( .A(n_1412), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1448 ( .A(n_1400), .B(n_1368), .Y(n_1448) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_1411), .B(n_1361), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1407), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1407), .Y(n_1451) );
OR2x2_ASAP7_75t_L g1452 ( .A(n_1413), .B(n_1369), .Y(n_1452) );
INVx1_ASAP7_75t_L g1453 ( .A(n_1435), .Y(n_1453) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_1402), .A2(n_1383), .B1(n_1358), .B2(n_1382), .Y(n_1454) );
INVxp67_ASAP7_75t_L g1455 ( .A(n_1439), .Y(n_1455) );
INVx2_ASAP7_75t_L g1456 ( .A(n_1425), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1411), .B(n_1361), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1413), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1397), .B(n_1369), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1416), .B(n_1382), .Y(n_1460) );
OR2x2_ASAP7_75t_L g1461 ( .A(n_1421), .B(n_1365), .Y(n_1461) );
HB1xp67_ASAP7_75t_L g1462 ( .A(n_1424), .Y(n_1462) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1425), .Y(n_1463) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1391), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1416), .B(n_1365), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1391), .Y(n_1466) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1397), .B(n_1366), .Y(n_1467) );
INVx1_ASAP7_75t_L g1468 ( .A(n_1395), .Y(n_1468) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1395), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1440), .B(n_1366), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1399), .B(n_1380), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1440), .B(n_1377), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1409), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1399), .B(n_1380), .Y(n_1474) );
INVxp67_ASAP7_75t_SL g1475 ( .A(n_1393), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1424), .B(n_1384), .Y(n_1476) );
AOI21xp33_ASAP7_75t_SL g1477 ( .A1(n_1396), .A2(n_1363), .B(n_1236), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1419), .B(n_1377), .Y(n_1478) );
AOI22xp5_ASAP7_75t_L g1479 ( .A1(n_1398), .A2(n_1383), .B1(n_1341), .B2(n_1346), .Y(n_1479) );
NOR2xp33_ASAP7_75t_L g1480 ( .A(n_1404), .B(n_1169), .Y(n_1480) );
NOR2x1_ASAP7_75t_L g1481 ( .A(n_1443), .B(n_1392), .Y(n_1481) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_1479), .A2(n_1392), .B1(n_1373), .B2(n_1427), .Y(n_1482) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1462), .Y(n_1483) );
AOI21xp5_ASAP7_75t_L g1484 ( .A1(n_1446), .A2(n_1333), .B(n_1334), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1485 ( .A(n_1460), .B(n_1419), .Y(n_1485) );
O2A1O1Ixp33_ASAP7_75t_SL g1486 ( .A1(n_1477), .A2(n_1387), .B(n_1334), .C(n_1406), .Y(n_1486) );
AOI211xp5_ASAP7_75t_L g1487 ( .A1(n_1446), .A2(n_1388), .B(n_1436), .C(n_1430), .Y(n_1487) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1445), .Y(n_1488) );
INVx1_ASAP7_75t_SL g1489 ( .A(n_1447), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1445), .Y(n_1490) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1453), .Y(n_1491) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1453), .B(n_1422), .Y(n_1492) );
AOI221xp5_ASAP7_75t_L g1493 ( .A1(n_1475), .A2(n_1394), .B1(n_1405), .B2(n_1433), .C(n_1432), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1494 ( .A(n_1467), .B(n_1422), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1464), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1441), .B(n_1426), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1464), .Y(n_1497) );
AOI211xp5_ASAP7_75t_L g1498 ( .A1(n_1454), .A2(n_1421), .B(n_1430), .C(n_1417), .Y(n_1498) );
AOI21xp33_ASAP7_75t_L g1499 ( .A1(n_1480), .A2(n_1232), .B(n_1273), .Y(n_1499) );
AOI332xp33_ASAP7_75t_L g1500 ( .A1(n_1450), .A2(n_1434), .A3(n_1420), .B1(n_1408), .B2(n_1410), .B3(n_1414), .C1(n_1415), .C2(n_1418), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1441), .B(n_1426), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1466), .Y(n_1502) );
NAND2xp5_ASAP7_75t_L g1503 ( .A(n_1467), .B(n_1428), .Y(n_1503) );
HB1xp67_ASAP7_75t_L g1504 ( .A(n_1442), .Y(n_1504) );
OAI21xp33_ASAP7_75t_L g1505 ( .A1(n_1442), .A2(n_1437), .B(n_1429), .Y(n_1505) );
INVx2_ASAP7_75t_L g1506 ( .A(n_1456), .Y(n_1506) );
OAI22xp33_ASAP7_75t_L g1507 ( .A1(n_1452), .A2(n_1293), .B1(n_1381), .B2(n_1320), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1508 ( .A(n_1452), .B(n_1417), .Y(n_1508) );
INVxp67_ASAP7_75t_L g1509 ( .A(n_1489), .Y(n_1509) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1508), .Y(n_1510) );
AOI211xp5_ASAP7_75t_L g1511 ( .A1(n_1486), .A2(n_1455), .B(n_1236), .C(n_1458), .Y(n_1511) );
A2O1A1Ixp33_ASAP7_75t_L g1512 ( .A1(n_1500), .A2(n_1345), .B(n_1476), .C(n_1444), .Y(n_1512) );
INVxp67_ASAP7_75t_SL g1513 ( .A(n_1481), .Y(n_1513) );
AOI221xp5_ASAP7_75t_L g1514 ( .A1(n_1498), .A2(n_1451), .B1(n_1470), .B2(n_1459), .C(n_1457), .Y(n_1514) );
AOI21xp33_ASAP7_75t_L g1515 ( .A1(n_1487), .A2(n_1178), .B(n_1230), .Y(n_1515) );
OAI211xp5_ASAP7_75t_L g1516 ( .A1(n_1486), .A2(n_1279), .B(n_1274), .C(n_1194), .Y(n_1516) );
NAND2xp5_ASAP7_75t_L g1517 ( .A(n_1493), .B(n_1459), .Y(n_1517) );
NOR3xp33_ASAP7_75t_L g1518 ( .A(n_1499), .B(n_1194), .C(n_1189), .Y(n_1518) );
AOI222xp33_ASAP7_75t_L g1519 ( .A1(n_1504), .A2(n_1316), .B1(n_1476), .B2(n_1474), .C1(n_1471), .C2(n_1437), .Y(n_1519) );
AOI21xp5_ASAP7_75t_L g1520 ( .A1(n_1484), .A2(n_1478), .B(n_1472), .Y(n_1520) );
AOI22xp5_ASAP7_75t_L g1521 ( .A1(n_1505), .A2(n_1431), .B1(n_1429), .B2(n_1428), .Y(n_1521) );
OAI221xp5_ASAP7_75t_L g1522 ( .A1(n_1482), .A2(n_1448), .B1(n_1444), .B2(n_1461), .C(n_1449), .Y(n_1522) );
A2O1A1Ixp33_ASAP7_75t_L g1523 ( .A1(n_1508), .A2(n_1345), .B(n_1448), .C(n_1461), .Y(n_1523) );
OAI221xp5_ASAP7_75t_L g1524 ( .A1(n_1483), .A2(n_1465), .B1(n_1381), .B2(n_1469), .C(n_1468), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1525 ( .A(n_1496), .B(n_1471), .Y(n_1525) );
AOI22xp5_ASAP7_75t_L g1526 ( .A1(n_1507), .A2(n_1431), .B1(n_1474), .B2(n_1346), .Y(n_1526) );
AOI22xp5_ASAP7_75t_L g1527 ( .A1(n_1485), .A2(n_1346), .B1(n_1329), .B2(n_1466), .Y(n_1527) );
NOR2xp33_ASAP7_75t_L g1528 ( .A(n_1494), .B(n_1256), .Y(n_1528) );
NOR3xp33_ASAP7_75t_L g1529 ( .A(n_1516), .B(n_1189), .C(n_1251), .Y(n_1529) );
AOI22xp5_ASAP7_75t_L g1530 ( .A1(n_1514), .A2(n_1491), .B1(n_1488), .B2(n_1490), .Y(n_1530) );
OAI222xp33_ASAP7_75t_L g1531 ( .A1(n_1513), .A2(n_1492), .B1(n_1503), .B2(n_1501), .C1(n_1496), .C2(n_1497), .Y(n_1531) );
HB1xp67_ASAP7_75t_L g1532 ( .A(n_1509), .Y(n_1532) );
OAI211xp5_ASAP7_75t_L g1533 ( .A1(n_1511), .A2(n_1251), .B(n_1231), .C(n_1329), .Y(n_1533) );
OAI21xp33_ASAP7_75t_L g1534 ( .A1(n_1512), .A2(n_1502), .B(n_1497), .Y(n_1534) );
INVx2_ASAP7_75t_SL g1535 ( .A(n_1510), .Y(n_1535) );
AOI211x1_ASAP7_75t_SL g1536 ( .A1(n_1515), .A2(n_1506), .B(n_1463), .C(n_1456), .Y(n_1536) );
AOI211xp5_ASAP7_75t_L g1537 ( .A1(n_1518), .A2(n_1251), .B(n_1299), .C(n_1501), .Y(n_1537) );
NOR2xp33_ASAP7_75t_R g1538 ( .A(n_1528), .B(n_1401), .Y(n_1538) );
NAND3xp33_ASAP7_75t_L g1539 ( .A(n_1518), .B(n_1502), .C(n_1495), .Y(n_1539) );
OAI221xp5_ASAP7_75t_L g1540 ( .A1(n_1522), .A2(n_1495), .B1(n_1506), .B2(n_1473), .C(n_1373), .Y(n_1540) );
NOR2xp67_ASAP7_75t_L g1541 ( .A(n_1526), .B(n_1463), .Y(n_1541) );
NAND4xp25_ASAP7_75t_L g1542 ( .A(n_1519), .B(n_1299), .C(n_1231), .D(n_1275), .Y(n_1542) );
NAND2xp5_ASAP7_75t_L g1543 ( .A(n_1532), .B(n_1517), .Y(n_1543) );
OAI221xp5_ASAP7_75t_L g1544 ( .A1(n_1537), .A2(n_1523), .B1(n_1524), .B2(n_1520), .C(n_1527), .Y(n_1544) );
OR2x6_ASAP7_75t_L g1545 ( .A(n_1535), .B(n_1533), .Y(n_1545) );
NAND2xp5_ASAP7_75t_SL g1546 ( .A(n_1538), .B(n_1521), .Y(n_1546) );
AOI211xp5_ASAP7_75t_L g1547 ( .A1(n_1529), .A2(n_1299), .B(n_1525), .C(n_1215), .Y(n_1547) );
OAI211xp5_ASAP7_75t_L g1548 ( .A1(n_1534), .A2(n_1318), .B(n_1218), .C(n_1215), .Y(n_1548) );
NOR2x1_ASAP7_75t_L g1549 ( .A(n_1531), .B(n_1539), .Y(n_1549) );
NOR3xp33_ASAP7_75t_L g1550 ( .A(n_1531), .B(n_1265), .C(n_1323), .Y(n_1550) );
NAND4xp25_ASAP7_75t_L g1551 ( .A(n_1536), .B(n_1275), .C(n_1320), .D(n_1364), .Y(n_1551) );
NAND2xp5_ASAP7_75t_SL g1552 ( .A(n_1541), .B(n_1323), .Y(n_1552) );
INVx1_ASAP7_75t_SL g1553 ( .A(n_1543), .Y(n_1553) );
AND4x1_ASAP7_75t_L g1554 ( .A(n_1547), .B(n_1530), .C(n_1540), .D(n_1542), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1549), .B(n_1473), .Y(n_1555) );
NOR3xp33_ASAP7_75t_L g1556 ( .A(n_1546), .B(n_1180), .C(n_1323), .Y(n_1556) );
NAND3xp33_ASAP7_75t_SL g1557 ( .A(n_1548), .B(n_1241), .C(n_1228), .Y(n_1557) );
BUFx2_ASAP7_75t_L g1558 ( .A(n_1545), .Y(n_1558) );
NOR3xp33_ASAP7_75t_L g1559 ( .A(n_1544), .B(n_1180), .C(n_1265), .Y(n_1559) );
INVx2_ASAP7_75t_SL g1560 ( .A(n_1558), .Y(n_1560) );
INVx3_ASAP7_75t_L g1561 ( .A(n_1554), .Y(n_1561) );
INVx2_ASAP7_75t_L g1562 ( .A(n_1553), .Y(n_1562) );
BUFx2_ASAP7_75t_L g1563 ( .A(n_1555), .Y(n_1563) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1556), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1559), .Y(n_1565) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1560), .Y(n_1566) );
INVx2_ASAP7_75t_L g1567 ( .A(n_1560), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1562), .Y(n_1568) );
INVx1_ASAP7_75t_L g1569 ( .A(n_1562), .Y(n_1569) );
OAI22x1_ASAP7_75t_L g1570 ( .A1(n_1561), .A2(n_1552), .B1(n_1545), .B2(n_1557), .Y(n_1570) );
CKINVDCx20_ASAP7_75t_R g1571 ( .A(n_1566), .Y(n_1571) );
OAI22xp5_ASAP7_75t_L g1572 ( .A1(n_1567), .A2(n_1561), .B1(n_1562), .B2(n_1564), .Y(n_1572) );
AOI211xp5_ASAP7_75t_L g1573 ( .A1(n_1568), .A2(n_1561), .B(n_1565), .C(n_1564), .Y(n_1573) );
XOR2xp5_ASAP7_75t_L g1574 ( .A(n_1571), .B(n_1569), .Y(n_1574) );
AOI222xp33_ASAP7_75t_SL g1575 ( .A1(n_1572), .A2(n_1565), .B1(n_1563), .B2(n_1570), .C1(n_1550), .C2(n_1551), .Y(n_1575) );
AOI222xp33_ASAP7_75t_L g1576 ( .A1(n_1573), .A2(n_1563), .B1(n_1170), .B2(n_1187), .C1(n_1197), .C2(n_1345), .Y(n_1576) );
INVx2_ASAP7_75t_L g1577 ( .A(n_1574), .Y(n_1577) );
OA21x2_ASAP7_75t_L g1578 ( .A1(n_1575), .A2(n_1170), .B(n_1378), .Y(n_1578) );
OAI21xp33_ASAP7_75t_L g1579 ( .A1(n_1577), .A2(n_1576), .B(n_1387), .Y(n_1579) );
AOI22xp5_ASAP7_75t_L g1580 ( .A1(n_1579), .A2(n_1578), .B1(n_1346), .B2(n_1374), .Y(n_1580) );
endmodule