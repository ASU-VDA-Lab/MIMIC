module fake_jpeg_25499_n_107 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_52),
.Y(n_55)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_43),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_36),
.B1(n_43),
.B2(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_18),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_59),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_61),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_40),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_5),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_62)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_20),
.B1(n_32),
.B2(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_51),
.B(n_1),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_6),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_63),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_76),
.B(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_2),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_73),
.A2(n_77),
.B(n_80),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_6),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_79),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_11),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_15),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_75),
.C(n_73),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_96),
.B1(n_89),
.B2(n_88),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_74),
.B1(n_69),
.B2(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_89),
.B1(n_84),
.B2(n_83),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_86),
.B(n_87),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_92),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_99),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_84),
.C(n_24),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_25),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_26),
.C(n_27),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_28),
.Y(n_107)
);


endmodule