module fake_jpeg_1190_n_187 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_13),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_13),
.B(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_15),
.A2(n_3),
.B(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_4),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_56),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_50),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_56),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_23),
.A2(n_4),
.B(n_6),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_18),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_78),
.B1(n_74),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_26),
.B1(n_27),
.B2(n_20),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_80),
.B1(n_54),
.B2(n_63),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_32),
.A2(n_26),
.B1(n_24),
.B2(n_20),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_61),
.B1(n_71),
.B2(n_73),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_30),
.A2(n_26),
.B1(n_24),
.B2(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_35),
.B(n_27),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_75),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_68),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_22),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g71 ( 
.A1(n_33),
.A2(n_19),
.B1(n_21),
.B2(n_8),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_21),
.B1(n_7),
.B2(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_6),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_31),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_9),
.B1(n_10),
.B2(n_42),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_10),
.B1(n_46),
.B2(n_23),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_89),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_92),
.B(n_107),
.Y(n_132)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_110),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_83),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_100),
.A2(n_73),
.B1(n_67),
.B2(n_71),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_83),
.B(n_82),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_113),
.B(n_71),
.Y(n_123)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_83),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_73),
.C(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_85),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_69),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_90),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_130),
.B1(n_131),
.B2(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_71),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_127),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_111),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_128),
.C(n_129),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_97),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_84),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_87),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_87),
.B1(n_60),
.B2(n_64),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_60),
.B1(n_64),
.B2(n_72),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_91),
.A2(n_70),
.B1(n_72),
.B2(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_122),
.A2(n_102),
.B(n_95),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_137),
.A2(n_115),
.B(n_133),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_118),
.A2(n_95),
.B(n_102),
.C(n_107),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_134),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_129),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_140),
.C(n_147),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_112),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_109),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_144),
.B(n_126),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_99),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_155),
.B(n_147),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_132),
.B1(n_130),
.B2(n_131),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_125),
.B(n_114),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_135),
.A3(n_136),
.B1(n_137),
.B2(n_140),
.C1(n_119),
.C2(n_139),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_159),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_155),
.B(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_119),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_169),
.B(n_171),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_154),
.B1(n_145),
.B2(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_154),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_172),
.B(n_173),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_145),
.C(n_164),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_167),
.C(n_166),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_174),
.Y(n_178)
);

AOI31xp67_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_169),
.A3(n_165),
.B(n_161),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_117),
.B1(n_108),
.B2(n_97),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_146),
.C(n_156),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_96),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_96),
.B(n_70),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_186),
.B(n_180),
.Y(n_187)
);


endmodule