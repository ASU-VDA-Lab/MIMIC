module fake_jpeg_31113_n_45 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_16),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_25),
.Y(n_26)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_0),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_20),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_20),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_20),
.C(n_8),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.C(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_28),
.B1(n_26),
.B2(n_5),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_1),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_38),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_4),
.C(n_6),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_38),
.B1(n_7),
.B2(n_37),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_40),
.C(n_11),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_10),
.B(n_12),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_14),
.Y(n_45)
);


endmodule