module real_aes_7054_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_792;
wire n_386;
wire n_503;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_889;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_867;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_756;
wire n_713;
wire n_598;
wire n_288;
wire n_735;
wire n_404;
wire n_728;
wire n_334;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_712;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_SL g572 ( .A1(n_0), .A2(n_241), .B1(n_521), .B2(n_559), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_1), .A2(n_275), .B1(n_553), .B2(n_554), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_2), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_3), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_4), .A2(n_234), .B1(n_333), .B2(n_336), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_5), .A2(n_127), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_6), .A2(n_23), .B1(n_398), .B2(n_399), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_7), .A2(n_70), .B1(n_369), .B2(n_432), .Y(n_431) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_8), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_9), .A2(n_249), .B1(n_867), .B2(n_868), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_10), .A2(n_80), .B1(n_326), .B2(n_681), .Y(n_869) );
INVx1_ASAP7_75t_L g535 ( .A(n_11), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_12), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_13), .A2(n_139), .B1(n_406), .B2(n_653), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_14), .A2(n_266), .B1(n_598), .B2(n_862), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_15), .A2(n_182), .B1(n_372), .B2(n_549), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_16), .A2(n_111), .B1(n_364), .B2(n_598), .Y(n_897) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_17), .A2(n_158), .B1(n_409), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_18), .A2(n_238), .B1(n_440), .B2(n_611), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_19), .A2(n_125), .B1(n_367), .B2(n_550), .Y(n_863) );
INVx1_ASAP7_75t_L g893 ( .A(n_20), .Y(n_893) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_21), .A2(n_169), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_22), .A2(n_184), .B1(n_483), .B2(n_485), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_24), .A2(n_150), .B1(n_361), .B2(n_364), .Y(n_360) );
INVx1_ASAP7_75t_L g456 ( .A(n_25), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g751 ( .A1(n_26), .A2(n_63), .B1(n_553), .B2(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_27), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_28), .A2(n_152), .B1(n_550), .B2(n_605), .Y(n_894) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_29), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_30), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_31), .A2(n_179), .B1(n_611), .B2(n_648), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_32), .A2(n_278), .B1(n_324), .B2(n_407), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_33), .A2(n_240), .B1(n_394), .B2(n_437), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_34), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_35), .A2(n_133), .B1(n_350), .B2(n_561), .Y(n_721) );
AO22x2_ASAP7_75t_L g313 ( .A1(n_36), .A2(n_97), .B1(n_314), .B2(n_315), .Y(n_313) );
INVx1_ASAP7_75t_L g850 ( .A(n_36), .Y(n_850) );
NAND2xp5_ASAP7_75t_SL g825 ( .A(n_37), .B(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_38), .A2(n_218), .B1(n_399), .B2(n_515), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_39), .A2(n_168), .B1(n_356), .B2(n_490), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_40), .A2(n_172), .B1(n_446), .B2(n_570), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_41), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_42), .A2(n_260), .B1(n_440), .B2(n_441), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g900 ( .A1(n_43), .A2(n_224), .B1(n_479), .B2(n_485), .Y(n_900) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_44), .A2(n_202), .B1(n_253), .B2(n_377), .C1(n_380), .C2(n_384), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_45), .Y(n_493) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_46), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_47), .A2(n_142), .B1(n_488), .B2(n_492), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g749 ( .A1(n_48), .A2(n_198), .B1(n_549), .B2(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_49), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_50), .Y(n_603) );
INVx1_ASAP7_75t_L g434 ( .A(n_51), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_52), .Y(n_730) );
AO22x2_ASAP7_75t_L g317 ( .A1(n_53), .A2(n_100), .B1(n_314), .B2(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g851 ( .A(n_53), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_54), .A2(n_144), .B1(n_373), .B2(n_385), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_55), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_56), .A2(n_156), .B1(n_712), .B2(n_713), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_57), .A2(n_186), .B1(n_369), .B2(n_750), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_58), .A2(n_272), .B1(n_401), .B2(n_402), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_59), .A2(n_171), .B1(n_446), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_60), .A2(n_230), .B1(n_380), .B2(n_811), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_61), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_62), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g755 ( .A1(n_64), .A2(n_71), .B1(n_677), .B2(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_65), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_66), .A2(n_257), .B1(n_384), .B2(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_67), .A2(n_136), .B1(n_670), .B2(n_671), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_68), .A2(n_854), .B1(n_873), .B2(n_874), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_68), .Y(n_873) );
AOI222xp33_ASAP7_75t_L g815 ( .A1(n_69), .A2(n_197), .B1(n_265), .B2(n_377), .C1(n_515), .C2(n_605), .Y(n_815) );
AOI22xp5_ASAP7_75t_SL g569 ( .A1(n_72), .A2(n_165), .B1(n_342), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_73), .A2(n_258), .B1(n_441), .B2(n_488), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_74), .A2(n_270), .B1(n_744), .B2(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_75), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_76), .Y(n_626) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_77), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_78), .A2(n_280), .B1(n_333), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_79), .A2(n_203), .B1(n_561), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_81), .A2(n_193), .B1(n_409), .B2(n_574), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_82), .A2(n_208), .B1(n_333), .B2(n_409), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_83), .A2(n_201), .B1(n_367), .B2(n_550), .Y(n_728) );
AOI22xp5_ASAP7_75t_SL g568 ( .A1(n_84), .A2(n_151), .B1(n_441), .B2(n_485), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_85), .A2(n_227), .B1(n_365), .B2(n_401), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_86), .Y(n_632) );
AO22x2_ASAP7_75t_L g622 ( .A1(n_87), .A2(n_623), .B1(n_654), .B2(n_655), .Y(n_622) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_87), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_88), .A2(n_237), .B1(n_647), .B2(n_648), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_89), .A2(n_173), .B1(n_687), .B2(n_688), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_90), .Y(n_594) );
AOI211xp5_ASAP7_75t_L g591 ( .A1(n_91), .A2(n_592), .B(n_593), .C(n_600), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_92), .A2(n_244), .B1(n_666), .B2(n_667), .Y(n_665) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_93), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_94), .A2(n_159), .B1(n_406), .B2(n_407), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g757 ( .A1(n_95), .A2(n_116), .B1(n_653), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g449 ( .A(n_96), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_98), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_99), .A2(n_276), .B1(n_342), .B2(n_344), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_101), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_102), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_103), .A2(n_212), .B1(n_334), .B2(n_356), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_104), .A2(n_772), .B1(n_798), .B2(n_799), .Y(n_771) );
INVx1_ASAP7_75t_L g798 ( .A(n_104), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_105), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_106), .Y(n_816) );
INVx1_ASAP7_75t_L g294 ( .A(n_107), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_108), .A2(n_267), .B1(n_350), .B2(n_355), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_109), .A2(n_210), .B1(n_409), .B2(n_411), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_110), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_112), .A2(n_214), .B1(n_448), .B2(n_490), .Y(n_609) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_113), .Y(n_673) );
INVx1_ASAP7_75t_L g292 ( .A(n_114), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_115), .A2(n_178), .B1(n_415), .B2(n_417), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_117), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_118), .Y(n_783) );
XOR2x2_ASAP7_75t_L g303 ( .A(n_119), .B(n_304), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_120), .A2(n_242), .B1(n_440), .B2(n_564), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g822 ( .A1(n_121), .A2(n_157), .B1(n_385), .B2(n_515), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_122), .B(n_402), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_123), .A2(n_131), .B1(n_574), .B2(n_648), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_124), .A2(n_229), .B1(n_712), .B2(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g508 ( .A(n_126), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_128), .A2(n_164), .B1(n_750), .B2(n_811), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g583 ( .A(n_129), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g759 ( .A1(n_130), .A2(n_681), .B(n_760), .C(n_765), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_132), .A2(n_163), .B1(n_561), .B2(n_791), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_134), .B(n_692), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g685 ( .A(n_135), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_137), .A2(n_226), .B1(n_558), .B2(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_138), .B(n_402), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_140), .A2(n_213), .B1(n_795), .B2(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g536 ( .A(n_141), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_143), .A2(n_243), .B1(n_367), .B2(n_372), .Y(n_366) );
INVx1_ASAP7_75t_L g883 ( .A(n_145), .Y(n_883) );
AOI22xp5_ASAP7_75t_SL g887 ( .A1(n_145), .A2(n_883), .B1(n_888), .B2(n_889), .Y(n_887) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_146), .A2(n_192), .B1(n_373), .B2(n_394), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_147), .A2(n_220), .B1(n_549), .B2(n_550), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_148), .A2(n_188), .B1(n_481), .B2(n_681), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_149), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_153), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_154), .B(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g295 ( .A(n_155), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_160), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_161), .A2(n_191), .B1(n_350), .B2(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g601 ( .A(n_162), .Y(n_601) );
AND2x6_ASAP7_75t_L g291 ( .A(n_166), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g844 ( .A(n_166), .Y(n_844) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_167), .A2(n_235), .B1(n_314), .B2(n_318), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g589 ( .A(n_170), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_174), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_175), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_176), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_177), .A2(n_211), .B1(n_440), .B2(n_485), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_180), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_181), .Y(n_524) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_183), .A2(n_262), .B1(n_411), .B2(n_446), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_185), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g782 ( .A(n_187), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_189), .A2(n_703), .B1(n_734), .B2(n_735), .Y(n_702) );
INVx1_ASAP7_75t_L g734 ( .A(n_189), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g419 ( .A(n_190), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_194), .A2(n_264), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI22xp33_ASAP7_75t_SL g832 ( .A1(n_195), .A2(n_254), .B1(n_406), .B2(n_407), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_196), .Y(n_472) );
AO22x2_ASAP7_75t_L g323 ( .A1(n_199), .A2(n_251), .B1(n_314), .B2(n_315), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_200), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_204), .A2(n_255), .B1(n_605), .B2(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g619 ( .A(n_205), .Y(n_619) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_206), .Y(n_682) );
INVx1_ASAP7_75t_L g505 ( .A(n_207), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_209), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_215), .A2(n_281), .B1(n_436), .B2(n_437), .Y(n_435) );
INVx1_ASAP7_75t_L g532 ( .A(n_216), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_217), .B(n_361), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_219), .A2(n_256), .B1(n_485), .B2(n_570), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_221), .B(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_222), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_223), .A2(n_252), .B1(n_356), .B2(n_647), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_225), .A2(n_274), .B1(n_479), .B2(n_481), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_228), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g615 ( .A(n_231), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g442 ( .A1(n_232), .A2(n_239), .B1(n_443), .B2(n_444), .Y(n_442) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_233), .A2(n_287), .B(n_296), .C(n_852), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_235), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_236), .B(n_402), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_245), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g628 ( .A(n_246), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_247), .A2(n_259), .B1(n_402), .B2(n_598), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_248), .A2(n_661), .B1(n_662), .B2(n_694), .Y(n_660) );
INVx1_ASAP7_75t_L g694 ( .A(n_248), .Y(n_694) );
XNOR2xp5_ASAP7_75t_L g738 ( .A(n_250), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g847 ( .A(n_251), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_261), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_263), .A2(n_285), .B1(n_479), .B2(n_483), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_268), .A2(n_273), .B1(n_307), .B2(n_324), .Y(n_306) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_269), .Y(n_780) );
INVx1_ASAP7_75t_L g314 ( .A(n_271), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_271), .Y(n_316) );
INVx1_ASAP7_75t_L g461 ( .A(n_277), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_279), .A2(n_284), .B1(n_791), .B2(n_792), .Y(n_790) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_282), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_283), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_292), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_293), .A2(n_842), .B(n_882), .Y(n_881) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_698), .B1(n_837), .B2(n_838), .C(n_839), .Y(n_296) );
INVx1_ASAP7_75t_L g837 ( .A(n_297), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_496), .B1(n_696), .B2(n_697), .Y(n_297) );
INVx1_ASAP7_75t_L g696 ( .A(n_298), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B1(n_422), .B2(n_495), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AO22x1_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_387), .B1(n_420), .B2(n_421), .Y(n_302) );
INVx1_ASAP7_75t_L g420 ( .A(n_303), .Y(n_420) );
NAND4xp75_ASAP7_75t_L g304 ( .A(n_305), .B(n_340), .C(n_359), .D(n_376), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_332), .Y(n_305) );
INVx4_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx3_ASAP7_75t_L g485 ( .A(n_308), .Y(n_485) );
INVx4_ASAP7_75t_L g564 ( .A(n_308), .Y(n_564) );
INVx2_ASAP7_75t_SL g795 ( .A(n_308), .Y(n_795) );
INVx11_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx11_ASAP7_75t_L g412 ( .A(n_309), .Y(n_412) );
AND2x6_ASAP7_75t_L g309 ( .A(n_310), .B(n_319), .Y(n_309) );
AND2x4_ASAP7_75t_L g363 ( .A(n_310), .B(n_335), .Y(n_363) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g459 ( .A(n_311), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_317), .Y(n_311) );
AND2x2_ASAP7_75t_L g330 ( .A(n_312), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g348 ( .A(n_312), .B(n_317), .Y(n_348) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g371 ( .A(n_313), .B(n_321), .Y(n_371) );
AND2x2_ASAP7_75t_L g375 ( .A(n_313), .B(n_317), .Y(n_375) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g318 ( .A(n_316), .Y(n_318) );
INVx2_ASAP7_75t_L g331 ( .A(n_317), .Y(n_331) );
INVx1_ASAP7_75t_L g358 ( .A(n_317), .Y(n_358) );
AND2x2_ASAP7_75t_L g343 ( .A(n_319), .B(n_330), .Y(n_343) );
AND2x4_ASAP7_75t_L g347 ( .A(n_319), .B(n_348), .Y(n_347) );
AND2x6_ASAP7_75t_L g379 ( .A(n_319), .B(n_375), .Y(n_379) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g335 ( .A(n_320), .B(n_323), .Y(n_335) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g328 ( .A(n_321), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_321), .B(n_323), .Y(n_339) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g329 ( .A(n_323), .Y(n_329) );
INVx1_ASAP7_75t_L g383 ( .A(n_323), .Y(n_383) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g406 ( .A(n_327), .Y(n_406) );
BUFx3_ASAP7_75t_L g446 ( .A(n_327), .Y(n_446) );
BUFx3_ASAP7_75t_L g480 ( .A(n_327), .Y(n_480) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
AND2x2_ASAP7_75t_L g354 ( .A(n_328), .B(n_348), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_328), .B(n_348), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_328), .B(n_330), .Y(n_533) );
INVx1_ASAP7_75t_L g374 ( .A(n_329), .Y(n_374) );
AND2x4_ASAP7_75t_L g334 ( .A(n_330), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g337 ( .A(n_330), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g382 ( .A(n_331), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g475 ( .A(n_331), .Y(n_475) );
BUFx2_ASAP7_75t_L g717 ( .A(n_333), .Y(n_717) );
BUFx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g443 ( .A(n_334), .Y(n_443) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_334), .Y(n_492) );
INVx2_ASAP7_75t_L g518 ( .A(n_334), .Y(n_518) );
BUFx3_ASAP7_75t_L g574 ( .A(n_334), .Y(n_574) );
AND2x6_ASAP7_75t_L g365 ( .A(n_335), .B(n_348), .Y(n_365) );
INVx1_ASAP7_75t_L g460 ( .A(n_335), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_335), .B(n_348), .Y(n_463) );
INVx2_ASAP7_75t_L g668 ( .A(n_336), .Y(n_668) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx3_ASAP7_75t_L g407 ( .A(n_337), .Y(n_407) );
BUFx2_ASAP7_75t_L g448 ( .A(n_337), .Y(n_448) );
BUFx2_ASAP7_75t_SL g481 ( .A(n_337), .Y(n_481) );
INVx1_ASAP7_75t_L g528 ( .A(n_337), .Y(n_528) );
BUFx3_ASAP7_75t_L g559 ( .A(n_337), .Y(n_559) );
BUFx3_ASAP7_75t_L g653 ( .A(n_337), .Y(n_653) );
BUFx2_ASAP7_75t_SL g868 ( .A(n_337), .Y(n_868) );
AND2x2_ASAP7_75t_L g521 ( .A(n_338), .B(n_475), .Y(n_521) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x6_ASAP7_75t_L g357 ( .A(n_339), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_349), .Y(n_340) );
BUFx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g410 ( .A(n_343), .Y(n_410) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_343), .Y(n_484) );
BUFx2_ASAP7_75t_SL g681 ( .A(n_343), .Y(n_681) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx6_ASAP7_75t_L g416 ( .A(n_347), .Y(n_416) );
BUFx3_ASAP7_75t_L g570 ( .A(n_347), .Y(n_570) );
BUFx3_ASAP7_75t_L g677 ( .A(n_347), .Y(n_677) );
INVx3_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx6f_ASAP7_75t_L g670 ( .A(n_352), .Y(n_670) );
INVx4_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx5_ASAP7_75t_L g417 ( .A(n_353), .Y(n_417) );
INVx3_ASAP7_75t_L g441 ( .A(n_353), .Y(n_441) );
INVx1_ASAP7_75t_L g611 ( .A(n_353), .Y(n_611) );
INVx2_ASAP7_75t_L g647 ( .A(n_353), .Y(n_647) );
INVx8_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g648 ( .A(n_356), .Y(n_648) );
BUFx2_ASAP7_75t_L g671 ( .A(n_356), .Y(n_671) );
BUFx4f_ASAP7_75t_SL g792 ( .A(n_356), .Y(n_792) );
INVx6_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g444 ( .A(n_357), .Y(n_444) );
INVx1_ASAP7_75t_SL g561 ( .A(n_357), .Y(n_561) );
INVx1_ASAP7_75t_L g370 ( .A(n_358), .Y(n_370) );
AND2x2_ASAP7_75t_SL g359 ( .A(n_360), .B(n_366), .Y(n_359) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx5_ASAP7_75t_L g401 ( .A(n_362), .Y(n_401) );
INVx2_ASAP7_75t_L g598 ( .A(n_362), .Y(n_598) );
INVx2_ASAP7_75t_L g826 ( .A(n_362), .Y(n_826) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx4f_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_SL g555 ( .A(n_365), .Y(n_555) );
BUFx2_ASAP7_75t_L g862 ( .A(n_365), .Y(n_862) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
BUFx2_ASAP7_75t_L g549 ( .A(n_369), .Y(n_549) );
BUFx2_ASAP7_75t_L g811 ( .A(n_369), .Y(n_811) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AND2x4_ASAP7_75t_L g381 ( .A(n_371), .B(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g385 ( .A(n_371), .B(n_386), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_371), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g551 ( .A(n_372), .Y(n_551) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_SL g395 ( .A(n_373), .Y(n_395) );
BUFx2_ASAP7_75t_SL g437 ( .A(n_373), .Y(n_437) );
BUFx3_ASAP7_75t_L g750 ( .A(n_373), .Y(n_750) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g643 ( .A(n_374), .Y(n_643) );
INVx1_ASAP7_75t_L g642 ( .A(n_375), .Y(n_642) );
INVx2_ASAP7_75t_L g892 ( .A(n_377), .Y(n_892) );
INVx4_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI21xp5_ASAP7_75t_SL g684 ( .A1(n_378), .A2(n_685), .B(n_686), .Y(n_684) );
INVx4_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g392 ( .A(n_379), .Y(n_392) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_379), .Y(n_467) );
INVx2_ASAP7_75t_SL g512 ( .A(n_379), .Y(n_512) );
INVx2_ASAP7_75t_L g578 ( .A(n_379), .Y(n_578) );
BUFx3_ASAP7_75t_L g592 ( .A(n_379), .Y(n_592) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx4f_ASAP7_75t_SL g398 ( .A(n_381), .Y(n_398) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_381), .Y(n_515) );
BUFx2_ASAP7_75t_L g635 ( .A(n_381), .Y(n_635) );
INVx1_ASAP7_75t_L g386 ( .A(n_383), .Y(n_386) );
BUFx4f_ASAP7_75t_L g688 ( .A(n_384), .Y(n_688) );
INVx1_ASAP7_75t_L g746 ( .A(n_384), .Y(n_746) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx12f_ASAP7_75t_L g394 ( .A(n_385), .Y(n_394) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_385), .Y(n_436) );
INVx3_ASAP7_75t_SL g421 ( .A(n_387), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_387), .A2(n_421), .B1(n_451), .B2(n_452), .Y(n_450) );
XOR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_419), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_389), .B(n_403), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_396), .Y(n_389) );
OAI21xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B(n_393), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_392), .A2(n_434), .B(n_435), .Y(n_433) );
OAI21xp5_ASAP7_75t_SL g820 ( .A1(n_392), .A2(n_821), .B(n_822), .Y(n_820) );
OAI21xp5_ASAP7_75t_SL g856 ( .A1(n_392), .A2(n_857), .B(n_858), .Y(n_856) );
INVx2_ASAP7_75t_L g606 ( .A(n_394), .Y(n_606) );
BUFx4f_ASAP7_75t_SL g859 ( .A(n_394), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_401), .Y(n_553) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_401), .Y(n_692) );
INVx1_ASAP7_75t_L g753 ( .A(n_402), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_413), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI22xp5_ASAP7_75t_SL g522 ( .A1(n_410), .A2(n_416), .B1(n_523), .B2(n_524), .Y(n_522) );
INVx3_ASAP7_75t_L g650 ( .A(n_410), .Y(n_650) );
INVx1_ASAP7_75t_L g674 ( .A(n_411), .Y(n_674) );
INVx5_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_412), .B(n_535), .Y(n_534) );
INVx2_ASAP7_75t_SL g652 ( .A(n_412), .Y(n_652) );
INVx1_ASAP7_75t_L g707 ( .A(n_412), .Y(n_707) );
INVx2_ASAP7_75t_L g867 ( .A(n_412), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .Y(n_413) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
INVx2_ASAP7_75t_L g488 ( .A(n_416), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_416), .A2(n_613), .B1(n_614), .B2(n_615), .Y(n_612) );
INVx2_ASAP7_75t_L g796 ( .A(n_416), .Y(n_796) );
BUFx6f_ASAP7_75t_L g791 ( .A(n_417), .Y(n_791) );
INVx2_ASAP7_75t_L g495 ( .A(n_422), .Y(n_495) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OA22x2_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_450), .B2(n_494), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
XOR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_449), .Y(n_425) );
NAND4xp75_ASAP7_75t_SL g426 ( .A(n_427), .B(n_438), .C(n_445), .D(n_447), .Y(n_426) );
NOR2xp67_ASAP7_75t_SL g427 ( .A(n_428), .B(n_433), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .C(n_431), .Y(n_428) );
INVx1_ASAP7_75t_L g602 ( .A(n_432), .Y(n_602) );
BUFx6f_ASAP7_75t_L g744 ( .A(n_432), .Y(n_744) );
INVx2_ASAP7_75t_L g732 ( .A(n_436), .Y(n_732) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_442), .Y(n_438) );
BUFx2_ASAP7_75t_L g756 ( .A(n_446), .Y(n_756) );
INVx1_ASAP7_75t_L g494 ( .A(n_450), .Y(n_494) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
XNOR2x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_493), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_476), .Y(n_453) );
NOR3xp33_ASAP7_75t_L g454 ( .A(n_455), .B(n_464), .C(n_469), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_461), .B2(n_462), .Y(n_455) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g627 ( .A(n_458), .Y(n_627) );
INVx2_ASAP7_75t_L g724 ( .A(n_458), .Y(n_724) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_459), .A2(n_505), .B(n_506), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_462), .A2(n_474), .B1(n_508), .B2(n_509), .Y(n_507) );
INVx2_ASAP7_75t_L g596 ( .A(n_462), .Y(n_596) );
BUFx3_ASAP7_75t_L g726 ( .A(n_462), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_462), .A2(n_627), .B1(n_775), .B2(n_776), .Y(n_774) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g630 ( .A(n_463), .Y(n_630) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_468), .Y(n_464) );
OAI222xp33_ASAP7_75t_L g777 ( .A1(n_466), .A2(n_514), .B1(n_732), .B2(n_778), .C1(n_779), .C2(n_780), .Y(n_777) );
INVx2_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_469) );
OAI222xp33_ASAP7_75t_L g729 ( .A1(n_471), .A2(n_512), .B1(n_730), .B2(n_731), .C1(n_732), .C2(n_733), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_473), .A2(n_782), .B1(n_783), .B2(n_784), .Y(n_781) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx4_ASAP7_75t_L g639 ( .A(n_474), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_482), .Y(n_477) );
BUFx4f_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g714 ( .A(n_480), .Y(n_714) );
INVx1_ASAP7_75t_L g719 ( .A(n_481), .Y(n_719) );
INVx1_ASAP7_75t_SL g618 ( .A(n_483), .Y(n_618) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g712 ( .A(n_484), .Y(n_712) );
INVx1_ASAP7_75t_L g614 ( .A(n_485), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
INVx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g666 ( .A(n_491), .Y(n_666) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g697 ( .A(n_496), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_584), .B1(n_585), .B2(n_695), .Y(n_496) );
INVx1_ASAP7_75t_SL g695 ( .A(n_497), .Y(n_695) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
XNOR2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_537), .Y(n_499) );
BUFx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
XNOR2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_536), .Y(n_501) );
AND3x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_516), .C(n_525), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .C(n_510), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_510) );
INVx3_ASAP7_75t_L g687 ( .A(n_514), .Y(n_687) );
INVx4_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g546 ( .A(n_515), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_517), .B(n_522), .Y(n_516) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_519), .B(n_520), .Y(n_517) );
INVx2_ASAP7_75t_L g558 ( .A(n_518), .Y(n_558) );
INVx1_ASAP7_75t_L g789 ( .A(n_518), .Y(n_789) );
NOR3xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_531), .C(n_534), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_529), .B2(n_530), .Y(n_526) );
BUFx2_ASAP7_75t_R g761 ( .A(n_530), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g621 ( .A(n_533), .Y(n_621) );
XOR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_566), .Y(n_537) );
XNOR2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_556), .C(n_562), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_547), .Y(n_541) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_544), .B(n_545), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_560), .Y(n_556) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g767 ( .A(n_564), .Y(n_767) );
XOR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_583), .Y(n_566) );
NAND4xp75_ASAP7_75t_SL g567 ( .A(n_568), .B(n_569), .C(n_571), .D(n_575), .Y(n_567) );
INVx1_ASAP7_75t_L g709 ( .A(n_570), .Y(n_709) );
AND2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_574), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_580), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B(n_579), .Y(n_576) );
OAI222xp33_ASAP7_75t_L g741 ( .A1(n_578), .A2(n_742), .B1(n_743), .B2(n_745), .C1(n_746), .C2(n_747), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
XNOR2xp5_ASAP7_75t_SL g585 ( .A(n_586), .B(n_658), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_622), .B1(n_656), .B2(n_657), .Y(n_587) );
INVx2_ASAP7_75t_L g656 ( .A(n_588), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_607), .Y(n_590) );
INVx3_ASAP7_75t_L g633 ( .A(n_592), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B(n_597), .C(n_599), .Y(n_593) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_612), .C(n_616), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_619), .B2(n_620), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_620), .A2(n_679), .B1(n_680), .B2(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g657 ( .A(n_622), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g659 ( .A(n_622), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g654 ( .A(n_623), .Y(n_654) );
AND2x2_ASAP7_75t_SL g623 ( .A(n_624), .B(n_644), .Y(n_623) );
NOR3xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_631), .C(n_636), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_628), .B2(n_629), .Y(n_625) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OAI21xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_634), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B1(n_640), .B2(n_641), .Y(n_636) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
CKINVDCx16_ASAP7_75t_R g785 ( .A(n_641), .Y(n_785) );
OR2x6_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
AND4x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .C(n_649), .D(n_651), .Y(n_644) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_663), .B(n_683), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_664), .B(n_672), .C(n_678), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_669), .Y(n_664) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g763 ( .A(n_671), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_675), .B2(n_676), .Y(n_672) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_689), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .C(n_693), .Y(n_689) );
INVx1_ASAP7_75t_L g838 ( .A(n_698), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B1(n_768), .B2(n_836), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI22xp5_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_702), .B1(n_736), .B2(n_737), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g735 ( .A(n_703), .Y(n_735) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_722), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_705), .B(n_715), .Y(n_704) );
OAI221xp5_ASAP7_75t_SL g705 ( .A1(n_706), .A2(n_708), .B1(n_709), .B2(n_710), .C(n_711), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI221xp5_ASAP7_75t_SL g715 ( .A1(n_716), .A2(n_718), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NOR2xp33_ASAP7_75t_SL g722 ( .A(n_723), .B(n_729), .Y(n_722) );
OAI221xp5_ASAP7_75t_SL g723 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_727), .C(n_728), .Y(n_723) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NAND3x1_ASAP7_75t_L g739 ( .A(n_740), .B(n_754), .C(n_759), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_748), .Y(n_740) );
INVx2_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g754 ( .A(n_755), .B(n_757), .Y(n_754) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx3_ASAP7_75t_L g836 ( .A(n_768), .Y(n_836) );
BUFx3_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_800), .B2(n_801), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g799 ( .A(n_772), .Y(n_799) );
AND2x2_ASAP7_75t_L g772 ( .A(n_773), .B(n_786), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_774), .B(n_777), .C(n_781), .Y(n_773) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_793), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_794), .B(n_797), .Y(n_793) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
AO22x2_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_803), .B1(n_817), .B2(n_835), .Y(n_801) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
XOR2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_816), .Y(n_803) );
NAND4xp75_ASAP7_75t_L g804 ( .A(n_805), .B(n_808), .C(n_812), .D(n_815), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_SL g808 ( .A(n_809), .B(n_810), .Y(n_808) );
AND2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx4_ASAP7_75t_SL g835 ( .A(n_817), .Y(n_835) );
XOR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_834), .Y(n_817) );
NAND3x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_828), .C(n_831), .Y(n_818) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_823), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .C(n_827), .Y(n_823) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
INVx1_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
NOR2x1_ASAP7_75t_L g840 ( .A(n_841), .B(n_845), .Y(n_840) );
OR2x2_ASAP7_75t_SL g907 ( .A(n_841), .B(n_846), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_842), .B(n_844), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g875 ( .A(n_843), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_843), .B(n_879), .Y(n_882) );
CKINVDCx16_ASAP7_75t_R g879 ( .A(n_844), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g845 ( .A(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
OAI322xp33_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_875), .A3(n_876), .B1(n_880), .B2(n_883), .C1(n_884), .C2(n_905), .Y(n_852) );
INVx2_ASAP7_75t_SL g874 ( .A(n_854), .Y(n_874) );
AND2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_864), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_861), .B(n_863), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_870), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_869), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
CKINVDCx20_ASAP7_75t_R g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_SL g888 ( .A(n_889), .Y(n_888) );
NAND2xp5_ASAP7_75t_SL g889 ( .A(n_890), .B(n_898), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g890 ( .A(n_891), .B(n_895), .Y(n_890) );
OAI21xp5_ASAP7_75t_SL g891 ( .A1(n_892), .A2(n_893), .B(n_894), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_897), .Y(n_895) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_902), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_901), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g905 ( .A(n_906), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_907), .Y(n_906) );
endmodule