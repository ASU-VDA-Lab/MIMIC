module fake_jpeg_27327_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_23),
.B1(n_40),
.B2(n_39),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_51),
.B1(n_49),
.B2(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_41),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_52),
.B1(n_47),
.B2(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_63),
.A2(n_64),
.B1(n_3),
.B2(n_6),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_54),
.B1(n_55),
.B2(n_48),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_8),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_72),
.B(n_74),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_73),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_77),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_6),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_90),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_14),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_82),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_98),
.B(n_86),
.CON(n_105),
.SN(n_105)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_31),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_101),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_85),
.Y(n_104)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_105),
.A2(n_107),
.B1(n_93),
.B2(n_96),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_32),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_105),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_115),
.C(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_117),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_109),
.Y(n_121)
);

AOI21x1_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_112),
.B(n_94),
.Y(n_122)
);

AOI322xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_89),
.A3(n_84),
.B1(n_106),
.B2(n_36),
.C1(n_37),
.C2(n_33),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_34),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_35),
.Y(n_125)
);


endmodule