module real_jpeg_19053_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

OAI32xp33_ASAP7_75t_L g32 ( 
.A1(n_0),
.A2(n_33),
.A3(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_32)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_35),
.B1(n_38),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_3),
.A2(n_33),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_3),
.B(n_75),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_24),
.B(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_3),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_3),
.A2(n_26),
.B1(n_109),
.B2(n_110),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_3),
.B(n_69),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_5),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_91)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_5),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_35),
.B1(n_38),
.B2(n_49),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_49),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_8),
.A2(n_35),
.B1(n_38),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_58),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_58),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_10),
.A2(n_25),
.B1(n_35),
.B2(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_76),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_87),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_86),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_61),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_18),
.B(n_61),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.C(n_50),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_19),
.A2(n_20),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_32),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_32),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_22),
.A2(n_26),
.B1(n_30),
.B2(n_96),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_23),
.A2(n_24),
.B1(n_54),
.B2(n_55),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_113),
.Y(n_112)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_26),
.A2(n_94),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_40),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_37),
.B(n_44),
.C(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_35),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_35),
.A2(n_40),
.B(n_55),
.C(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_40),
.B(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_40),
.B(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_41),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_56),
.B1(n_59),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_52),
.A2(n_56),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_52),
.A2(n_56),
.B1(n_57),
.B2(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_79),
.B2(n_80),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_127),
.B(n_132),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_117),
.B(n_126),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_105),
.B(n_116),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_97),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_101),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_111),
.B(n_115),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_108),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_119),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_125),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_124),
.C(n_125),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_129),
.Y(n_132)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_130),
.Y(n_131)
);


endmodule