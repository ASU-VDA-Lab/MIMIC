module fake_jpeg_2354_n_121 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_16),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_45),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_1),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_49),
.B(n_43),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_39),
.B1(n_34),
.B2(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_58),
.B(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_2),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_42),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_39),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_71),
.A2(n_40),
.B1(n_53),
.B2(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_17),
.B1(n_29),
.B2(n_27),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_83),
.Y(n_86)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_3),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_3),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_13),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_91),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_40),
.B1(n_19),
.B2(n_20),
.Y(n_87)
);

AOI21x1_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_73),
.B(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_12),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_14),
.B1(n_26),
.B2(n_24),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_9),
.B1(n_22),
.B2(n_23),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_7),
.Y(n_102)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_8),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_32),
.C(n_9),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_110),
.A2(n_88),
.B(n_87),
.Y(n_112)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_106),
.C(n_97),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_114),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_116),
.A2(n_107),
.B(n_109),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_92),
.B(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_94),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_100),
.B(n_105),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_109),
.Y(n_121)
);


endmodule