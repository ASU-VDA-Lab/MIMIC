module fake_jpeg_21458_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_5),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_16),
.B1(n_15),
.B2(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_22),
.Y(n_23)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_25),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_16),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_21),
.C(n_14),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_18),
.B(n_11),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_32),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_31),
.C(n_35),
.Y(n_38)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_17),
.B1(n_12),
.B2(n_9),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_15),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_12),
.B1(n_8),
.B2(n_10),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_26),
.B2(n_27),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_1),
.C(n_2),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_24),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_31),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_38),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_24),
.C(n_26),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_38),
.C(n_39),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_37),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_45),
.B(n_4),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_48),
.C(n_24),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_1),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_48),
.C(n_24),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_4),
.B1(n_6),
.B2(n_43),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_6),
.Y(n_55)
);


endmodule