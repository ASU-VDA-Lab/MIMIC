module fake_jpeg_6762_n_180 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_22),
.Y(n_49)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_31),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_39),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_27),
.C(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_27),
.B1(n_20),
.B2(n_23),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_21),
.B1(n_15),
.B2(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_19),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_53),
.B1(n_30),
.B2(n_16),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_54),
.B(n_56),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_49),
.B1(n_43),
.B2(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_32),
.B1(n_19),
.B2(n_22),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_45),
.B(n_52),
.C(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_65),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_15),
.B1(n_28),
.B2(n_25),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_81),
.B1(n_83),
.B2(n_1),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_78),
.Y(n_90)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_65),
.B(n_48),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_76),
.A2(n_87),
.B(n_3),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_51),
.B1(n_16),
.B2(n_45),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_12),
.B(n_4),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_40),
.B1(n_31),
.B2(n_26),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_59),
.A3(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_88),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_38),
.B1(n_26),
.B2(n_10),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_62),
.B1(n_2),
.B2(n_3),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_38),
.C(n_13),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_58),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_96),
.A2(n_73),
.B1(n_75),
.B2(n_12),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_104),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_11),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_79),
.B(n_4),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_106),
.A2(n_99),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_74),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_106),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_79),
.C(n_71),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_93),
.C(n_96),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_75),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_131),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_90),
.A3(n_118),
.B1(n_117),
.B2(n_107),
.C1(n_102),
.C2(n_100),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_109),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_104),
.B1(n_94),
.B2(n_90),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_109),
.C(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_132),
.C(n_129),
.Y(n_147)
);

XOR2x2_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_134),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_136),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_111),
.B1(n_116),
.B2(n_108),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_142),
.A2(n_127),
.B1(n_130),
.B2(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_131),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_149),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_113),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_155),
.C(n_145),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_139),
.A2(n_141),
.B(n_135),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_152),
.A2(n_142),
.B1(n_111),
.B2(n_73),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_135),
.C(n_121),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_140),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_159),
.B(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_149),
.B(n_153),
.C(n_67),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_3),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_157),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_162),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_165),
.A2(n_166),
.B(n_167),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_85),
.B1(n_57),
.B2(n_6),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_169),
.A2(n_172),
.B(n_168),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_85),
.B(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_170),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_175),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_85),
.C(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_5),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_176),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_6),
.Y(n_180)
);


endmodule