module real_aes_17990_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_863, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_863;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g856 ( .A(n_0), .B(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_1), .A2(n_35), .B1(n_138), .B2(n_161), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_2), .A2(n_9), .B1(n_180), .B2(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g857 ( .A(n_3), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_4), .Y(n_136) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_5), .A2(n_11), .B1(n_197), .B2(n_200), .Y(n_196) );
OR2x2_ASAP7_75t_L g116 ( .A(n_6), .B(n_31), .Y(n_116) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_7), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_8), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_10), .Y(n_832) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_12), .B(n_141), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_13), .A2(n_101), .B1(n_180), .B2(n_181), .Y(n_179) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_14), .A2(n_32), .B1(n_146), .B2(n_213), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_15), .A2(n_18), .B1(n_806), .B2(n_807), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_15), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_16), .B(n_141), .Y(n_140) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_17), .A2(n_48), .B(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g807 ( .A(n_18), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_19), .B(n_504), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_20), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_21), .A2(n_39), .B1(n_166), .B2(n_167), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_22), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_23), .A2(n_46), .B1(n_167), .B2(n_180), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_24), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_25), .B(n_146), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_26), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_27), .B(n_198), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_28), .A2(n_105), .B1(n_852), .B2(n_858), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_29), .B(n_155), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_30), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_33), .A2(n_85), .B1(n_138), .B2(n_236), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_34), .A2(n_38), .B1(n_137), .B2(n_138), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_36), .A2(n_51), .B1(n_180), .B2(n_184), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_37), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g844 ( .A1(n_40), .A2(n_831), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_41), .B(n_141), .Y(n_487) );
INVx2_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_43), .A2(n_54), .B1(n_819), .B2(n_820), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_43), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_44), .B(n_142), .Y(n_499) );
BUFx3_ASAP7_75t_L g114 ( .A(n_45), .Y(n_114) );
INVx1_ASAP7_75t_L g829 ( .A(n_45), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_47), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g547 ( .A(n_49), .B(n_507), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_50), .B(n_214), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_52), .B(n_198), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_53), .B(n_166), .Y(n_623) );
INVx1_ASAP7_75t_L g819 ( .A(n_54), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_55), .A2(n_72), .B1(n_166), .B2(n_184), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_56), .A2(n_75), .B1(n_137), .B2(n_138), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_57), .B(n_532), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_58), .A2(n_239), .B(n_488), .C(n_541), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_59), .A2(n_97), .B1(n_180), .B2(n_200), .Y(n_226) );
INVx1_ASAP7_75t_L g133 ( .A(n_60), .Y(n_133) );
AND2x4_ASAP7_75t_L g152 ( .A(n_61), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_62), .A2(n_63), .B1(n_167), .B2(n_217), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_64), .B(n_155), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_65), .B(n_507), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_66), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_67), .B(n_167), .Y(n_492) );
INVx1_ASAP7_75t_L g153 ( .A(n_68), .Y(n_153) );
INVx1_ASAP7_75t_L g830 ( .A(n_69), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_70), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_71), .B(n_155), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_73), .B(n_138), .Y(n_527) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_74), .B(n_142), .C(n_161), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_76), .B(n_138), .Y(n_554) );
INVx2_ASAP7_75t_L g143 ( .A(n_77), .Y(n_143) );
CKINVDCx14_ASAP7_75t_R g474 ( .A(n_78), .Y(n_474) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_78), .A2(n_474), .B1(n_818), .B2(n_821), .Y(n_817) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_79), .B(n_203), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_80), .B(n_141), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_81), .B(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_82), .A2(n_98), .B1(n_167), .B2(n_239), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_83), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_84), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_86), .A2(n_91), .B1(n_198), .B2(n_511), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_87), .B(n_141), .Y(n_620) );
NAND2xp33_ASAP7_75t_SL g572 ( .A(n_88), .B(n_147), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_89), .B(n_182), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_90), .B(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_92), .Y(n_207) );
INVx1_ASAP7_75t_L g471 ( .A(n_93), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_93), .B(n_828), .Y(n_827) );
OAI22x1_ASAP7_75t_SL g803 ( .A1(n_94), .A2(n_804), .B1(n_805), .B2(n_808), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g808 ( .A(n_94), .Y(n_808) );
NAND2xp33_ASAP7_75t_L g148 ( .A(n_95), .B(n_141), .Y(n_148) );
NAND2xp33_ASAP7_75t_L g555 ( .A(n_96), .B(n_147), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_99), .B(n_507), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_100), .B(n_147), .C(n_203), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_102), .B(n_138), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_103), .B(n_198), .Y(n_530) );
AO21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_117), .B(n_811), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx12f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x6_ASAP7_75t_SL g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx3_ASAP7_75t_L g843 ( .A(n_111), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_111), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NOR2x1_ASAP7_75t_L g851 ( .A(n_114), .B(n_116), .Y(n_851) );
AND2x6_ASAP7_75t_SL g826 ( .A(n_115), .B(n_827), .Y(n_826) );
AND3x2_ASAP7_75t_L g839 ( .A(n_115), .B(n_801), .C(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_802), .B(n_809), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_119), .B(n_810), .Y(n_809) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_472), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g120 ( .A(n_121), .B(n_467), .Y(n_120) );
NAND2x1p5_ASAP7_75t_L g121 ( .A(n_122), .B(n_411), .Y(n_121) );
NOR3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_329), .C(n_366), .Y(n_122) );
NAND4xp75_ASAP7_75t_L g123 ( .A(n_124), .B(n_249), .C(n_283), .D(n_313), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI32xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_171), .A3(n_221), .B1(n_230), .B2(n_244), .Y(n_125) );
OR2x2_ASAP7_75t_L g230 ( .A(n_126), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g440 ( .A1(n_127), .A2(n_441), .B(n_443), .Y(n_440) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_156), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_128), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g312 ( .A(n_128), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g407 ( .A(n_128), .B(n_223), .Y(n_407) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx2_ASAP7_75t_L g256 ( .A(n_129), .Y(n_256) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_129) );
OAI21x1_ASAP7_75t_L g289 ( .A1(n_130), .A2(n_134), .B(n_154), .Y(n_289) );
INVx2_ASAP7_75t_SL g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g155 ( .A(n_131), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_131), .B(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g218 ( .A(n_131), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_131), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_131), .B(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g483 ( .A(n_131), .Y(n_483) );
AND2x4_ASAP7_75t_SL g562 ( .A(n_131), .B(n_493), .Y(n_562) );
INVx1_ASAP7_75t_SL g565 ( .A(n_131), .Y(n_565) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_144), .B(n_150), .Y(n_134) );
O2A1O1Ixp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_137), .B(n_140), .C(n_142), .Y(n_135) );
INVx4_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g200 ( .A(n_138), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_138), .A2(n_167), .B1(n_545), .B2(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_139), .Y(n_141) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
INVx1_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
INVx1_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVx1_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
INVx2_ASAP7_75t_L g237 ( .A(n_139), .Y(n_237) );
INVx1_ASAP7_75t_L g239 ( .A(n_139), .Y(n_239) );
INVx3_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVx1_ASAP7_75t_L g504 ( .A(n_141), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_141), .A2(n_568), .B(n_569), .Y(n_567) );
INVx6_ASAP7_75t_L g149 ( .A(n_142), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_142), .A2(n_491), .B(n_492), .Y(n_490) );
O2A1O1Ixp5_ASAP7_75t_L g618 ( .A1(n_142), .A2(n_181), .B(n_619), .C(n_620), .Y(n_618) );
BUFx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g164 ( .A(n_143), .Y(n_164) );
INVx1_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
INVx1_ASAP7_75t_L g489 ( .A(n_143), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_149), .Y(n_144) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_149), .A2(n_160), .B1(n_162), .B2(n_165), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g178 ( .A1(n_149), .A2(n_162), .B1(n_179), .B2(n_183), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_149), .A2(n_196), .B1(n_201), .B2(n_202), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_149), .A2(n_162), .B1(n_212), .B2(n_215), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_149), .A2(n_202), .B1(n_226), .B2(n_227), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_149), .A2(n_235), .B1(n_238), .B2(n_240), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_149), .A2(n_162), .B1(n_274), .B2(n_275), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_149), .A2(n_162), .B1(n_510), .B2(n_512), .Y(n_509) );
INVx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_SL g241 ( .A(n_151), .Y(n_241) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx10_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
BUFx10_ASAP7_75t_L g493 ( .A(n_152), .Y(n_493) );
INVx2_ASAP7_75t_L g168 ( .A(n_155), .Y(n_168) );
INVx2_ASAP7_75t_L g280 ( .A(n_156), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_156), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_157), .Y(n_267) );
INVx1_ASAP7_75t_L g311 ( .A(n_157), .Y(n_311) );
AND2x2_ASAP7_75t_L g355 ( .A(n_157), .B(n_289), .Y(n_355) );
OR2x2_ASAP7_75t_L g409 ( .A(n_157), .B(n_233), .Y(n_409) );
AO31x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .A3(n_168), .B(n_169), .Y(n_157) );
INVx2_ASAP7_75t_L g177 ( .A(n_158), .Y(n_177) );
AO31x2_ASAP7_75t_L g194 ( .A1(n_158), .A2(n_195), .A3(n_204), .B(n_206), .Y(n_194) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_158), .A2(n_211), .A3(n_218), .B(n_219), .Y(n_210) );
AO31x2_ASAP7_75t_L g508 ( .A1(n_158), .A2(n_187), .A3(n_509), .B(n_513), .Y(n_508) );
INVx2_ASAP7_75t_L g532 ( .A(n_161), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_162), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g533 ( .A(n_163), .Y(n_533) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g559 ( .A(n_164), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_167), .A2(n_499), .B(n_500), .Y(n_498) );
INVx2_ASAP7_75t_L g511 ( .A(n_167), .Y(n_511) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_172), .A2(n_335), .B1(n_427), .B2(n_429), .Y(n_426) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_192), .Y(n_172) );
INVx4_ASAP7_75t_L g252 ( .A(n_173), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_173), .A2(n_232), .B1(n_264), .B2(n_266), .Y(n_263) );
OR2x2_ASAP7_75t_L g269 ( .A(n_173), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g388 ( .A(n_173), .B(n_287), .Y(n_388) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g308 ( .A(n_174), .B(n_193), .Y(n_308) );
AND2x2_ASAP7_75t_L g399 ( .A(n_174), .B(n_271), .Y(n_399) );
AND2x2_ASAP7_75t_L g454 ( .A(n_174), .B(n_210), .Y(n_454) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
AND2x4_ASAP7_75t_L g375 ( .A(n_175), .B(n_271), .Y(n_375) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .A3(n_185), .B(n_189), .Y(n_175) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_176), .A2(n_204), .A3(n_225), .B(n_228), .Y(n_224) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp67_ASAP7_75t_SL g538 ( .A(n_177), .B(n_186), .Y(n_538) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_185), .A2(n_241), .A3(n_273), .B(n_276), .Y(n_272) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_SL g206 ( .A(n_187), .B(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_187), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g191 ( .A(n_188), .Y(n_191) );
INVx2_ASAP7_75t_L g205 ( .A(n_188), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_191), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g507 ( .A(n_191), .Y(n_507) );
INVx2_ASAP7_75t_L g534 ( .A(n_191), .Y(n_534) );
NAND2x1_ASAP7_75t_L g251 ( .A(n_192), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_192), .B(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_208), .Y(n_192) );
INVx2_ASAP7_75t_L g246 ( .A(n_193), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_193), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g294 ( .A(n_193), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_193), .B(n_296), .Y(n_321) );
AND2x2_ASAP7_75t_L g324 ( .A(n_193), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g384 ( .A(n_193), .Y(n_384) );
INVx4_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_194), .B(n_209), .Y(n_262) );
BUFx2_ASAP7_75t_L g300 ( .A(n_194), .Y(n_300) );
AND2x2_ASAP7_75t_L g349 ( .A(n_194), .B(n_210), .Y(n_349) );
AND2x2_ASAP7_75t_L g391 ( .A(n_194), .B(n_272), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_194), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
INVx1_ASAP7_75t_L g505 ( .A(n_203), .Y(n_505) );
BUFx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_205), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_210), .B(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g302 ( .A(n_210), .B(n_272), .Y(n_302) );
INVx1_ASAP7_75t_L g325 ( .A(n_210), .Y(n_325) );
INVx2_ASAP7_75t_L g345 ( .A(n_210), .Y(n_345) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_210), .Y(n_390) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AO31x2_ASAP7_75t_L g233 ( .A1(n_218), .A2(n_234), .A3(n_241), .B(n_242), .Y(n_233) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g309 ( .A(n_222), .B(n_310), .Y(n_309) );
NOR2x1p5_ASAP7_75t_L g415 ( .A(n_222), .B(n_409), .Y(n_415) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x4_ASAP7_75t_L g232 ( .A(n_223), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g265 ( .A(n_223), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_223), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_223), .B(n_341), .Y(n_340) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g257 ( .A(n_224), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g315 ( .A(n_224), .B(n_233), .Y(n_315) );
BUFx2_ASAP7_75t_L g428 ( .A(n_224), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_230), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g466 ( .A(n_230), .Y(n_466) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g402 ( .A(n_232), .Y(n_402) );
AND2x4_ASAP7_75t_L g425 ( .A(n_232), .B(n_355), .Y(n_425) );
AND2x2_ASAP7_75t_L g449 ( .A(n_232), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g258 ( .A(n_233), .Y(n_258) );
BUFx2_ASAP7_75t_L g282 ( .A(n_233), .Y(n_282) );
INVx1_ASAP7_75t_L g338 ( .A(n_233), .Y(n_338) );
OR2x2_ASAP7_75t_L g460 ( .A(n_233), .B(n_317), .Y(n_460) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_237), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g560 ( .A(n_239), .Y(n_560) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g306 ( .A(n_246), .Y(n_306) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_247), .Y(n_323) );
INVx1_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g268 ( .A(n_248), .Y(n_268) );
OR2x2_ASAP7_75t_L g305 ( .A(n_248), .B(n_297), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B(n_259), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_254), .A2(n_348), .B1(n_350), .B2(n_353), .Y(n_347) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
OR2x2_ASAP7_75t_L g393 ( .A(n_256), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g401 ( .A(n_256), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_256), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g376 ( .A(n_257), .B(n_355), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .B1(n_269), .B2(n_278), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g328 ( .A(n_262), .Y(n_328) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x4_ASAP7_75t_L g286 ( .A(n_265), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g354 ( .A(n_265), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g363 ( .A(n_265), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_265), .B(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_266), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
AND2x2_ASAP7_75t_L g351 ( .A(n_268), .B(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g365 ( .A(n_268), .Y(n_365) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g297 ( .A(n_272), .Y(n_297) );
AND2x4_ASAP7_75t_L g344 ( .A(n_272), .B(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_272), .Y(n_360) );
INVx1_ASAP7_75t_L g424 ( .A(n_272), .Y(n_424) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x4_ASAP7_75t_L g316 ( .A(n_280), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g333 ( .A(n_280), .Y(n_333) );
INVx1_ASAP7_75t_L g291 ( .A(n_282), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_292), .B1(n_303), .B2(n_309), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_286), .B(n_290), .Y(n_285) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_SL g341 ( .A(n_288), .Y(n_341) );
INVx1_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_298), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_294), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g446 ( .A(n_295), .Y(n_446) );
INVx1_ASAP7_75t_L g465 ( .A(n_295), .Y(n_465) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_299), .B(n_365), .Y(n_442) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g458 ( .A(n_300), .Y(n_458) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_307), .Y(n_303) );
INVx2_ASAP7_75t_L g396 ( .A(n_304), .Y(n_396) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx2_ASAP7_75t_L g385 ( .A(n_305), .Y(n_385) );
AND2x4_ASAP7_75t_L g387 ( .A(n_306), .B(n_344), .Y(n_387) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_310), .A2(n_456), .B1(n_459), .B2(n_461), .Y(n_455) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g380 ( .A(n_311), .Y(n_380) );
INVx1_ASAP7_75t_L g334 ( .A(n_312), .Y(n_334) );
AND2x4_ASAP7_75t_L g427 ( .A(n_312), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g435 ( .A(n_312), .B(n_436), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_318), .Y(n_313) );
AND2x4_ASAP7_75t_SL g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_SL g378 ( .A(n_315), .Y(n_378) );
INVx2_ASAP7_75t_L g394 ( .A(n_315), .Y(n_394) );
INVx1_ASAP7_75t_L g421 ( .A(n_316), .Y(n_421) );
AND2x2_ASAP7_75t_L g452 ( .A(n_316), .B(n_363), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_322), .C(n_326), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_323), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g364 ( .A(n_324), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_324), .B(n_399), .Y(n_432) );
INVx1_ASAP7_75t_L g352 ( .A(n_325), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_327), .B(n_391), .Y(n_417) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_346), .C(n_356), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B(n_342), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g450 ( .A(n_333), .Y(n_450) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_339), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AOI32xp33_ASAP7_75t_L g386 ( .A1(n_337), .A2(n_387), .A3(n_388), .B1(n_389), .B2(n_392), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_337), .B(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g370 ( .A(n_344), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_344), .B(n_365), .Y(n_405) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_349), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g410 ( .A(n_349), .B(n_359), .Y(n_410) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g438 ( .A(n_352), .Y(n_438) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g356 ( .A1(n_354), .A2(n_357), .B1(n_361), .B2(n_364), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_355), .B(n_363), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_357), .A2(n_415), .B1(n_452), .B2(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g453 ( .A(n_359), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_361), .A2(n_404), .B1(n_406), .B2(n_410), .Y(n_403) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g445 ( .A(n_365), .Y(n_445) );
NAND4xp25_ASAP7_75t_L g366 ( .A(n_367), .B(n_386), .C(n_395), .D(n_403), .Y(n_366) );
O2A1O1Ixp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_373), .B(n_376), .C(n_377), .Y(n_367) );
NOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g431 ( .A(n_375), .B(n_390), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_375), .B(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_382), .A2(n_420), .B1(n_422), .B2(n_425), .Y(n_419) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_387), .A2(n_392), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_400), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_R g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_410), .A2(n_427), .B1(n_464), .B2(n_466), .Y(n_463) );
NOR3x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_433), .C(n_447), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_426), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g439 ( .A(n_414), .Y(n_439) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g462 ( .A(n_424), .Y(n_462) );
INVx1_ASAP7_75t_L g436 ( .A(n_428), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_430), .A2(n_434), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g447 ( .A(n_448), .B(n_451), .C(n_455), .D(n_463), .Y(n_447) );
AND2x2_ASAP7_75t_L g461 ( .A(n_454), .B(n_462), .Y(n_461) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVxp67_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx4_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx12f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g850 ( .A(n_470), .B(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g801 ( .A(n_471), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_798), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
BUFx2_ASAP7_75t_L g815 ( .A(n_475), .Y(n_815) );
NAND2x1p5_ASAP7_75t_SL g475 ( .A(n_476), .B(n_732), .Y(n_475) );
NOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_668), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_590), .C(n_629), .D(n_658), .Y(n_477) );
O2A1O1Ixp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_515), .B(n_522), .C(n_574), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_495), .Y(n_479) );
INVx2_ASAP7_75t_L g518 ( .A(n_480), .Y(n_518) );
AND2x2_ASAP7_75t_L g656 ( .A(n_480), .B(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_480), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_480), .B(n_576), .Y(n_751) );
OR2x2_ASAP7_75t_L g787 ( .A(n_480), .B(n_703), .Y(n_787) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g684 ( .A(n_481), .B(n_496), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g710 ( .A(n_481), .B(n_520), .Y(n_710) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g645 ( .A(n_482), .Y(n_645) );
OAI21x1_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B(n_494), .Y(n_482) );
OAI21x1_ASAP7_75t_L g496 ( .A1(n_483), .A2(n_497), .B(n_506), .Y(n_496) );
OAI21x1_ASAP7_75t_L g578 ( .A1(n_483), .A2(n_484), .B(n_494), .Y(n_578) );
OA21x2_ASAP7_75t_L g613 ( .A1(n_483), .A2(n_497), .B(n_506), .Y(n_613) );
OAI21x1_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_490), .B(n_493), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_488), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_488), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_488), .A2(n_554), .B(n_555), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_488), .A2(n_571), .B(n_572), .Y(n_570) );
BUFx4f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI21x1_ASAP7_75t_L g497 ( .A1(n_493), .A2(n_498), .B(n_501), .Y(n_497) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_493), .A2(n_526), .B(n_529), .Y(n_525) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_493), .A2(n_567), .B(n_570), .Y(n_566) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_493), .A2(n_618), .B(n_621), .Y(n_617) );
AND2x2_ASAP7_75t_L g584 ( .A(n_495), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_495), .B(n_614), .Y(n_628) );
AND2x2_ASAP7_75t_L g636 ( .A(n_495), .B(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_495), .Y(n_659) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_508), .Y(n_495) );
INVx1_ASAP7_75t_L g520 ( .A(n_496), .Y(n_520) );
INVx1_ASAP7_75t_L g576 ( .A(n_496), .Y(n_576) );
AND2x2_ASAP7_75t_L g646 ( .A(n_496), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g707 ( .A(n_496), .B(n_615), .Y(n_707) );
AOI21x1_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g521 ( .A(n_508), .Y(n_521) );
AND2x2_ASAP7_75t_L g577 ( .A(n_508), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_508), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_508), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g690 ( .A(n_508), .B(n_645), .Y(n_690) );
OR2x2_ASAP7_75t_L g703 ( .A(n_508), .B(n_613), .Y(n_703) );
OR2x2_ASAP7_75t_L g713 ( .A(n_508), .B(n_578), .Y(n_713) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_518), .B(n_729), .Y(n_775) );
INVx1_ASAP7_75t_L g631 ( .A(n_519), .Y(n_631) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_L g715 ( .A(n_521), .B(n_578), .Y(n_715) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_548), .Y(n_522) );
AND2x2_ASAP7_75t_L g588 ( .A(n_523), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g650 ( .A(n_523), .Y(n_650) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_536), .Y(n_523) );
BUFx2_ASAP7_75t_L g757 ( .A(n_524), .Y(n_757) );
OAI21xp33_ASAP7_75t_SL g524 ( .A1(n_525), .A2(n_534), .B(n_535), .Y(n_524) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_525), .A2(n_534), .B(n_535), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B(n_533), .Y(n_529) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_534), .A2(n_617), .B(n_624), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g647 ( .A1(n_534), .A2(n_617), .B(n_624), .Y(n_647) );
AND2x2_ASAP7_75t_L g596 ( .A(n_536), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g582 ( .A(n_537), .B(n_564), .Y(n_582) );
INVx2_ASAP7_75t_L g608 ( .A(n_537), .Y(n_608) );
AOI21x1_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B(n_547), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
AND2x2_ASAP7_75t_L g754 ( .A(n_548), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_563), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g581 ( .A(n_550), .Y(n_581) );
BUFx2_ASAP7_75t_L g589 ( .A(n_550), .Y(n_589) );
OR2x2_ASAP7_75t_L g593 ( .A(n_550), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g653 ( .A(n_550), .B(n_597), .Y(n_653) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
OAI21x1_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_556), .B(n_562), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_559), .B1(n_560), .B2(n_561), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_558), .A2(n_622), .B(n_623), .Y(n_621) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g640 ( .A(n_563), .Y(n_640) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_563), .Y(n_654) );
INVx2_ASAP7_75t_L g679 ( .A(n_563), .Y(n_679) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g594 ( .A(n_564), .Y(n_594) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_566), .B(n_573), .Y(n_564) );
OAI22xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_579), .B1(n_583), .B2(n_587), .Y(n_574) );
INVx1_ASAP7_75t_L g664 ( .A(n_575), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx2_ASAP7_75t_L g675 ( .A(n_576), .Y(n_675) );
AND2x2_ASAP7_75t_L g692 ( .A(n_577), .B(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_577), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g586 ( .A(n_578), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_579), .B(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_580), .B(n_596), .Y(n_687) );
AND2x2_ASAP7_75t_L g695 ( .A(n_580), .B(n_661), .Y(n_695) );
AND2x2_ASAP7_75t_L g771 ( .A(n_580), .B(n_718), .Y(n_771) );
BUFx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g606 ( .A(n_581), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g627 ( .A(n_581), .B(n_597), .Y(n_627) );
OR2x2_ASAP7_75t_L g639 ( .A(n_581), .B(n_640), .Y(n_639) );
NAND2x1_ASAP7_75t_L g673 ( .A(n_581), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g678 ( .A(n_581), .Y(n_678) );
INVx2_ASAP7_75t_L g672 ( .A(n_582), .Y(n_672) );
AND2x2_ASAP7_75t_L g698 ( .A(n_582), .B(n_662), .Y(n_698) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_585), .Y(n_634) );
INVx1_ASAP7_75t_L g701 ( .A(n_585), .Y(n_701) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g685 ( .A(n_586), .B(n_615), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_587), .A2(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g758 ( .A(n_589), .B(n_698), .Y(n_758) );
INVx1_ASAP7_75t_L g794 ( .A(n_589), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_599), .B(n_603), .Y(n_590) );
AOI322xp5_ASAP7_75t_L g742 ( .A1(n_591), .A2(n_638), .A3(n_743), .B1(n_744), .B2(n_745), .C1(n_746), .C2(n_749), .Y(n_742) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
NOR3xp33_ASAP7_75t_L g730 ( .A(n_593), .B(n_595), .C(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g609 ( .A(n_594), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g738 ( .A(n_594), .B(n_739), .Y(n_738) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_594), .Y(n_790) );
OR2x2_ASAP7_75t_L g686 ( .A(n_595), .B(n_639), .Y(n_686) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g674 ( .A(n_597), .Y(n_674) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g610 ( .A(n_598), .Y(n_610) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_SL g735 ( .A(n_600), .Y(n_735) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g706 ( .A(n_601), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g769 ( .A(n_602), .B(n_729), .Y(n_769) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_611), .B(n_625), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_605), .B(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
AND2x2_ASAP7_75t_L g661 ( .A(n_607), .B(n_662), .Y(n_661) );
AND3x2_ASAP7_75t_L g705 ( .A(n_607), .B(n_609), .C(n_678), .Y(n_705) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g667 ( .A(n_608), .Y(n_667) );
AND2x2_ASAP7_75t_L g718 ( .A(n_608), .B(n_679), .Y(n_718) );
INVx2_ASAP7_75t_L g741 ( .A(n_608), .Y(n_741) );
AND2x2_ASAP7_75t_L g745 ( .A(n_609), .B(n_741), .Y(n_745) );
INVx2_ASAP7_75t_L g662 ( .A(n_610), .Y(n_662) );
OR2x2_ASAP7_75t_L g796 ( .A(n_610), .B(n_679), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_611), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g748 ( .A(n_612), .Y(n_748) );
AND2x2_ASAP7_75t_L g657 ( .A(n_613), .B(n_647), .Y(n_657) );
AND2x2_ASAP7_75t_L g693 ( .A(n_613), .B(n_615), .Y(n_693) );
AND2x2_ASAP7_75t_L g689 ( .A(n_614), .B(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_614), .B(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g761 ( .A(n_614), .Y(n_761) );
BUFx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g632 ( .A(n_615), .Y(n_632) );
INVxp67_ASAP7_75t_SL g637 ( .A(n_615), .Y(n_637) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_615), .Y(n_683) );
INVx1_ASAP7_75t_L g729 ( .A(n_615), .Y(n_729) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_638), .B(n_641), .Y(n_629) );
OAI31xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .A3(n_633), .B(n_635), .Y(n_630) );
INVx1_ASAP7_75t_L g712 ( .A(n_632), .Y(n_712) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_633), .A2(n_642), .A3(n_671), .B1(n_675), .B2(n_676), .Y(n_670) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g663 ( .A(n_639), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_648), .B1(n_651), .B2(n_655), .Y(n_641) );
OAI22xp33_ASAP7_75t_SL g726 ( .A1(n_642), .A2(n_687), .B1(n_727), .B2(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx2_ASAP7_75t_L g784 ( .A(n_644), .Y(n_784) );
BUFx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g739 ( .A(n_647), .Y(n_739) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx3_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
AND2x2_ASAP7_75t_L g665 ( .A(n_653), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g740 ( .A(n_653), .B(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g791 ( .A(n_653), .Y(n_791) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g731 ( .A(n_657), .Y(n_731) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_664), .B2(n_665), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_660), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
AND2x2_ASAP7_75t_L g717 ( .A(n_662), .B(n_678), .Y(n_717) );
AOI211xp5_ASAP7_75t_L g722 ( .A1(n_665), .A2(n_723), .B(n_726), .C(n_730), .Y(n_722) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
HB1xp67_ASAP7_75t_L g780 ( .A(n_667), .Y(n_780) );
INVx1_ASAP7_75t_L g797 ( .A(n_667), .Y(n_797) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_669), .B(n_691), .C(n_704), .D(n_722), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_680), .Y(n_669) );
OR2x6_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_674), .B(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g779 ( .A(n_677), .B(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_680) );
NOR2xp33_ASAP7_75t_SL g681 ( .A(n_682), .B(n_685), .Y(n_681) );
BUFx2_ASAP7_75t_L g694 ( .A(n_682), .Y(n_694) );
AND2x4_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_688), .B(n_774), .Y(n_773) );
INVx3_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g743 ( .A(n_690), .B(n_729), .Y(n_743) );
O2A1O1Ixp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_694), .B(n_695), .C(n_696), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_693), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g753 ( .A(n_700), .B(n_754), .Y(n_753) );
AND2x4_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_708), .B2(n_716), .C(n_719), .Y(n_704) );
AND2x2_ASAP7_75t_L g783 ( .A(n_707), .B(n_784), .Y(n_783) );
NAND3xp33_ASAP7_75t_SL g708 ( .A(n_709), .B(n_711), .C(n_714), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OR2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_712), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_712), .B(n_748), .Y(n_778) );
INVx1_ASAP7_75t_L g721 ( .A(n_713), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_713), .Y(n_725) );
AND2x2_ASAP7_75t_L g766 ( .A(n_715), .B(n_755), .Y(n_766) );
NAND2xp33_ASAP7_75t_SL g767 ( .A(n_715), .B(n_737), .Y(n_767) );
AND2x4_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g727 ( .A(n_718), .Y(n_727) );
NOR3x1_ASAP7_75t_L g732 ( .A(n_733), .B(n_762), .C(n_781), .Y(n_732) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_742), .C(n_752), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
AND2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g755 ( .A(n_739), .Y(n_755) );
INVx2_ASAP7_75t_L g744 ( .A(n_741), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_743), .A2(n_786), .B1(n_793), .B2(n_863), .Y(n_792) );
O2A1O1Ixp5_ASAP7_75t_L g764 ( .A1(n_744), .A2(n_756), .B(n_765), .C(n_767), .Y(n_764) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AO21x1_ASAP7_75t_L g768 ( .A1(n_747), .A2(n_769), .B(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OR2x2_ASAP7_75t_L g760 ( .A(n_751), .B(n_761), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_756), .B1(n_758), .B2(n_759), .Y(n_752) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND4xp75_ASAP7_75t_L g762 ( .A(n_763), .B(n_768), .C(n_772), .D(n_776), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_779), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
NAND3xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .C(n_792), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_788), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVxp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
AND2x4_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NOR2x1p5_ASAP7_75t_SL g795 ( .A(n_796), .B(n_797), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx2_ASAP7_75t_SL g802 ( .A(n_803), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_803), .Y(n_810) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI21xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_842), .B(n_844), .Y(n_811) );
OAI21xp5_ASAP7_75t_SL g812 ( .A1(n_813), .A2(n_822), .B(n_834), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g834 ( .A1(n_814), .A2(n_815), .B1(n_816), .B2(n_817), .C(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_818), .Y(n_821) );
AO21x1_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_830), .B(n_831), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
CKINVDCx8_ASAP7_75t_R g833 ( .A(n_826), .Y(n_833) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_829), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g836 ( .A1(n_830), .A2(n_837), .B(n_841), .Y(n_836) );
INVxp67_ASAP7_75t_L g841 ( .A(n_831), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_833), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
INVx3_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx4_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
BUFx10_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
AND2x6_ASAP7_75t_L g855 ( .A(n_850), .B(n_856), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
BUFx3_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_855), .Y(n_861) );
BUFx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
endmodule