module fake_jpeg_22740_n_280 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_24),
.Y(n_54)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_65),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_27),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_22),
.B1(n_38),
.B2(n_29),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_58),
.A2(n_25),
.B(n_44),
.C(n_5),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_23),
.B1(n_18),
.B2(n_35),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_67),
.B1(n_32),
.B2(n_30),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_46),
.B1(n_39),
.B2(n_41),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_77),
.B1(n_28),
.B2(n_26),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_64),
.Y(n_95)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_66),
.B(n_79),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_23),
.B1(n_21),
.B2(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_69),
.B(n_1),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_70),
.A2(n_26),
.B1(n_20),
.B2(n_30),
.Y(n_84)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_72),
.Y(n_106)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_42),
.B(n_36),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_33),
.B(n_35),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_92),
.C(n_109),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_3),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_84),
.A2(n_85),
.B1(n_96),
.B2(n_104),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_34),
.B1(n_18),
.B2(n_33),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_27),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_34),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_SL g131 ( 
.A(n_90),
.B(n_91),
.C(n_50),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_18),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_63),
.A2(n_32),
.B(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_44),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_56),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_112),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_53),
.B(n_25),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_74),
.B1(n_68),
.B2(n_57),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_99),
.B1(n_103),
.B2(n_100),
.Y(n_156)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_128),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_68),
.B1(n_57),
.B2(n_72),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_137),
.B1(n_113),
.B2(n_131),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_92),
.C(n_80),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_95),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_123),
.B(n_91),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_90),
.A2(n_3),
.B(n_4),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_124),
.A2(n_134),
.B(n_140),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_109),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_74),
.B1(n_73),
.B2(n_51),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_135),
.B1(n_139),
.B2(n_105),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_3),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_141),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_94),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_50),
.B1(n_17),
.B2(n_10),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_6),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_93),
.Y(n_168)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_152),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_157),
.C(n_163),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_151),
.B(n_172),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_101),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_162),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_119),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_91),
.B1(n_103),
.B2(n_81),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_154),
.B(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_158),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_157),
.B1(n_129),
.B2(n_132),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_119),
.A2(n_115),
.B1(n_130),
.B2(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_160),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_81),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_87),
.B(n_89),
.Y(n_182)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_168),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_123),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_100),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_93),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_124),
.A2(n_99),
.B(n_102),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_179),
.B1(n_171),
.B2(n_169),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_127),
.B1(n_126),
.B2(n_102),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_86),
.B(n_82),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_185),
.B(n_189),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_164),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_193),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_89),
.B(n_98),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_187),
.B(n_190),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_151),
.C(n_146),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_147),
.A2(n_97),
.B(n_88),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_197),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_204),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_162),
.B1(n_145),
.B2(n_154),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_199),
.A2(n_200),
.B1(n_181),
.B2(n_188),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_151),
.B1(n_148),
.B2(n_152),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_209),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_144),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_208),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_211),
.A2(n_216),
.B1(n_196),
.B2(n_190),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_214),
.C(n_9),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_215),
.B(n_198),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_144),
.C(n_158),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_167),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_192),
.A2(n_160),
.B1(n_117),
.B2(n_136),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_217),
.A2(n_185),
.B1(n_191),
.B2(n_182),
.Y(n_230)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_173),
.B1(n_174),
.B2(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_180),
.B(n_195),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_229),
.B(n_210),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_174),
.B1(n_179),
.B2(n_176),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_228),
.B1(n_234),
.B2(n_230),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_207),
.A2(n_186),
.B1(n_195),
.B2(n_178),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_217),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_230),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_206),
.A2(n_181),
.B1(n_178),
.B2(n_190),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_214),
.C(n_212),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_234)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_241),
.C(n_244),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_246),
.B(n_247),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_200),
.C(n_203),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_242),
.A2(n_232),
.B1(n_234),
.B2(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_203),
.B1(n_215),
.B2(n_218),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_220),
.B1(n_228),
.B2(n_222),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_208),
.C(n_202),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_221),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_241),
.B1(n_11),
.B2(n_12),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_229),
.C(n_223),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_243),
.B(n_204),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_255),
.A2(n_257),
.B(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_235),
.Y(n_259)
);

OAI31xp33_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_232),
.A3(n_205),
.B(n_12),
.Y(n_257)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_258),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_248),
.A2(n_246),
.B1(n_238),
.B2(n_236),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_264),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_249),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_237),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_258),
.A2(n_254),
.B(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_266),
.B(n_261),
.Y(n_270)
);

NOR4xp25_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_257),
.C(n_253),
.D(n_13),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_255),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_273),
.B(n_268),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_250),
.C(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_12),
.C(n_13),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_275),
.A2(n_276),
.B(n_9),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_277),
.A2(n_278),
.B(n_14),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_14),
.Y(n_280)
);


endmodule