module fake_netlist_6_4699_n_461 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_461);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_461;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_209;
wire n_367;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_350;
wire n_392;
wire n_442;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_443;
wire n_246;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_389;
wire n_415;
wire n_230;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_372;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_375;
wire n_338;
wire n_360;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_371;
wire n_189;
wire n_405;
wire n_213;
wire n_294;
wire n_302;
wire n_380;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_397;
wire n_155;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_381;
wire n_236;
wire n_172;
wire n_270;
wire n_239;
wire n_414;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_460;
wire n_417;
wire n_446;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_293;
wire n_334;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_456;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_356;
wire n_166;
wire n_184;
wire n_216;
wire n_455;
wire n_363;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_152;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_406;
wire n_204;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_292;
wire n_164;
wire n_307;
wire n_433;
wire n_291;
wire n_219;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_282;
wire n_436;
wire n_211;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_311;
wire n_403;
wire n_253;
wire n_136;
wire n_249;
wire n_201;
wire n_386;
wire n_159;
wire n_157;
wire n_162;
wire n_241;
wire n_275;
wire n_276;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_277;
wire n_418;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_328;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_288;
wire n_427;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_187;
wire n_361;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_37),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_42),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVxp67_ASAP7_75t_SL g136 ( 
.A(n_17),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_50),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_126),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_44),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_38),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_27),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_46),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_71),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_14),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_108),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_1),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_56),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_33),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_40),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_48),
.Y(n_158)
);

INVxp33_ASAP7_75t_SL g159 ( 
.A(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_23),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_43),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_77),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

INVxp33_ASAP7_75t_SL g166 ( 
.A(n_107),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_73),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_62),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_103),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_4),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_32),
.Y(n_176)
);

NOR2xp67_ASAP7_75t_L g177 ( 
.A(n_21),
.B(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_0),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g181 ( 
.A(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_78),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_53),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_102),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_2),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_61),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_65),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_49),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_10),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_2),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_64),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_93),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_110),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_22),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_52),
.Y(n_198)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_87),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_129),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g201 ( 
.A(n_25),
.Y(n_201)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_57),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_101),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_51),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_59),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_131),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_143),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_133),
.B(n_0),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_139),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_154),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_141),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_161),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_133),
.B(n_1),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_176),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_R g226 ( 
.A(n_138),
.B(n_12),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_138),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_132),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_196),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_143),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_134),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_134),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

NAND2x1p5_ASAP7_75t_L g237 ( 
.A(n_142),
.B(n_18),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_148),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_135),
.B(n_3),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_166),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_148),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_230),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_163),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_146),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_140),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_140),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_168),
.Y(n_261)
);

AND2x6_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_190),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_168),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_222),
.B(n_136),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_209),
.A2(n_153),
.B1(n_193),
.B2(n_175),
.Y(n_267)
);

AND2x4_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_228),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_223),
.Y(n_270)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_218),
.B(n_162),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_218),
.Y(n_273)
);

INVx4_ASAP7_75t_SL g274 ( 
.A(n_236),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_232),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_188),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_159),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_220),
.B(n_159),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_244),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_242),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_199),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_219),
.Y(n_286)
);

NAND2x1_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_190),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_194),
.B1(n_197),
.B2(n_206),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_259),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_278),
.A2(n_194),
.B(n_197),
.C(n_206),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_241),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_255),
.A2(n_200),
.B(n_201),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_191),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_202),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_278),
.A2(n_182),
.B1(n_151),
.B2(n_152),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_247),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_225),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_SL g306 ( 
.A(n_279),
.B(n_239),
.C(n_184),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

AOI211xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_177),
.B(n_155),
.C(n_156),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_203),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_280),
.A2(n_181),
.B1(n_237),
.B2(n_233),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_268),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_150),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_248),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_157),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_240),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_SL g324 ( 
.A(n_277),
.B(n_205),
.C(n_204),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_270),
.B(n_158),
.Y(n_325)
);

BUFx8_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_308),
.Y(n_327)
);

O2A1O1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_260),
.B(n_160),
.C(n_185),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_261),
.Y(n_329)
);

AND2x4_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_252),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_312),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_286),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_290),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_SL g334 ( 
.A1(n_292),
.A2(n_245),
.B(n_181),
.Y(n_334)
);

OA21x2_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_260),
.B(n_164),
.Y(n_335)
);

O2A1O1Ixp5_ASAP7_75t_SL g336 ( 
.A1(n_309),
.A2(n_189),
.B(n_169),
.C(n_170),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_297),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_252),
.B(n_267),
.C(n_167),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_317),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_258),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_299),
.A2(n_192),
.B(n_173),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_172),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_314),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_297),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_314),
.A2(n_245),
.B1(n_262),
.B2(n_174),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_299),
.B(n_262),
.Y(n_350)
);

A2O1A1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_288),
.A2(n_267),
.B(n_198),
.C(n_195),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_245),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_321),
.A2(n_315),
.B1(n_325),
.B2(n_306),
.Y(n_353)
);

INVx4_ASAP7_75t_SL g354 ( 
.A(n_320),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_293),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_347),
.A2(n_178),
.B1(n_180),
.B2(n_183),
.Y(n_359)
);

AOI222xp33_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_310),
.B1(n_298),
.B2(n_307),
.C1(n_304),
.C2(n_303),
.Y(n_360)
);

OAI22xp33_ASAP7_75t_L g361 ( 
.A1(n_344),
.A2(n_300),
.B1(n_289),
.B2(n_284),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_294),
.B(n_313),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_335),
.A2(n_248),
.B1(n_287),
.B2(n_289),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_352),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_333),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_291),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_337),
.Y(n_367)
);

A2O1A1Ixp33_ASAP7_75t_L g368 ( 
.A1(n_351),
.A2(n_328),
.B(n_353),
.C(n_347),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_274),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_327),
.B(n_338),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_3),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_338),
.B(n_274),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_335),
.A2(n_248),
.B1(n_8),
.B2(n_9),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_7),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_356),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_330),
.B(n_19),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_354),
.B(n_20),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_345),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

OR2x6_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_341),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_343),
.Y(n_385)
);

BUFx4f_ASAP7_75t_SL g386 ( 
.A(n_382),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

AO21x2_ASAP7_75t_L g388 ( 
.A1(n_362),
.A2(n_349),
.B(n_334),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_379),
.Y(n_390)
);

AO21x2_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_336),
.B(n_355),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_381),
.A2(n_346),
.B1(n_11),
.B2(n_24),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_26),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_28),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_381),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g397 ( 
.A(n_386),
.B(n_380),
.Y(n_397)
);

NAND4xp25_ASAP7_75t_SL g398 ( 
.A(n_392),
.B(n_374),
.C(n_368),
.D(n_359),
.Y(n_398)
);

OAI221xp5_ASAP7_75t_SL g399 ( 
.A1(n_392),
.A2(n_374),
.B1(n_378),
.B2(n_361),
.C(n_376),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_360),
.C(n_366),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_396),
.A2(n_361),
.B1(n_377),
.B2(n_358),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

NAND3xp33_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_395),
.C(n_393),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g405 ( 
.A1(n_388),
.A2(n_377),
.B1(n_379),
.B2(n_383),
.Y(n_405)
);

AO21x2_ASAP7_75t_L g406 ( 
.A1(n_391),
.A2(n_369),
.B(n_363),
.Y(n_406)
);

OAI31xp33_ASAP7_75t_L g407 ( 
.A1(n_394),
.A2(n_372),
.A3(n_380),
.B(n_363),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_372),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_384),
.B(n_35),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_R g410 ( 
.A(n_390),
.B(n_36),
.Y(n_410)
);

NOR2x2_ASAP7_75t_L g411 ( 
.A(n_384),
.B(n_39),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_406),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_408),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_403),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_404),
.B(n_388),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_405),
.B(n_128),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_398),
.A2(n_402),
.B1(n_405),
.B2(n_407),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_41),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_401),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_403),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_397),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_411),
.Y(n_425)
);

INVx6_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_426),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_414),
.B(n_402),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_413),
.B(n_417),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_47),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_66),
.Y(n_431)
);

NOR4xp25_ASAP7_75t_SL g432 ( 
.A(n_422),
.B(n_67),
.C(n_68),
.D(n_69),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_70),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_R g434 ( 
.A(n_426),
.B(n_127),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_72),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_426),
.B(n_74),
.Y(n_437)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_419),
.B(n_75),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_415),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_415),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_420),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_436),
.B(n_421),
.Y(n_443)
);

OAI322xp33_ASAP7_75t_L g444 ( 
.A1(n_436),
.A2(n_418),
.A3(n_424),
.B1(n_412),
.B2(n_416),
.C1(n_421),
.C2(n_83),
.Y(n_444)
);

AOI31xp33_ASAP7_75t_L g445 ( 
.A1(n_438),
.A2(n_76),
.A3(n_79),
.B(n_80),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_440),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_441),
.Y(n_447)
);

NOR3xp33_ASAP7_75t_SL g448 ( 
.A(n_444),
.B(n_431),
.C(n_437),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_447),
.B(n_446),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_442),
.C(n_443),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_433),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_449),
.A2(n_434),
.B1(n_427),
.B2(n_430),
.Y(n_452)
);

AOI221xp5_ASAP7_75t_SL g453 ( 
.A1(n_451),
.A2(n_445),
.B1(n_439),
.B2(n_432),
.C(n_89),
.Y(n_453)
);

AOI222xp33_ASAP7_75t_L g454 ( 
.A1(n_452),
.A2(n_125),
.B1(n_82),
.B2(n_86),
.C1(n_90),
.C2(n_91),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_453),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_454),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_456)
);

NOR4xp25_ASAP7_75t_L g457 ( 
.A(n_455),
.B(n_97),
.C(n_98),
.D(n_99),
.Y(n_457)
);

OAI221xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_456),
.B1(n_105),
.B2(n_109),
.C(n_111),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_458),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_460),
.A2(n_123),
.B(n_124),
.Y(n_461)
);


endmodule