module fake_jpeg_1720_n_206 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx10_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_SL g61 ( 
.A(n_30),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_41),
.Y(n_64)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_29),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_83),
.Y(n_85)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_1),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_64),
.Y(n_91)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_84),
.A2(n_56),
.B1(n_61),
.B2(n_76),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_79),
.A2(n_58),
.B1(n_66),
.B2(n_71),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_97),
.B1(n_80),
.B2(n_70),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_77),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_81),
.A2(n_58),
.B(n_62),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_70),
.C(n_53),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_76),
.B1(n_75),
.B2(n_55),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_84),
.B1(n_80),
.B2(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_71),
.B1(n_76),
.B2(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_104),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_103),
.Y(n_118)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_100),
.Y(n_130)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_54),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

OR2x4_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_60),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_102),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_90),
.B(n_72),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_115),
.Y(n_131)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_113),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_110),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_75),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_84),
.B1(n_53),
.B2(n_89),
.Y(n_122)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_25),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_102),
.A2(n_70),
.B1(n_53),
.B2(n_69),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_128),
.B1(n_119),
.B2(n_130),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_21),
.B1(n_28),
.B2(n_32),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_134),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_60),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_137),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_69),
.B1(n_63),
.B2(n_3),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_126),
.B1(n_8),
.B2(n_9),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_63),
.B1(n_2),
.B2(n_3),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_27),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_26),
.C(n_49),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_139),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_117),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_129),
.A2(n_105),
.B1(n_112),
.B2(n_22),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_143),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_144),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_4),
.B(n_7),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_7),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_153),
.B1(n_154),
.B2(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_12),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_15),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_18),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_33),
.B(n_34),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_127),
.B(n_19),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_159),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_140),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_156),
.B1(n_52),
.B2(n_48),
.Y(n_180)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_42),
.B1(n_43),
.B2(n_47),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_150),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_161),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_141),
.B(n_158),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_181),
.B(n_175),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_182),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_150),
.B(n_169),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_183),
.B(n_168),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_166),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_190),
.C(n_175),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_177),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_179),
.B1(n_165),
.B2(n_184),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_194),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_193),
.B(n_195),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_199),
.B(n_191),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_197),
.C(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_192),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_204),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_167),
.Y(n_206)
);


endmodule