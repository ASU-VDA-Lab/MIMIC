module fake_ibex_283_n_34 (n_7, n_11, n_3, n_1, n_5, n_4, n_2, n_0, n_9, n_6, n_8, n_10, n_34);

input n_7;
input n_11;
input n_3;
input n_1;
input n_5;
input n_4;
input n_2;
input n_0;
input n_9;
input n_6;
input n_8;
input n_10;

output n_34;



endmodule