module fake_jpeg_16395_n_215 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_33),
.B(n_40),
.Y(n_44)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_41),
.Y(n_57)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_0),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_22),
.B1(n_31),
.B2(n_20),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_21),
.B1(n_17),
.B2(n_27),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_60),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_35),
.B(n_22),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_24),
.B1(n_39),
.B2(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_32),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_62),
.Y(n_74)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_43),
.Y(n_77)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_43),
.B1(n_42),
.B2(n_29),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_75),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_35),
.B(n_18),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_27),
.C(n_42),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_80),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_22),
.B1(n_31),
.B2(n_39),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_48),
.B1(n_62),
.B2(n_50),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_76),
.Y(n_95)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_24),
.B1(n_17),
.B2(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_44),
.Y(n_85)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_82),
.B1(n_83),
.B2(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_19),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_19),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_64),
.B1(n_62),
.B2(n_50),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_93),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_69),
.B1(n_71),
.B2(n_79),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_92),
.B1(n_103),
.B2(n_82),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_52),
.B1(n_46),
.B2(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_52),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_56),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_88),
.C(n_85),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_101),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_21),
.Y(n_101)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_1),
.C(n_2),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_72),
.C(n_73),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_49),
.B1(n_23),
.B2(n_26),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_75),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_71),
.B(n_68),
.C(n_76),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_107),
.A2(n_120),
.B(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_108),
.B(n_113),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_91),
.B(n_105),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_110),
.A2(n_117),
.B(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_119),
.A2(n_90),
.B1(n_65),
.B2(n_104),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_76),
.B(n_73),
.C(n_80),
.D(n_78),
.Y(n_121)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_26),
.A3(n_49),
.B1(n_16),
.B2(n_23),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_78),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_94),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_131),
.C(n_133),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_108),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_87),
.C(n_96),
.Y(n_131)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_137),
.B(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_87),
.C(n_89),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_95),
.B(n_100),
.Y(n_137)
);

NAND2x1_ASAP7_75t_SL g138 ( 
.A(n_121),
.B(n_95),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_101),
.B(n_92),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_125),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_103),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_145),
.C(n_117),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_112),
.B1(n_106),
.B2(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_118),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_26),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_127),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_156),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_123),
.B1(n_113),
.B2(n_119),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_157),
.B1(n_139),
.B2(n_129),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_154),
.C(n_158),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_106),
.C(n_124),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_146),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_112),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_142),
.B(n_23),
.C(n_49),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_160),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_16),
.C(n_3),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_140),
.C(n_137),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_165),
.C(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_166),
.B(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_133),
.C(n_145),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_152),
.A2(n_130),
.B(n_138),
.C(n_141),
.Y(n_174)
);

OAI31xp33_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_16),
.A3(n_4),
.B(n_5),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_132),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_16),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_146),
.B1(n_153),
.B2(n_148),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_184),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_158),
.B1(n_154),
.B2(n_162),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_183),
.Y(n_194)
);

OA21x2_ASAP7_75t_SL g180 ( 
.A1(n_176),
.A2(n_16),
.B(n_3),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_6),
.B(n_7),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_4),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_187),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_196),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_163),
.C(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_164),
.C(n_173),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_167),
.C(n_169),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_186),
.C(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_187),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_194),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_181),
.B1(n_180),
.B2(n_183),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_201),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g202 ( 
.A1(n_194),
.A2(n_181),
.B(n_179),
.C(n_9),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_192),
.B(n_11),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_197),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_10),
.C(n_12),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_207),
.A2(n_202),
.B1(n_200),
.B2(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_14),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_202),
.B(n_11),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_210),
.B(n_211),
.C(n_206),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_212),
.A2(n_10),
.B(n_13),
.C(n_175),
.Y(n_214)
);


endmodule