module fake_netlist_6_1415_n_607 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_607);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_607;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_599;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_596;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_41),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_16),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_14),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_0),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_53),
.Y(n_136)
);

BUFx2_ASAP7_75t_SL g137 ( 
.A(n_23),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_0),
.Y(n_140)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_59),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_55),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_73),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_70),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_107),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_87),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_11),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_4),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_26),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_5),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_9),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_66),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_45),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_103),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_78),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_42),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_30),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_110),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_34),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_62),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_85),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_49),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_47),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_104),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_65),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_43),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_10),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_18),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_75),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_21),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_2),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_48),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_77),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_101),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_102),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_22),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_111),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_114),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_127),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_132),
.B(n_1),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_130),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_133),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_159),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_134),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_138),
.B(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_144),
.B(n_2),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_156),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_143),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_145),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_136),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_139),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_155),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_157),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_168),
.B(n_3),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_153),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_161),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

AND2x4_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_190),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_171),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_231),
.B(n_195),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_237),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_198),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_171),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_201),
.B(n_174),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_205),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_190),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_212),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_193),
.B(n_197),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_198),
.B(n_190),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_194),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_200),
.B(n_128),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_149),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_192),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_L g278 ( 
.A(n_200),
.B(n_182),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_219),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_232),
.B(n_160),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_215),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_207),
.B(n_191),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_224),
.Y(n_286)
);

AND2x2_ASAP7_75t_R g287 ( 
.A(n_229),
.B(n_3),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_238),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_249),
.A2(n_187),
.B1(n_186),
.B2(n_184),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_276),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_279),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_137),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_141),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_162),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_163),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g302 ( 
.A(n_275),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_272),
.Y(n_303)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_240),
.B(n_164),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_254),
.Y(n_306)
);

BUFx8_ASAP7_75t_SL g307 ( 
.A(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_254),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_281),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_245),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_246),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_255),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_165),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_275),
.Y(n_315)
);

AND2x2_ASAP7_75t_SL g316 ( 
.A(n_278),
.B(n_4),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_240),
.B(n_166),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_251),
.B(n_167),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_258),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_275),
.B(n_169),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_260),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

INVx4_ASAP7_75t_SL g328 ( 
.A(n_253),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

AND2x6_ASAP7_75t_L g330 ( 
.A(n_276),
.B(n_243),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

NOR2x1p5_ASAP7_75t_L g333 ( 
.A(n_261),
.B(n_170),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_277),
.B(n_172),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_269),
.B(n_264),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_262),
.B(n_249),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_252),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_173),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_262),
.B(n_175),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_271),
.B(n_176),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_257),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_247),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_252),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_248),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_265),
.B(n_182),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_266),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_282),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_248),
.Y(n_353)
);

OAI221xp5_ASAP7_75t_L g354 ( 
.A1(n_302),
.A2(n_267),
.B1(n_247),
.B2(n_286),
.C(n_270),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_248),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_306),
.A2(n_288),
.B1(n_287),
.B2(n_285),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_250),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_328),
.Y(n_359)
);

AO22x2_ASAP7_75t_L g360 ( 
.A1(n_308),
.A2(n_285),
.B1(n_6),
.B2(n_7),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

NAND2x1p5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_285),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_335),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_316),
.A2(n_182),
.B1(n_250),
.B2(n_284),
.Y(n_365)
);

OAI221xp5_ASAP7_75t_L g366 ( 
.A1(n_305),
.A2(n_182),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_366)
);

AO22x2_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_15),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_12),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_312),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_17),
.Y(n_375)
);

AO22x2_ASAP7_75t_L g376 ( 
.A1(n_290),
.A2(n_297),
.B1(n_296),
.B2(n_322),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_325),
.Y(n_380)
);

OAI221xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.C(n_25),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_351),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_318),
.Y(n_384)
);

AO22x2_ASAP7_75t_L g385 ( 
.A1(n_344),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_35),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_346),
.B(n_36),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_323),
.Y(n_388)
);

AO22x2_ASAP7_75t_L g389 ( 
.A1(n_317),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_294),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_317),
.Y(n_392)
);

AO22x2_ASAP7_75t_L g393 ( 
.A1(n_324),
.A2(n_40),
.B1(n_46),
.B2(n_50),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_51),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_333),
.Y(n_395)
);

OAI221xp5_ASAP7_75t_L g396 ( 
.A1(n_341),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.C(n_57),
.Y(n_396)
);

AO22x2_ASAP7_75t_L g397 ( 
.A1(n_326),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_293),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_340),
.B(n_71),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_320),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_336),
.B(n_74),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_340),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_338),
.B(n_83),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g406 ( 
.A1(n_326),
.A2(n_343),
.B1(n_347),
.B2(n_334),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_303),
.B(n_84),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_L g410 ( 
.A1(n_352),
.A2(n_88),
.B(n_89),
.Y(n_410)
);

NAND2xp33_ASAP7_75t_SL g411 ( 
.A(n_359),
.B(n_289),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_388),
.B(n_332),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_384),
.B(n_332),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_378),
.B(n_371),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_309),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_395),
.B(n_310),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_386),
.B(n_332),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_390),
.B(n_365),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_369),
.B(n_291),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_SL g420 ( 
.A(n_373),
.B(n_301),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_309),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_355),
.B(n_353),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_358),
.B(n_361),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_370),
.B(n_301),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_403),
.B(n_350),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_372),
.B(n_291),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_353),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_SL g428 ( 
.A(n_394),
.B(n_291),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_SL g429 ( 
.A(n_377),
.B(n_349),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_379),
.B(n_327),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_380),
.B(n_327),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_383),
.B(n_362),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_398),
.B(n_327),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_400),
.B(n_304),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_404),
.B(n_304),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g436 ( 
.A(n_382),
.B(n_350),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_401),
.B(n_304),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_410),
.B(n_90),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_363),
.B(n_93),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_SL g440 ( 
.A(n_399),
.B(n_94),
.Y(n_440)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_375),
.B(n_96),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_376),
.B(n_97),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g443 ( 
.A(n_387),
.B(n_409),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_391),
.B(n_98),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_408),
.B(n_100),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_105),
.Y(n_446)
);

NAND2xp33_ASAP7_75t_SL g447 ( 
.A(n_405),
.B(n_106),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_422),
.A2(n_357),
.B(n_407),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_442),
.A2(n_446),
.B(n_414),
.Y(n_450)
);

AO21x1_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_438),
.B(n_440),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_415),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_406),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_423),
.Y(n_454)
);

NOR4xp25_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_366),
.C(n_381),
.D(n_396),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_SL g456 ( 
.A1(n_445),
.A2(n_402),
.B(n_354),
.C(n_389),
.Y(n_456)
);

OAI22x1_ASAP7_75t_L g457 ( 
.A1(n_421),
.A2(n_413),
.B1(n_432),
.B2(n_367),
.Y(n_457)
);

CKINVDCx11_ASAP7_75t_R g458 ( 
.A(n_415),
.Y(n_458)
);

OAI21xp33_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_368),
.B(n_367),
.Y(n_459)
);

AO31x2_ASAP7_75t_L g460 ( 
.A1(n_443),
.A2(n_385),
.A3(n_393),
.B(n_397),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_424),
.A2(n_385),
.B(n_393),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_428),
.A2(n_389),
.B(n_397),
.C(n_356),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_417),
.A2(n_360),
.B(n_109),
.Y(n_463)
);

AOI21x1_ASAP7_75t_SL g464 ( 
.A1(n_441),
.A2(n_360),
.B(n_112),
.Y(n_464)
);

AND3x2_ASAP7_75t_L g465 ( 
.A(n_425),
.B(n_108),
.C(n_113),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_419),
.B(n_115),
.Y(n_467)
);

AOI21x1_ASAP7_75t_L g468 ( 
.A1(n_426),
.A2(n_116),
.B(n_118),
.Y(n_468)
);

AOI21x1_ASAP7_75t_L g469 ( 
.A1(n_439),
.A2(n_119),
.B(n_122),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_124),
.Y(n_470)
);

NAND2x1p5_ASAP7_75t_L g471 ( 
.A(n_430),
.B(n_125),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_444),
.A2(n_433),
.B(n_435),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_416),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

AOI22x1_ASAP7_75t_L g475 ( 
.A1(n_457),
.A2(n_447),
.B1(n_429),
.B2(n_420),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_454),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_473),
.A2(n_431),
.B1(n_434),
.B2(n_470),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_452),
.B(n_467),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_459),
.A2(n_450),
.B(n_462),
.C(n_463),
.Y(n_479)
);

NAND2x1p5_ASAP7_75t_L g480 ( 
.A(n_452),
.B(n_467),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_459),
.C(n_456),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_468),
.B(n_469),
.Y(n_482)
);

OAI21x1_ASAP7_75t_L g483 ( 
.A1(n_472),
.A2(n_451),
.B(n_453),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_448),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_449),
.Y(n_485)
);

CKINVDCx6p67_ASAP7_75t_R g486 ( 
.A(n_465),
.Y(n_486)
);

AO21x2_ASAP7_75t_L g487 ( 
.A1(n_455),
.A2(n_461),
.B(n_449),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_471),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_455),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_460),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_448),
.Y(n_491)
);

A2O1A1Ixp33_ASAP7_75t_L g492 ( 
.A1(n_459),
.A2(n_436),
.B(n_371),
.C(n_450),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_458),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_454),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_458),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_448),
.B(n_292),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_478),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_496),
.B(n_484),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_494),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_484),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_478),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

AO31x2_ASAP7_75t_L g506 ( 
.A1(n_485),
.A2(n_492),
.A3(n_479),
.B(n_491),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_495),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_489),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_489),
.B(n_481),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_483),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_479),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

CKINVDCx8_ASAP7_75t_R g513 ( 
.A(n_478),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_487),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_480),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_482),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_480),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_493),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_474),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_493),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_R g523 ( 
.A(n_498),
.B(n_486),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_520),
.Y(n_524)
);

AND2x4_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_488),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_R g526 ( 
.A(n_518),
.B(n_486),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_477),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_475),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_503),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_520),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_517),
.B(n_519),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_497),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_497),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_505),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_497),
.B(n_504),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_500),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_R g537 ( 
.A(n_518),
.B(n_515),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_522),
.Y(n_538)
);

OR2x6_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_519),
.Y(n_539)
);

BUFx10_ASAP7_75t_L g540 ( 
.A(n_521),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_504),
.B(n_522),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_499),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_513),
.B(n_504),
.Y(n_543)
);

CKINVDCx8_ASAP7_75t_R g544 ( 
.A(n_504),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_504),
.B(n_513),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_534),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_536),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_542),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_538),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_527),
.A2(n_511),
.B1(n_508),
.B2(n_512),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_511),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_533),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_528),
.B(n_510),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_505),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_541),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_506),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_512),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_528),
.B(n_506),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_527),
.B(n_506),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_546),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_551),
.B(n_539),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_553),
.B(n_543),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_557),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_547),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_551),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_514),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_554),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_561),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_555),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_552),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_562),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_565),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_557),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_567),
.B(n_558),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_572),
.B(n_540),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_572),
.A2(n_563),
.B1(n_523),
.B2(n_537),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_571),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_575),
.B(n_560),
.Y(n_579)
);

INVxp33_ASAP7_75t_SL g580 ( 
.A(n_574),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_578),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_576),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_579),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_577),
.B(n_564),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_580),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_581),
.Y(n_586)
);

AOI221xp5_ASAP7_75t_L g587 ( 
.A1(n_582),
.A2(n_573),
.B1(n_569),
.B2(n_563),
.C(n_549),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_585),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_588),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_586),
.Y(n_590)
);

INVxp33_ASAP7_75t_SL g591 ( 
.A(n_589),
.Y(n_591)
);

OAI211xp5_ASAP7_75t_SL g592 ( 
.A1(n_591),
.A2(n_590),
.B(n_582),
.C(n_587),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_592),
.A2(n_584),
.B(n_583),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_593),
.B(n_531),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_594),
.B(n_530),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_595),
.Y(n_596)
);

NAND2x1p5_ASAP7_75t_L g597 ( 
.A(n_596),
.B(n_560),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_597),
.Y(n_598)
);

AOI31xp33_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_526),
.A3(n_524),
.B(n_539),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_599),
.A2(n_564),
.B1(n_570),
.B2(n_525),
.Y(n_600)
);

OAI322xp33_ASAP7_75t_L g601 ( 
.A1(n_599),
.A2(n_545),
.A3(n_524),
.B1(n_549),
.B2(n_556),
.C1(n_548),
.C2(n_555),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_600),
.A2(n_570),
.B1(n_525),
.B2(n_554),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_601),
.B(n_548),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_603),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_602),
.Y(n_605)
);

OAI221xp5_ASAP7_75t_R g606 ( 
.A1(n_604),
.A2(n_605),
.B1(n_550),
.B2(n_544),
.C(n_567),
.Y(n_606)
);

AOI211xp5_ASAP7_75t_L g607 ( 
.A1(n_606),
.A2(n_559),
.B(n_516),
.C(n_514),
.Y(n_607)
);


endmodule