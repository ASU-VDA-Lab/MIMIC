module fake_jpeg_23553_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx12_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_14),
.B(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

NAND2xp33_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_16),
.A2(n_18),
.B(n_20),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_7),
.C(n_8),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_1),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_25),
.B(n_26),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_10),
.C(n_11),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_8),
.B(n_11),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_14),
.A2(n_8),
.B1(n_10),
.B2(n_1),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_17),
.B1(n_1),
.B2(n_20),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_19),
.B1(n_13),
.B2(n_10),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.C(n_3),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_23),
.A3(n_25),
.B1(n_22),
.B2(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_2),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_36),
.C(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.C(n_36),
.Y(n_39)
);

NAND3xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_29),
.C(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);


endmodule