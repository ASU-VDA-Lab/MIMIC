module fake_jpeg_12797_n_201 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_201);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_201;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_35),
.B(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_42),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_60),
.Y(n_97)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

AND2x4_ASAP7_75t_SL g89 ( 
.A(n_78),
.B(n_24),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_22),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_75),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_89),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_100),
.B(n_71),
.C(n_61),
.D(n_80),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_78),
.B1(n_82),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_102),
.B1(n_109),
.B2(n_74),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_79),
.C(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_67),
.B1(n_74),
.B2(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_107),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_0),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_80),
.B1(n_73),
.B2(n_59),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_112),
.Y(n_133)
);

AO22x2_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_89),
.B1(n_91),
.B2(n_57),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_125),
.B1(n_101),
.B2(n_25),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_110),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_76),
.B1(n_81),
.B2(n_86),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_126),
.B(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_92),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_87),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_127),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_91),
.B1(n_72),
.B2(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_66),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_101),
.B(n_64),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_119),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_138),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_140),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_144),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_147),
.B1(n_149),
.B2(n_19),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_3),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_8),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_10),
.B(n_11),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_15),
.B(n_18),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_12),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_167),
.B(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_157),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_26),
.B(n_28),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_169),
.B(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_29),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_143),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_30),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_56),
.C(n_39),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_32),
.B(n_41),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_170),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_43),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_171),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_175),
.Y(n_184)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_136),
.B(n_140),
.Y(n_178)
);

AOI211xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_167),
.B(n_45),
.C(n_55),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_136),
.B1(n_47),
.B2(n_48),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_183),
.B1(n_159),
.B2(n_160),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_158),
.A2(n_136),
.B1(n_50),
.B2(n_53),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_186),
.Y(n_190)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_158),
.B1(n_157),
.B2(n_168),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_182),
.B1(n_183),
.B2(n_178),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_180),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_179),
.C(n_190),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_177),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_186),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_197),
.B(n_174),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_192),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_199),
.A2(n_192),
.B(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_189),
.C(n_188),
.Y(n_201)
);


endmodule