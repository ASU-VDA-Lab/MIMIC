module real_aes_6966_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_729;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
INVx1_ASAP7_75t_L g528 ( .A(n_1), .Y(n_528) );
INVx1_ASAP7_75t_L g143 ( .A(n_2), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_3), .A2(n_38), .B1(n_168), .B2(n_474), .Y(n_497) );
AOI21xp33_ASAP7_75t_L g175 ( .A1(n_4), .A2(n_159), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_5), .B(n_157), .Y(n_540) );
AND2x6_ASAP7_75t_L g136 ( .A(n_6), .B(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_7), .A2(n_246), .B(n_247), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_8), .B(n_39), .Y(n_110) );
INVx1_ASAP7_75t_L g181 ( .A(n_9), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_10), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g128 ( .A(n_11), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_12), .B(n_149), .Y(n_483) );
INVx1_ASAP7_75t_L g252 ( .A(n_13), .Y(n_252) );
INVx1_ASAP7_75t_L g522 ( .A(n_14), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_15), .B(n_124), .Y(n_511) );
AO32x2_ASAP7_75t_L g495 ( .A1(n_16), .A2(n_123), .A3(n_157), .B1(n_476), .B2(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_17), .B(n_168), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_18), .B(n_164), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_19), .B(n_124), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_20), .A2(n_49), .B1(n_168), .B2(n_474), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_21), .B(n_159), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_22), .A2(n_97), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_22), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g475 ( .A1(n_23), .A2(n_75), .B1(n_149), .B2(n_168), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_24), .B(n_168), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_25), .B(n_171), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g249 ( .A1(n_26), .A2(n_250), .B(n_251), .C(n_253), .Y(n_249) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_28), .B(n_154), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_29), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_30), .B(n_104), .Y(n_430) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_31), .A2(n_87), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_31), .Y(n_114) );
INVx1_ASAP7_75t_L g196 ( .A(n_32), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_33), .B(n_154), .Y(n_467) );
INVx2_ASAP7_75t_L g134 ( .A(n_34), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_35), .B(n_168), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_36), .B(n_154), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_37), .A2(n_136), .B(n_139), .C(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g194 ( .A(n_40), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_41), .B(n_147), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_42), .B(n_168), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_43), .A2(n_85), .B1(n_216), .B2(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_44), .B(n_168), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_45), .B(n_168), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g197 ( .A(n_46), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_47), .B(n_527), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_48), .B(n_159), .Y(n_240) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_50), .A2(n_60), .B1(n_149), .B2(n_168), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g727 ( .A1(n_51), .A2(n_728), .B1(n_729), .B2(n_732), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_51), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_52), .A2(n_139), .B1(n_149), .B2(n_192), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_53), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_54), .B(n_168), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_55), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_56), .B(n_168), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_57), .A2(n_167), .B(n_179), .C(n_180), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g229 ( .A(n_58), .Y(n_229) );
INVx1_ASAP7_75t_L g177 ( .A(n_59), .Y(n_177) );
INVx1_ASAP7_75t_L g137 ( .A(n_61), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_62), .B(n_168), .Y(n_529) );
INVx1_ASAP7_75t_L g127 ( .A(n_63), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_64), .Y(n_435) );
AO32x2_ASAP7_75t_L g471 ( .A1(n_65), .A2(n_157), .A3(n_232), .B1(n_472), .B2(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g547 ( .A(n_66), .Y(n_547) );
INVx1_ASAP7_75t_L g462 ( .A(n_67), .Y(n_462) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_68), .A2(n_103), .B1(n_431), .B2(n_439), .C1(n_738), .C2(n_743), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_68), .A2(n_112), .B1(n_428), .B2(n_429), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_68), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_SL g163 ( .A1(n_69), .A2(n_164), .B(n_165), .C(n_167), .Y(n_163) );
INVxp67_ASAP7_75t_L g166 ( .A(n_70), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_71), .B(n_149), .Y(n_463) );
INVx1_ASAP7_75t_L g438 ( .A(n_72), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_73), .Y(n_199) );
INVx1_ASAP7_75t_L g222 ( .A(n_74), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_76), .A2(n_136), .B(n_139), .C(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_77), .B(n_474), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_78), .B(n_149), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_79), .B(n_144), .Y(n_212) );
INVx2_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_81), .B(n_164), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_82), .B(n_149), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_83), .A2(n_136), .B(n_139), .C(n_142), .Y(n_138) );
OR2x2_ASAP7_75t_L g106 ( .A(n_84), .B(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g444 ( .A(n_84), .B(n_108), .Y(n_444) );
INVx2_ASAP7_75t_L g449 ( .A(n_84), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_86), .A2(n_101), .B1(n_149), .B2(n_150), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_87), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_88), .B(n_154), .Y(n_182) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_89), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_90), .A2(n_136), .B(n_139), .C(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_91), .Y(n_242) );
INVx1_ASAP7_75t_L g162 ( .A(n_92), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g248 ( .A(n_93), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_94), .B(n_144), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_95), .B(n_149), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_96), .B(n_157), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_97), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_98), .A2(n_159), .B(n_160), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_99), .B(n_438), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g440 ( .A1(n_100), .A2(n_441), .B1(n_726), .B2(n_727), .C1(n_733), .C2(n_736), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_111), .B(n_430), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g742 ( .A(n_106), .Y(n_742) );
BUFx2_ASAP7_75t_L g745 ( .A(n_106), .Y(n_745) );
NOR2x2_ASAP7_75t_L g735 ( .A(n_107), .B(n_449), .Y(n_735) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g448 ( .A(n_108), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g429 ( .A(n_112), .Y(n_429) );
XNOR2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
INVx1_ASAP7_75t_L g445 ( .A(n_116), .Y(n_445) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_116), .A2(n_446), .B1(n_451), .B2(n_737), .Y(n_736) );
NAND2x1_ASAP7_75t_L g116 ( .A(n_117), .B(n_344), .Y(n_116) );
NOR5xp2_ASAP7_75t_L g117 ( .A(n_118), .B(n_267), .C(n_299), .D(n_314), .E(n_331), .Y(n_117) );
A2O1A1Ixp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_183), .B(n_204), .C(n_255), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_155), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_120), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_120), .B(n_319), .Y(n_382) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_121), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_121), .B(n_201), .Y(n_268) );
AND2x2_ASAP7_75t_L g309 ( .A(n_121), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_121), .B(n_278), .Y(n_313) );
OR2x2_ASAP7_75t_L g350 ( .A(n_121), .B(n_189), .Y(n_350) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g188 ( .A(n_122), .B(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g258 ( .A(n_122), .Y(n_258) );
OR2x2_ASAP7_75t_L g421 ( .A(n_122), .B(n_261), .Y(n_421) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_129), .B(n_151), .Y(n_122) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_123), .A2(n_190), .B(n_198), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_123), .B(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g217 ( .A(n_123), .Y(n_217) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
AND2x2_ASAP7_75t_SL g154 ( .A(n_125), .B(n_126), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
OAI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B(n_138), .Y(n_129) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_131), .A2(n_169), .B1(n_191), .B2(n_197), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_131), .A2(n_222), .B(n_223), .Y(n_221) );
NAND2x1p5_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
AND2x4_ASAP7_75t_L g159 ( .A(n_132), .B(n_136), .Y(n_159) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g527 ( .A(n_133), .Y(n_527) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g150 ( .A(n_134), .Y(n_150) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx3_ASAP7_75t_L g145 ( .A(n_135), .Y(n_145) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_135), .Y(n_147) );
INVx1_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
INVx4_ASAP7_75t_SL g169 ( .A(n_136), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_136), .A2(n_461), .B(n_464), .Y(n_460) );
BUFx3_ASAP7_75t_L g476 ( .A(n_136), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_136), .A2(n_481), .B(n_485), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_136), .A2(n_521), .B(n_525), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_136), .A2(n_534), .B(n_537), .Y(n_533) );
INVx5_ASAP7_75t_L g161 ( .A(n_139), .Y(n_161) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
BUFx3_ASAP7_75t_L g216 ( .A(n_140), .Y(n_216) );
INVx1_ASAP7_75t_L g474 ( .A(n_140), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_146), .C(n_148), .Y(n_142) );
O2A1O1Ixp5_ASAP7_75t_SL g461 ( .A1(n_144), .A2(n_167), .B(n_462), .C(n_463), .Y(n_461) );
INVx2_ASAP7_75t_L g498 ( .A(n_144), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_144), .A2(n_535), .B(n_536), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_144), .A2(n_544), .B(n_545), .Y(n_543) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_145), .B(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_145), .B(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g472 ( .A1(n_145), .A2(n_147), .B1(n_473), .B2(n_475), .Y(n_472) );
INVx2_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
INVx4_ASAP7_75t_L g238 ( .A(n_147), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_147), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_147), .A2(n_498), .B1(n_514), .B2(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_148), .A2(n_522), .B(n_523), .C(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_153), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_153), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_154), .A2(n_245), .B(n_254), .Y(n_244) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_154), .A2(n_460), .B(n_467), .Y(n_459) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_154), .A2(n_480), .B(n_488), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g323 ( .A1(n_155), .A2(n_324), .B1(n_325), .B2(n_328), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_155), .B(n_258), .Y(n_407) );
AND2x2_ASAP7_75t_L g155 ( .A(n_156), .B(n_173), .Y(n_155) );
AND2x2_ASAP7_75t_L g203 ( .A(n_156), .B(n_189), .Y(n_203) );
AND2x2_ASAP7_75t_L g260 ( .A(n_156), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g265 ( .A(n_156), .Y(n_265) );
INVx3_ASAP7_75t_L g278 ( .A(n_156), .Y(n_278) );
OR2x2_ASAP7_75t_L g298 ( .A(n_156), .B(n_261), .Y(n_298) );
AND2x2_ASAP7_75t_L g317 ( .A(n_156), .B(n_174), .Y(n_317) );
BUFx2_ASAP7_75t_L g349 ( .A(n_156), .Y(n_349) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_170), .Y(n_156) );
INVx4_ASAP7_75t_L g172 ( .A(n_157), .Y(n_172) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_157), .A2(n_533), .B(n_540), .Y(n_532) );
BUFx2_ASAP7_75t_L g246 ( .A(n_159), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .C(n_169), .Y(n_160) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_161), .A2(n_169), .B(n_177), .C(n_178), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_161), .A2(n_169), .B(n_248), .C(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g484 ( .A(n_164), .Y(n_484) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_171), .A2(n_175), .B(n_182), .Y(n_174) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g218 ( .A(n_172), .B(n_219), .Y(n_218) );
NAND3xp33_ASAP7_75t_L g512 ( .A(n_172), .B(n_476), .C(n_513), .Y(n_512) );
AO21x1_ASAP7_75t_L g602 ( .A1(n_172), .A2(n_513), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_L g264 ( .A(n_173), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
BUFx2_ASAP7_75t_L g187 ( .A(n_174), .Y(n_187) );
INVx2_ASAP7_75t_L g202 ( .A(n_174), .Y(n_202) );
OR2x2_ASAP7_75t_L g280 ( .A(n_174), .B(n_261), .Y(n_280) );
AND2x2_ASAP7_75t_L g310 ( .A(n_174), .B(n_189), .Y(n_310) );
AND2x2_ASAP7_75t_L g327 ( .A(n_174), .B(n_258), .Y(n_327) );
AND2x2_ASAP7_75t_L g367 ( .A(n_174), .B(n_278), .Y(n_367) );
AND2x2_ASAP7_75t_SL g403 ( .A(n_174), .B(n_203), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_179), .A2(n_486), .B(n_487), .Y(n_485) );
O2A1O1Ixp5_ASAP7_75t_L g546 ( .A1(n_179), .A2(n_526), .B(n_547), .C(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp33_ASAP7_75t_SL g184 ( .A(n_185), .B(n_200), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_186), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_187), .A2(n_203), .B(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_187), .B(n_189), .Y(n_397) );
AND2x2_ASAP7_75t_L g333 ( .A(n_188), .B(n_334), .Y(n_333) );
INVx3_ASAP7_75t_L g261 ( .A(n_189), .Y(n_261) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_189), .Y(n_359) );
OAI22xp5_ASAP7_75t_SL g192 ( .A1(n_193), .A2(n_194), .B1(n_195), .B2(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g195 ( .A(n_193), .Y(n_195) );
INVx4_ASAP7_75t_L g250 ( .A(n_193), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_200), .B(n_258), .Y(n_426) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_201), .A2(n_369), .B1(n_370), .B2(n_375), .Y(n_368) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AND2x2_ASAP7_75t_L g259 ( .A(n_202), .B(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g297 ( .A(n_202), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_SL g334 ( .A(n_202), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_203), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g388 ( .A(n_203), .Y(n_388) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_230), .Y(n_205) );
INVx4_ASAP7_75t_L g274 ( .A(n_206), .Y(n_274) );
AND2x2_ASAP7_75t_L g352 ( .A(n_206), .B(n_319), .Y(n_352) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_220), .Y(n_206) );
INVx3_ASAP7_75t_L g271 ( .A(n_207), .Y(n_271) );
AND2x2_ASAP7_75t_L g285 ( .A(n_207), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g289 ( .A(n_207), .Y(n_289) );
INVx2_ASAP7_75t_L g303 ( .A(n_207), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_207), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g360 ( .A(n_207), .B(n_355), .Y(n_360) );
AND2x2_ASAP7_75t_L g425 ( .A(n_207), .B(n_395), .Y(n_425) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_210), .B(n_217), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_214), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_214), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
INVx1_ASAP7_75t_L g227 ( .A(n_217), .Y(n_227) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_217), .A2(n_520), .B(n_530), .Y(n_519) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_217), .A2(n_542), .B(n_549), .Y(n_541) );
AND2x2_ASAP7_75t_L g266 ( .A(n_220), .B(n_244), .Y(n_266) );
INVx2_ASAP7_75t_L g286 ( .A(n_220), .Y(n_286) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_227), .B(n_228), .Y(n_220) );
INVx1_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
AND2x2_ASAP7_75t_L g337 ( .A(n_230), .B(n_285), .Y(n_337) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
INVx2_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
INVx1_ASAP7_75t_L g284 ( .A(n_231), .Y(n_284) );
AND2x2_ASAP7_75t_L g302 ( .A(n_231), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_231), .B(n_286), .Y(n_340) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_241), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_239), .Y(n_235) );
AND2x2_ASAP7_75t_L g319 ( .A(n_243), .B(n_276), .Y(n_319) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g272 ( .A(n_244), .Y(n_272) );
AND2x2_ASAP7_75t_L g355 ( .A(n_244), .B(n_286), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_250), .B(n_252), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_250), .A2(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g524 ( .A(n_250), .Y(n_524) );
OAI21xp5_ASAP7_75t_SL g255 ( .A1(n_256), .A2(n_262), .B(n_266), .Y(n_255) );
INVx1_ASAP7_75t_SL g300 ( .A(n_256), .Y(n_300) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_257), .B(n_264), .Y(n_357) );
INVx1_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g306 ( .A(n_258), .B(n_261), .Y(n_306) );
AND2x2_ASAP7_75t_L g335 ( .A(n_258), .B(n_279), .Y(n_335) );
OR2x2_ASAP7_75t_L g338 ( .A(n_258), .B(n_298), .Y(n_338) );
AOI222xp33_ASAP7_75t_L g402 ( .A1(n_259), .A2(n_351), .B1(n_403), .B2(n_404), .C1(n_406), .C2(n_408), .Y(n_402) );
BUFx2_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g305 ( .A(n_264), .B(n_306), .Y(n_305) );
INVx3_ASAP7_75t_SL g322 ( .A(n_264), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_264), .B(n_316), .Y(n_376) );
AND2x2_ASAP7_75t_L g311 ( .A(n_266), .B(n_271), .Y(n_311) );
INVx1_ASAP7_75t_L g330 ( .A(n_266), .Y(n_330) );
OAI221xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_269), .B1(n_273), .B2(n_277), .C(n_281), .Y(n_267) );
OR2x2_ASAP7_75t_L g339 ( .A(n_269), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AND2x2_ASAP7_75t_L g324 ( .A(n_271), .B(n_294), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_271), .B(n_284), .Y(n_364) );
AND2x2_ASAP7_75t_L g369 ( .A(n_271), .B(n_319), .Y(n_369) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_271), .Y(n_379) );
NAND2x1_ASAP7_75t_SL g390 ( .A(n_271), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g275 ( .A(n_272), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g295 ( .A(n_272), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_272), .B(n_290), .Y(n_321) );
INVx1_ASAP7_75t_L g387 ( .A(n_272), .Y(n_387) );
INVx1_ASAP7_75t_L g362 ( .A(n_273), .Y(n_362) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g374 ( .A(n_274), .Y(n_374) );
NOR2xp67_ASAP7_75t_L g386 ( .A(n_274), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g391 ( .A(n_275), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_275), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g294 ( .A(n_276), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_276), .B(n_286), .Y(n_307) );
INVx1_ASAP7_75t_L g373 ( .A(n_276), .Y(n_373) );
INVx1_ASAP7_75t_L g394 ( .A(n_277), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI21xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_287), .B(n_296), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
AND2x2_ASAP7_75t_L g427 ( .A(n_283), .B(n_360), .Y(n_427) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g395 ( .A(n_284), .B(n_355), .Y(n_395) );
AOI32xp33_ASAP7_75t_L g308 ( .A1(n_285), .A2(n_291), .A3(n_309), .B1(n_311), .B2(n_312), .Y(n_308) );
AOI322xp5_ASAP7_75t_L g410 ( .A1(n_285), .A2(n_317), .A3(n_400), .B1(n_411), .B2(n_412), .C1(n_413), .C2(n_415), .Y(n_410) );
INVx2_ASAP7_75t_L g290 ( .A(n_286), .Y(n_290) );
INVx1_ASAP7_75t_L g400 ( .A(n_286), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_291), .B1(n_292), .B2(n_293), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_288), .B(n_294), .Y(n_343) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_289), .B(n_355), .Y(n_405) );
INVx1_ASAP7_75t_L g292 ( .A(n_290), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_290), .B(n_319), .Y(n_409) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_298), .B(n_393), .Y(n_392) );
OAI221xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_301), .B1(n_304), .B2(n_307), .C(n_308), .Y(n_299) );
OR2x2_ASAP7_75t_L g320 ( .A(n_301), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g329 ( .A(n_301), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g354 ( .A(n_302), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g358 ( .A(n_312), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_318), .B1(n_320), .B2(n_322), .C(n_323), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_316), .A2(n_347), .B1(n_351), .B2(n_352), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_317), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_317), .Y(n_422) );
INVx1_ASAP7_75t_L g416 ( .A(n_319), .Y(n_416) );
INVx1_ASAP7_75t_SL g351 ( .A(n_320), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_322), .B(n_350), .Y(n_412) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_327), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g393 ( .A(n_327), .Y(n_393) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
OAI221xp5_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_336), .B1(n_338), .B2(n_339), .C(n_341), .Y(n_331) );
NOR2xp33_ASAP7_75t_SL g332 ( .A(n_333), .B(n_335), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_333), .A2(n_351), .B1(n_397), .B2(n_398), .Y(n_396) );
CKINVDCx14_ASAP7_75t_R g336 ( .A(n_337), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_338), .A2(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NOR3xp33_ASAP7_75t_SL g344 ( .A(n_345), .B(n_377), .C(n_401), .Y(n_344) );
NAND4xp25_ASAP7_75t_L g345 ( .A(n_346), .B(n_353), .C(n_361), .D(n_368), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
INVx1_ASAP7_75t_L g424 ( .A(n_349), .Y(n_424) );
INVx3_ASAP7_75t_SL g418 ( .A(n_350), .Y(n_418) );
OR2x2_ASAP7_75t_L g423 ( .A(n_350), .B(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B1(n_358), .B2(n_360), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_355), .B(n_373), .Y(n_414) );
INVxp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_363), .B(n_365), .Y(n_361) );
INVxp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI211xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_380), .B(n_383), .C(n_396), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g411 ( .A(n_382), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_388), .B1(n_389), .B2(n_392), .C1(n_394), .C2(n_395), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND4xp25_ASAP7_75t_SL g420 ( .A(n_393), .B(n_421), .C(n_422), .D(n_423), .Y(n_420) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND3xp33_ASAP7_75t_SL g401 ( .A(n_402), .B(n_410), .C(n_419), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_419) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NOR2xp33_ASAP7_75t_SL g740 ( .A(n_435), .B(n_437), .Y(n_740) );
OA21x2_ASAP7_75t_L g744 ( .A1(n_435), .A2(n_436), .B(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_446), .B2(n_450), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g737 ( .A(n_443), .Y(n_737) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_647), .Y(n_451) );
NAND3xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_596), .C(n_638), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_505), .B(n_550), .C(n_572), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_468), .B(n_489), .C(n_500), .Y(n_454) );
INVxp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_456), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g659 ( .A(n_456), .B(n_576), .Y(n_659) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g561 ( .A(n_457), .B(n_492), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_457), .B(n_479), .Y(n_678) );
INVx1_ASAP7_75t_L g696 ( .A(n_457), .Y(n_696) );
AND2x2_ASAP7_75t_L g705 ( .A(n_457), .B(n_593), .Y(n_705) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g588 ( .A(n_458), .B(n_479), .Y(n_588) );
AND2x2_ASAP7_75t_L g646 ( .A(n_458), .B(n_593), .Y(n_646) );
INVx1_ASAP7_75t_L g690 ( .A(n_458), .Y(n_690) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g567 ( .A(n_459), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g575 ( .A(n_459), .Y(n_575) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_459), .Y(n_615) );
INVxp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_477), .Y(n_469) );
AND2x2_ASAP7_75t_L g554 ( .A(n_470), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g587 ( .A(n_470), .Y(n_587) );
OR2x2_ASAP7_75t_L g713 ( .A(n_470), .B(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_470), .B(n_479), .Y(n_717) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
INVx1_ASAP7_75t_L g503 ( .A(n_471), .Y(n_503) );
AND2x2_ASAP7_75t_L g576 ( .A(n_471), .B(n_494), .Y(n_576) );
AND2x2_ASAP7_75t_L g616 ( .A(n_471), .B(n_495), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_476), .A2(n_543), .B(n_546), .Y(n_542) );
INVxp67_ASAP7_75t_L g658 ( .A(n_477), .Y(n_658) );
AND2x4_ASAP7_75t_L g683 ( .A(n_477), .B(n_576), .Y(n_683) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_SL g574 ( .A(n_478), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g493 ( .A(n_479), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g562 ( .A(n_479), .B(n_495), .Y(n_562) );
INVx1_ASAP7_75t_L g568 ( .A(n_479), .Y(n_568) );
INVx2_ASAP7_75t_L g594 ( .A(n_479), .Y(n_594) );
AND2x2_ASAP7_75t_L g610 ( .A(n_479), .B(n_611), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_490), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx2_ASAP7_75t_L g565 ( .A(n_492), .Y(n_565) );
AND2x2_ASAP7_75t_L g673 ( .A(n_492), .B(n_494), .Y(n_673) );
AND2x2_ASAP7_75t_L g590 ( .A(n_493), .B(n_575), .Y(n_590) );
AND2x2_ASAP7_75t_L g689 ( .A(n_493), .B(n_690), .Y(n_689) );
NOR2xp67_ASAP7_75t_L g611 ( .A(n_494), .B(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g714 ( .A(n_494), .B(n_575), .Y(n_714) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g504 ( .A(n_495), .Y(n_504) );
AND2x2_ASAP7_75t_L g593 ( .A(n_495), .B(n_594), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_498), .A2(n_526), .B(n_528), .C(n_529), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_498), .A2(n_538), .B(n_539), .Y(n_537) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_504), .Y(n_501) );
AND2x2_ASAP7_75t_L g639 ( .A(n_502), .B(n_574), .Y(n_639) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_503), .B(n_575), .Y(n_624) );
INVx2_ASAP7_75t_L g623 ( .A(n_504), .Y(n_623) );
OAI222xp33_ASAP7_75t_L g627 ( .A1(n_504), .A2(n_567), .B1(n_628), .B2(n_630), .C1(n_631), .C2(n_634), .Y(n_627) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
OR2x2_ASAP7_75t_L g663 ( .A(n_509), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g585 ( .A(n_510), .Y(n_585) );
NOR2x1_ASAP7_75t_L g636 ( .A(n_510), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g642 ( .A(n_510), .B(n_556), .Y(n_642) );
AND2x4_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g603 ( .A(n_511), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_516), .A2(n_606), .B1(n_645), .B2(n_646), .Y(n_644) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_531), .Y(n_516) );
INVx3_ASAP7_75t_L g578 ( .A(n_517), .Y(n_578) );
OR2x2_ASAP7_75t_L g711 ( .A(n_517), .B(n_587), .Y(n_711) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g584 ( .A(n_518), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g600 ( .A(n_518), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g608 ( .A(n_518), .B(n_556), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_518), .B(n_532), .Y(n_664) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g555 ( .A(n_519), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g559 ( .A(n_519), .B(n_532), .Y(n_559) );
AND2x2_ASAP7_75t_L g635 ( .A(n_519), .B(n_582), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_519), .B(n_541), .Y(n_675) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_531), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_552), .Y(n_591) );
AND2x2_ASAP7_75t_L g595 ( .A(n_531), .B(n_585), .Y(n_595) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_541), .Y(n_531) );
INVx3_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
AND2x2_ASAP7_75t_L g581 ( .A(n_532), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g716 ( .A(n_532), .B(n_699), .Y(n_716) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_541), .Y(n_570) );
INVx2_ASAP7_75t_L g582 ( .A(n_541), .Y(n_582) );
AND2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_602), .Y(n_626) );
INVx1_ASAP7_75t_L g669 ( .A(n_541), .Y(n_669) );
OR2x2_ASAP7_75t_L g700 ( .A(n_541), .B(n_602), .Y(n_700) );
AND2x2_ASAP7_75t_L g720 ( .A(n_541), .B(n_556), .Y(n_720) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_553), .B(n_557), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g558 ( .A(n_552), .B(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_552), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g677 ( .A(n_554), .Y(n_677) );
INVx2_ASAP7_75t_SL g571 ( .A(n_555), .Y(n_571) );
AND2x2_ASAP7_75t_L g691 ( .A(n_555), .B(n_585), .Y(n_691) );
INVx2_ASAP7_75t_L g637 ( .A(n_556), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_556), .B(n_669), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_560), .B1(n_563), .B2(n_569), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_559), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g725 ( .A(n_559), .Y(n_725) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g650 ( .A(n_561), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_561), .B(n_593), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_562), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g666 ( .A(n_562), .B(n_615), .Y(n_666) );
INVx2_ASAP7_75t_L g722 ( .A(n_562), .Y(n_722) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g592 ( .A(n_565), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_565), .B(n_610), .Y(n_643) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_567), .B(n_587), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g704 ( .A(n_570), .Y(n_704) );
O2A1O1Ixp33_ASAP7_75t_SL g654 ( .A1(n_571), .A2(n_655), .B(n_657), .C(n_660), .Y(n_654) );
OR2x2_ASAP7_75t_L g681 ( .A(n_571), .B(n_585), .Y(n_681) );
OAI221xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_577), .B1(n_579), .B2(n_586), .C(n_589), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_574), .B(n_623), .Y(n_630) );
AND2x2_ASAP7_75t_L g672 ( .A(n_574), .B(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g708 ( .A(n_574), .Y(n_708) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_575), .Y(n_599) );
INVx1_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
NOR2xp67_ASAP7_75t_L g632 ( .A(n_578), .B(n_633), .Y(n_632) );
INVxp67_ASAP7_75t_L g686 ( .A(n_578), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_578), .B(n_626), .Y(n_702) );
INVx2_ASAP7_75t_L g688 ( .A(n_579), .Y(n_688) );
OR2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g629 ( .A(n_581), .B(n_600), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_581), .A2(n_597), .B(n_639), .C(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g607 ( .A(n_582), .B(n_602), .Y(n_607) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_586), .B(n_685), .Y(n_684) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g655 ( .A(n_587), .B(n_656), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_592), .B2(n_595), .Y(n_589) );
INVx1_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
INVx1_ASAP7_75t_L g656 ( .A(n_593), .Y(n_656) );
INVx1_ASAP7_75t_L g707 ( .A(n_595), .Y(n_707) );
AOI211xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_600), .B(n_604), .C(n_627), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g619 ( .A(n_599), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g670 ( .A(n_600), .Y(n_670) );
AND2x2_ASAP7_75t_L g719 ( .A(n_600), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_609), .B(n_617), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g633 ( .A(n_607), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_607), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g625 ( .A(n_608), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g701 ( .A(n_608), .Y(n_701) );
OAI32xp33_ASAP7_75t_L g712 ( .A1(n_608), .A2(n_660), .A3(n_667), .B1(n_708), .B2(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_613), .Y(n_609) );
INVx1_ASAP7_75t_SL g680 ( .A(n_610), .Y(n_680) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_SL g620 ( .A(n_616), .Y(n_620) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_625), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_619), .A2(n_667), .B1(n_693), .B2(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_623), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g660 ( .A(n_626), .Y(n_660) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B(n_644), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_646), .A2(n_688), .B1(n_689), .B2(n_691), .C(n_692), .Y(n_687) );
NAND5xp2_ASAP7_75t_L g647 ( .A(n_648), .B(n_671), .C(n_687), .D(n_697), .E(n_715), .Y(n_647) );
AOI211xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_651), .B(n_654), .C(n_661), .Y(n_648) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g718 ( .A(n_655), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_665), .B2(n_667), .Y(n_661) );
INVx1_ASAP7_75t_SL g694 ( .A(n_664), .Y(n_694) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI322xp33_ASAP7_75t_L g676 ( .A1(n_667), .A2(n_677), .A3(n_678), .B1(n_679), .B2(n_680), .C1(n_681), .C2(n_682), .Y(n_676) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g679 ( .A(n_669), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_669), .B(n_694), .Y(n_693) );
AOI211xp5_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_674), .B(n_676), .C(n_684), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g706 ( .A1(n_680), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_706) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g723 ( .A(n_690), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_705), .B1(n_706), .B2(n_710), .C(n_712), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_701), .B(n_702), .C(n_703), .Y(n_698) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g724 ( .A(n_700), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B1(n_718), .B2(n_719), .C(n_721), .Y(n_715) );
AOI21xp33_ASAP7_75t_SL g721 ( .A1(n_722), .A2(n_723), .B(n_724), .Y(n_721) );
CKINVDCx16_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
NAND2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
endmodule