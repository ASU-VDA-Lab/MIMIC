module fake_jpeg_13451_n_551 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_551);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_551;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_10),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_57),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_59),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_61),
.Y(n_152)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_18),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_70),
.Y(n_128)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_17),
.Y(n_70)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_74),
.A2(n_39),
.B1(n_36),
.B2(n_34),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_25),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_86),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_41),
.B(n_30),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_25),
.B(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_106),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx5_ASAP7_75t_SL g118 ( 
.A(n_107),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_58),
.A2(n_29),
.B1(n_49),
.B2(n_48),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_112),
.A2(n_116),
.B1(n_129),
.B2(n_49),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_46),
.B1(n_52),
.B2(n_30),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_125),
.B(n_139),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_47),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_127),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_59),
.A2(n_46),
.B1(n_28),
.B2(n_39),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_94),
.B(n_28),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_167),
.B1(n_48),
.B2(n_24),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g143 ( 
.A1(n_57),
.A2(n_34),
.B(n_36),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_172),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_82),
.B(n_53),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_165),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_99),
.B(n_44),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_20),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_60),
.A2(n_24),
.B1(n_29),
.B2(n_49),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_61),
.B(n_44),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_171),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_63),
.B(n_51),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_104),
.B(n_51),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g272 ( 
.A1(n_173),
.A2(n_218),
.B1(n_152),
.B2(n_145),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_121),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_174),
.Y(n_253)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_112),
.A2(n_87),
.B1(n_88),
.B2(n_96),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_177),
.A2(n_178),
.B1(n_208),
.B2(n_219),
.Y(n_262)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_107),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_180),
.B(n_217),
.Y(n_285)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_181),
.Y(n_251)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_182),
.Y(n_256)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_42),
.B1(n_43),
.B2(n_92),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_185),
.A2(n_207),
.B1(n_226),
.B2(n_234),
.Y(n_242)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_216),
.Y(n_243)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_119),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_191),
.A2(n_182),
.B1(n_198),
.B2(n_200),
.Y(n_238)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_194),
.Y(n_277)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_196),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_197),
.Y(n_257)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_198),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_123),
.B(n_47),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_199),
.Y(n_288)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_200),
.Y(n_281)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_115),
.Y(n_201)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_202),
.Y(n_260)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_204),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_48),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_225),
.Y(n_250)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_159),
.Y(n_206)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_126),
.A2(n_91),
.B1(n_24),
.B2(n_29),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_128),
.A2(n_106),
.B1(n_105),
.B2(n_50),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_212),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_149),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_20),
.B1(n_50),
.B2(n_47),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_128),
.A2(n_50),
.B1(n_2),
.B2(n_4),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_220),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_164),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_222),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_120),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_124),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_223),
.B(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_122),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_158),
.B(n_1),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_156),
.A2(n_50),
.B1(n_5),
.B2(n_6),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_50),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_232),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_4),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_233),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_120),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_230),
.B(n_5),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_110),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_231),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_286)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_151),
.B(n_16),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_110),
.B(n_4),
.Y(n_233)
);

INVx3_ASAP7_75t_SL g234 ( 
.A(n_146),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_238),
.A2(n_240),
.B1(n_180),
.B2(n_220),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_191),
.A2(n_141),
.B1(n_161),
.B2(n_122),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_255),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_177),
.A2(n_146),
.B1(n_161),
.B2(n_141),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_248),
.A2(n_286),
.B1(n_189),
.B2(n_211),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_197),
.A2(n_111),
.B1(n_114),
.B2(n_169),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_254),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_203),
.A2(n_155),
.A3(n_152),
.B1(n_145),
.B2(n_142),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_180),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_199),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_267),
.B(n_215),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_193),
.B(n_166),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_270),
.B(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_203),
.B(n_166),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_233),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_232),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_193),
.B(n_6),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_234),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_279),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_176),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_228),
.B(n_184),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_184),
.B(n_9),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_232),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_289),
.B(n_302),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_290),
.B(n_314),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_291),
.B(n_304),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_184),
.B1(n_228),
.B2(n_205),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_294),
.A2(n_298),
.B(n_258),
.Y(n_376)
);

OA22x2_ASAP7_75t_L g361 ( 
.A1(n_295),
.A2(n_322),
.B1(n_257),
.B2(n_278),
.Y(n_361)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_299),
.B(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_301),
.A2(n_307),
.B1(n_321),
.B2(n_257),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_243),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_240),
.A2(n_232),
.B1(n_199),
.B2(n_192),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_303),
.A2(n_312),
.B1(n_315),
.B2(n_319),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_250),
.B(n_210),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_229),
.B(n_225),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_217),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_306),
.B(n_326),
.C(n_337),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_277),
.A2(n_183),
.B1(n_194),
.B2(n_222),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_250),
.B(n_212),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_308),
.B(n_316),
.Y(n_352)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_311),
.A2(n_313),
.B1(n_335),
.B2(n_284),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_271),
.A2(n_209),
.B1(n_188),
.B2(n_190),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_262),
.A2(n_196),
.B1(n_179),
.B2(n_186),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_202),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_262),
.A2(n_206),
.B1(n_214),
.B2(n_13),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_266),
.B(n_11),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_241),
.Y(n_318)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_255),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_237),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_320),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_242),
.A2(n_16),
.B1(n_13),
.B2(n_14),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_272),
.A2(n_14),
.B1(n_16),
.B2(n_288),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_246),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_237),
.Y(n_345)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_236),
.Y(n_324)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_324),
.Y(n_368)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_236),
.Y(n_325)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_261),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_288),
.A2(n_272),
.B1(n_285),
.B2(n_261),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_327),
.A2(n_268),
.B1(n_265),
.B2(n_252),
.Y(n_365)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_269),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_328),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_251),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_329),
.B(n_331),
.Y(n_341)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_330),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_263),
.B(n_239),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_273),
.B(n_287),
.Y(n_332)
);

OAI21xp33_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_265),
.B(n_268),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_280),
.B(n_249),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_333),
.A2(n_327),
.B(n_301),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_285),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_334),
.B(n_302),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_272),
.A2(n_286),
.B1(n_252),
.B2(n_259),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_283),
.B(n_273),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_303),
.B1(n_335),
.B2(n_313),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_342),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_284),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_297),
.B(n_260),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_344),
.B(n_347),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_345),
.B(n_350),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_260),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_314),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_353),
.A2(n_364),
.B(n_377),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_324),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_360),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_278),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_356),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_306),
.B(n_276),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_325),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_361),
.B(n_296),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_276),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_362),
.B(n_370),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_365),
.A2(n_328),
.B1(n_317),
.B2(n_300),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_366),
.B(n_376),
.C(n_339),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_337),
.B(n_244),
.Y(n_370)
);

OAI32xp33_ASAP7_75t_L g373 ( 
.A1(n_293),
.A2(n_244),
.A3(n_258),
.B1(n_294),
.B2(n_301),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_379),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_310),
.A2(n_333),
.B(n_334),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_378),
.B(n_341),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_312),
.B(n_330),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_364),
.A2(n_315),
.B1(n_319),
.B2(n_295),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_381),
.A2(n_387),
.B1(n_389),
.B2(n_405),
.Y(n_419)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_377),
.A2(n_336),
.B(n_310),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_386),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_363),
.A2(n_353),
.B(n_374),
.Y(n_386)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_390),
.Y(n_437)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_336),
.B(n_292),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_393),
.Y(n_438)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_392),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g393 ( 
.A(n_374),
.B(n_305),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_371),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_408),
.Y(n_439)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_395),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_409),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_320),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_347),
.Y(n_420)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_401),
.Y(n_423)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_402),
.Y(n_424)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_346),
.Y(n_403)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_403),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_338),
.A2(n_289),
.B1(n_309),
.B2(n_318),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_357),
.A2(n_299),
.B1(n_365),
.B2(n_355),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_407),
.A2(n_414),
.B1(n_344),
.B2(n_342),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_345),
.Y(n_408)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_343),
.A2(n_373),
.B1(n_370),
.B2(n_361),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_413),
.Y(n_418)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_359),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_343),
.B1(n_361),
.B2(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_415),
.B(n_367),
.Y(n_425)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_420),
.Y(n_462)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_359),
.Y(n_426)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_390),
.Y(n_427)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_367),
.Y(n_428)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_428),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_349),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_433),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_356),
.Y(n_430)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_430),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_431),
.A2(n_412),
.B1(n_411),
.B2(n_380),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_397),
.B(n_340),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_432),
.B(n_429),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_383),
.B(n_362),
.Y(n_433)
);

BUFx8_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_436),
.B(n_396),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_397),
.B(n_376),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_441),
.B(n_442),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_348),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_405),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_398),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_358),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_446),
.C(n_433),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_414),
.B(n_375),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g493 ( 
.A(n_447),
.B(n_459),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_386),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_448),
.B(n_451),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_452),
.B(n_442),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_418),
.A2(n_400),
.B1(n_411),
.B2(n_389),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_453),
.A2(n_457),
.B1(n_466),
.B2(n_461),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_435),
.A2(n_384),
.B(n_400),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_456),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_351),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_389),
.B1(n_385),
.B2(n_380),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_439),
.B(n_410),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_472),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_432),
.B(n_407),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_391),
.C(n_394),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_465),
.C(n_470),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_461),
.B(n_419),
.Y(n_476)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_463),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_SL g465 ( 
.A(n_438),
.B(n_352),
.C(n_403),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_382),
.B1(n_392),
.B2(n_395),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_402),
.C(n_401),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_388),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_425),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_454),
.Y(n_475)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_475),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_476),
.Y(n_505)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_479),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_480),
.B(n_488),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_451),
.A2(n_419),
.B1(n_440),
.B2(n_416),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_482),
.A2(n_484),
.B1(n_487),
.B2(n_492),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_428),
.Y(n_483)
);

AOI21x1_ASAP7_75t_SL g501 ( 
.A1(n_483),
.A2(n_494),
.B(n_489),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_453),
.A2(n_416),
.B1(n_446),
.B2(n_436),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_466),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_486),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_467),
.B(n_452),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_449),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_420),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_468),
.B(n_445),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_490),
.B(n_447),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_459),
.C(n_462),
.Y(n_507)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_469),
.B(n_417),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_498),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_491),
.B(n_468),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_470),
.C(n_460),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_507),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_448),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_493),
.Y(n_525)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_478),
.A2(n_465),
.B(n_455),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_503),
.A2(n_477),
.B(n_494),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_482),
.B(n_457),
.Y(n_504)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_504),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_462),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_484),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_474),
.B(n_436),
.C(n_422),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_511),
.C(n_499),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_474),
.B(n_421),
.C(n_423),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_511),
.B(n_481),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_513),
.B(n_522),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_525),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_495),
.B(n_483),
.Y(n_518)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_518),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_519),
.B(n_523),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_520),
.A2(n_501),
.B(n_504),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_477),
.C(n_480),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_521),
.B(n_496),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_502),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_505),
.B(n_427),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_473),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_524),
.A2(n_476),
.B(n_434),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_528),
.A2(n_520),
.B(n_516),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_531),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_424),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_524),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g537 ( 
.A1(n_532),
.A2(n_529),
.B1(n_531),
.B2(n_517),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_514),
.A2(n_496),
.B1(n_493),
.B2(n_509),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_533),
.B(n_535),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_SL g536 ( 
.A(n_527),
.B(n_515),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_536),
.A2(n_537),
.B(n_538),
.Y(n_542)
);

A2O1A1Ixp33_ASAP7_75t_SL g539 ( 
.A1(n_528),
.A2(n_519),
.B(n_521),
.C(n_525),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_526),
.C(n_512),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_540),
.B(n_530),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_543),
.B(n_544),
.Y(n_545)
);

O2A1O1Ixp33_ASAP7_75t_SL g546 ( 
.A1(n_542),
.A2(n_541),
.B(n_533),
.C(n_534),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_546),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g548 ( 
.A1(n_547),
.A2(n_545),
.B(n_526),
.Y(n_548)
);

MAJx2_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_512),
.C(n_498),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_549),
.B(n_500),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_497),
.C(n_437),
.Y(n_551)
);


endmodule