module fake_jpeg_26647_n_57 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_57);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_57;

wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_37),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_30),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_41),
.A2(n_32),
.B(n_34),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_28),
.CI(n_25),
.CON(n_42),
.SN(n_42)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_28),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_47),
.B(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_48),
.A2(n_38),
.B1(n_45),
.B2(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

AO21x1_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_51),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_41),
.Y(n_54)
);

AOI322xp5_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_7),
.A3(n_8),
.B1(n_10),
.B2(n_12),
.C1(n_13),
.C2(n_14),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_19),
.C1(n_21),
.C2(n_22),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_24),
.Y(n_57)
);


endmodule