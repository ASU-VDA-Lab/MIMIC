module fake_jpeg_30976_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_28),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_62),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_0),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_67),
.Y(n_81)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_48),
.B(n_1),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_2),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_53),
.B1(n_56),
.B2(n_42),
.Y(n_70)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_79),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_56),
.B1(n_42),
.B2(n_48),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_59),
.B1(n_55),
.B2(n_50),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_41),
.B1(n_43),
.B2(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_76),
.B1(n_71),
.B2(n_70),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_43),
.C(n_50),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_46),
.B1(n_58),
.B2(n_57),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_67),
.A2(n_49),
.B(n_51),
.C(n_47),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_93),
.B1(n_95),
.B2(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_96),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_94),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_23),
.B1(n_38),
.B2(n_37),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_2),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_72),
.B1(n_82),
.B2(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_3),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_11),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_4),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_6),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_27),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_89),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_95),
.B(n_83),
.C(n_92),
.D(n_84),
.Y(n_113)
);

NAND5xp2_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_120),
.C(n_40),
.D(n_20),
.E(n_22),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_114),
.B(n_117),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_30),
.C(n_36),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_119),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_12),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_31),
.C(n_34),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_26),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_122),
.A2(n_128),
.B1(n_105),
.B2(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_115),
.C(n_126),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_109),
.Y(n_136)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_132),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_122),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_140),
.B1(n_130),
.B2(n_138),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_107),
.B1(n_112),
.B2(n_113),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_140),
.A3(n_129),
.B1(n_102),
.B2(n_120),
.C1(n_108),
.C2(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_133),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_129),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_104),
.B1(n_134),
.B2(n_137),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_123),
.Y(n_146)
);


endmodule