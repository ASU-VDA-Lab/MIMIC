module fake_jpeg_10938_n_30 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_15;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

NAND3xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_1),
.C(n_2),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_13),
.B(n_9),
.C(n_8),
.D(n_7),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_10),
.B(n_13),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_19),
.C(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_14),
.B1(n_10),
.B2(n_11),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_24),
.B(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_28),
.B1(n_26),
.B2(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_3),
.Y(n_30)
);


endmodule