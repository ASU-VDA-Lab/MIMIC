module real_jpeg_1952_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_69),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_30),
.B1(n_37),
.B2(n_69),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_2),
.B(n_57),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_2),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_2),
.A2(n_57),
.B(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_2),
.B(n_78),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_2),
.A2(n_65),
.B(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_2),
.B(n_30),
.C(n_46),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_205),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_2),
.B(n_32),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_2),
.B(n_51),
.Y(n_260)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_4),
.A2(n_57),
.B1(n_58),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_4),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_179),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_179),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_4),
.A2(n_30),
.B1(n_37),
.B2(n_179),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_5),
.A2(n_30),
.B1(n_37),
.B2(n_75),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_7),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_30),
.B1(n_37),
.B2(n_50),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_7),
.A2(n_50),
.B1(n_57),
.B2(n_58),
.Y(n_306)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_67),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_9),
.A2(n_30),
.B1(n_37),
.B2(n_67),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_10),
.A2(n_36),
.B1(n_57),
.B2(n_58),
.Y(n_314)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_13),
.A2(n_64),
.B1(n_65),
.B2(n_125),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_125),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_13),
.A2(n_30),
.B1(n_37),
.B2(n_125),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_14),
.A2(n_57),
.B1(n_58),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_14),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_159),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_14),
.A2(n_30),
.B1(n_37),
.B2(n_159),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_16),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_16),
.A2(n_41),
.B1(n_64),
.B2(n_65),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_16),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_16),
.A2(n_30),
.B1(n_37),
.B2(n_41),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_311),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_298),
.B(n_310),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_139),
.B(n_295),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_126),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_99),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_23),
.B(n_99),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_70),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_24),
.B(n_85),
.C(n_97),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_52),
.B(n_53),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_25),
.A2(n_26),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_27),
.A2(n_52),
.B1(n_53),
.B2(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_27),
.A2(n_38),
.B1(n_39),
.B2(n_52),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B(n_34),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_28),
.A2(n_31),
.B1(n_113),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_28),
.A2(n_31),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_28),
.A2(n_31),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_29),
.A2(n_32),
.B1(n_35),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_29),
.A2(n_32),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_29),
.A2(n_32),
.B1(n_172),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_29),
.A2(n_32),
.B1(n_209),
.B2(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_29),
.A2(n_32),
.B1(n_205),
.B2(n_258),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_29),
.A2(n_32),
.B1(n_258),
.B2(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_37),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_30),
.B(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_40),
.A2(n_44),
.B1(n_51),
.B2(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_42),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

AO22x2_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_43),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_65),
.A3(n_79),
.B1(n_204),
.B2(n_206),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_42),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_43),
.B(n_80),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_44),
.A2(n_49),
.B1(n_51),
.B2(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_51),
.B(n_84),
.Y(n_91)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_44),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_44),
.A2(n_51),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_44),
.A2(n_51),
.B1(n_201),
.B2(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_44),
.A2(n_51),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_44),
.A2(n_51),
.B1(n_228),
.B2(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_48),
.A2(n_117),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_48),
.A2(n_152),
.B1(n_200),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_63),
.B1(n_68),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_54),
.A2(n_63),
.B1(n_66),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_54),
.A2(n_63),
.B1(n_88),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_54),
.A2(n_63),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_54),
.A2(n_63),
.B1(n_178),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_55),
.A2(n_124),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_55),
.A2(n_160),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_55),
.A2(n_160),
.B1(n_306),
.B2(n_314),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_63),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI32xp33_ASAP7_75t_L g168 ( 
.A1(n_58),
.A2(n_62),
.A3(n_65),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g170 ( 
.A(n_60),
.B(n_64),
.Y(n_170)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_65),
.B1(n_79),
.B2(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_64),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_85),
.B1(n_97),
.B2(n_98),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_71),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_72),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_83),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_76),
.B1(n_78),
.B2(n_82),
.Y(n_72)
);

INVxp33_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_74),
.A2(n_77),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_78),
.B1(n_82),
.B2(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_76),
.A2(n_78),
.B1(n_120),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_76),
.A2(n_78),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_77),
.A2(n_95),
.B1(n_121),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_77),
.A2(n_121),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_77),
.A2(n_121),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_77),
.A2(n_121),
.B1(n_175),
.B2(n_191),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_77),
.A2(n_121),
.B1(n_190),
.B2(n_237),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_79),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_87),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_87),
.B(n_91),
.C(n_93),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_87),
.B(n_130),
.C(n_137),
.Y(n_299)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_96),
.Y(n_90)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_96),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_91),
.B(n_133),
.C(n_135),
.Y(n_309)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_105),
.C(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_142)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_118),
.C(n_122),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_108),
.A2(n_109),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_122),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_126),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_138),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_127),
.B(n_138),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_134),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_136),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_161),
.B(n_294),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_141),
.B(n_143),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_148),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.C(n_157),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_150),
.B(n_153),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_157),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_184),
.B(n_293),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_182),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_163),
.B(n_182),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_181),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_164),
.B(n_181),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_166),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.C(n_177),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_167),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_171),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_174),
.B(n_177),
.Y(n_284)
);

AOI31xp33_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_278),
.A3(n_287),
.B(n_290),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_223),
.B(n_277),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_211),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_187),
.B(n_211),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_198),
.C(n_202),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_188),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_193),
.C(n_197),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_202),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_207),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_207),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_204),
.Y(n_238)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_211),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_211),
.B(n_288),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.CI(n_214),
.CON(n_211),
.SN(n_211)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_215),
.B(n_218),
.C(n_222),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_272),
.B(n_276),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_241),
.B(n_271),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_233),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_233),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_231),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_230),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_251),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_236),
.C(n_239),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_252),
.B(n_270),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_250),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_248),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_264),
.B(n_269),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_259),
.B(n_263),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_261),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_268),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_275),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_279),
.A2(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_282),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_309),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_304),
.B1(n_307),
.B2(n_308),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_307),
.C(n_309),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);


endmodule