module fake_jpeg_3257_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_33),
.Y(n_54)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_64),
.B1(n_66),
.B2(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_48),
.B1(n_41),
.B2(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_42),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_56),
.A2(n_47),
.B1(n_53),
.B2(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_34),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_78),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_69),
.B(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_77),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_79),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_38),
.B1(n_51),
.B2(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_0),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_76),
.A2(n_61),
.B1(n_60),
.B2(n_59),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_75),
.A2(n_60),
.B1(n_59),
.B2(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_88),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_84),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_1),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_86),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_14),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_92),
.B(n_22),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_18),
.C(n_28),
.Y(n_92)
);

AOI22x1_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_16),
.B1(n_27),
.B2(n_26),
.Y(n_94)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_83),
.B(n_91),
.C(n_89),
.D(n_93),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_31),
.C(n_24),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_5),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_107),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_23),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_10),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_7),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_109),
.B(n_11),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_111),
.B(n_19),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_118),
.C(n_120),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_101),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_119),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_98),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_15),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_13),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_12),
.B(n_13),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_96),
.B(n_95),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_97),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_123),
.B(n_121),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_117),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_128),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_126),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_120),
.Y(n_133)
);

INVxp33_ASAP7_75t_SL g135 ( 
.A(n_133),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_136),
.B(n_124),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_132),
.C(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_114),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_118),
.Y(n_140)
);


endmodule