module real_jpeg_11888_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_221;
wire n_215;
wire n_292;
wire n_288;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_290;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_259;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_244;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_29),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_1),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_1),
.A2(n_37),
.B1(n_60),
.B2(n_63),
.Y(n_287)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_29),
.B1(n_36),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_3),
.A2(n_53),
.B1(n_60),
.B2(n_63),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_5),
.A2(n_60),
.B1(n_63),
.B2(n_68),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_5),
.A2(n_29),
.B1(n_36),
.B2(n_68),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_29),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_7),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_8),
.A2(n_65),
.B1(n_66),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_8),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_8),
.A2(n_60),
.B1(n_63),
.B2(n_101),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_101),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_8),
.A2(n_29),
.B1(n_36),
.B2(n_101),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g131 ( 
.A1(n_9),
.A2(n_65),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_9),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_9),
.B(n_63),
.Y(n_189)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_134),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_9),
.A2(n_44),
.B(n_49),
.C(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_109),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_9),
.B(n_33),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_9),
.B(n_54),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_9),
.A2(n_63),
.B(n_189),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_10),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_60),
.B1(n_63),
.B2(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_136),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_29),
.B1(n_36),
.B2(n_136),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_14),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_14),
.A2(n_60),
.B1(n_63),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_70),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_14),
.A2(n_29),
.B1(n_36),
.B2(n_70),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_60),
.B1(n_63),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_15),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_78),
.Y(n_160)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_17),
.A2(n_46),
.B1(n_60),
.B2(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_17),
.A2(n_29),
.B1(n_36),
.B2(n_46),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_17),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_280)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_271),
.B1(n_293),
.B2(n_294),
.Y(n_19)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_20),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_124),
.B(n_270),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_102),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_22),
.B(n_102),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_80),
.C(n_86),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_23),
.B(n_80),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_55),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_24),
.B(n_57),
.C(n_71),
.Y(n_123)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_28),
.A2(n_33),
.B(n_38),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_28),
.A2(n_33),
.B1(n_92),
.B2(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_33),
.B1(n_148),
.B2(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_28),
.A2(n_33),
.B1(n_160),
.B2(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_28),
.A2(n_33),
.B1(n_192),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_28),
.A2(n_33),
.B1(n_134),
.B2(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_28),
.A2(n_33),
.B1(n_218),
.B2(n_225),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_29),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_32),
.A2(n_35),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_32),
.A2(n_90),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_36),
.A2(n_50),
.B(n_134),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_43),
.A2(n_51),
.B1(n_94),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_45),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_45),
.B1(n_74),
.B2(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_44),
.B(n_75),
.Y(n_190)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_45),
.A2(n_63),
.A3(n_74),
.B1(n_188),
.B2(n_190),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_84),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_47),
.A2(n_54),
.B1(n_84),
.B2(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_47),
.A2(n_54),
.B1(n_95),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_47),
.A2(n_54),
.B1(n_142),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_47),
.A2(n_54),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_47),
.A2(n_54),
.B1(n_204),
.B2(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_47),
.A2(n_54),
.B(n_111),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_51),
.A2(n_96),
.B1(n_183),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_71),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_59),
.B1(n_67),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_59),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_58),
.A2(n_59),
.B1(n_131),
.B2(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_58),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_58),
.A2(n_59),
.B1(n_120),
.B2(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_63),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_60),
.A2(n_62),
.A3(n_65),
.B1(n_133),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_63),
.Y(n_151)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_66),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_76),
.B1(n_77),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_72),
.A2(n_76),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_72),
.A2(n_76),
.B1(n_155),
.B2(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_85),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_81),
.A2(n_82),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_82),
.A2(n_119),
.B(n_121),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_86),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_97),
.C(n_99),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_87),
.A2(n_88),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_89),
.B(n_93),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_97),
.B(n_99),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_123),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B(n_112),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_109),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_107),
.A2(n_109),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_286),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_112),
.A2(n_277),
.B1(n_289),
.B2(n_290),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_112),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_113),
.B(n_122),
.C(n_123),
.Y(n_291)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_265),
.B(n_269),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_175),
.B(n_253),
.C(n_264),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_161),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_127),
.B(n_161),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_145),
.C(n_152),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_128),
.A2(n_129),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_138),
.C(n_144),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_143),
.B2(n_144),
.Y(n_137)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_139),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_145),
.B(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_159),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_163),
.B(n_164),
.C(n_165),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_174),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_167),
.B(n_170),
.C(n_174),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_252),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_196),
.B(n_251),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_193),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_178),
.B(n_193),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.C(n_184),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_179),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_181),
.A2(n_184),
.B1(n_185),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_181),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_186),
.A2(n_187),
.B1(n_191),
.B2(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_245),
.B(n_250),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_234),
.B(n_244),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_214),
.B(n_233),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_200),
.B(n_207),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_210),
.C(n_212),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_211),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_222),
.B(n_232),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_216),
.B(n_220),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_228),
.B(n_231),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_229),
.B(n_230),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_235),
.B(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_240),
.C(n_242),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_255),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_263),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_262),
.C(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_258),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_267),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_292),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_291),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_291),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_283),
.Y(n_288)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);


endmodule