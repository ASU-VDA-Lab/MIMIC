module fake_netlist_5_1656_n_2048 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2048);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2048;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1587;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1951;
wire n_1825;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_38),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_146),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_204),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_131),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_107),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_34),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_41),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_116),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_32),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_76),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_30),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_41),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_47),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_70),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_48),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_38),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_79),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_9),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_186),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_189),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_90),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_89),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_64),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_80),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_39),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_106),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_123),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_137),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_6),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_150),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_81),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_130),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_113),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_64),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_139),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_74),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_82),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_57),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_114),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_166),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_175),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_78),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_4),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_105),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_120),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_153),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_46),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_183),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_62),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_133),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_73),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_12),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_84),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_136),
.Y(n_283)
);

BUFx10_ASAP7_75t_L g284 ( 
.A(n_181),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_62),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_10),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_46),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_10),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_68),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_140),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_59),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_54),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_182),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_94),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_199),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_110),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_52),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_36),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_9),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_15),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_71),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_169),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_125),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_58),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_190),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_11),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_164),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_197),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_141),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_205),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_91),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_8),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_152),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_57),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_58),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_201),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_132),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_98),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_118),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_142),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_149),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_19),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_17),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_200),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_172),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_39),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_15),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_75),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_127),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_11),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_66),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_65),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_77),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_63),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_22),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_99),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_21),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_117),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_55),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_147),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_97),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_88),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_52),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_69),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_206),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_185),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_63),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_17),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_103),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_54),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_56),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_1),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_27),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_0),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_26),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_188),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_72),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_93),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_3),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_40),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_155),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_16),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_178),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_104),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_34),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_66),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

INVx4_ASAP7_75t_R g369 ( 
.A(n_28),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_23),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_44),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_12),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_31),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_161),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_129),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_85),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_27),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_194),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_86),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_16),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_87),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_18),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_5),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_35),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_111),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_13),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_151),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_202),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_24),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_121),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_60),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_203),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_3),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_7),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_50),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_192),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_92),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_36),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_47),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_48),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_135),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_32),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_173),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_25),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_13),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_19),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_51),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_7),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_33),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_144),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_0),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_253),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_258),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_262),
.Y(n_414)
);

INVxp33_ASAP7_75t_SL g415 ( 
.A(n_289),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_293),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g417 ( 
.A(n_292),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_215),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_215),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_215),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_211),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_215),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_215),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_215),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_215),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_215),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_218),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_267),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_268),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_327),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_327),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_327),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_327),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_229),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_274),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_327),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_244),
.Y(n_437)
);

BUFx6f_ASAP7_75t_SL g438 ( 
.A(n_284),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_250),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_327),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_400),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_309),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_327),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_256),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_327),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_275),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_277),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_207),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_292),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_305),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_305),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_285),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_406),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_286),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_244),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_302),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_381),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_406),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_406),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_220),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g463 ( 
.A(n_207),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_223),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_224),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_290),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_225),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_223),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_233),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_390),
.Y(n_470)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_216),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_270),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_401),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_230),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_231),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_298),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_245),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_280),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_301),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_330),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_233),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_254),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_287),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_288),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_299),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_255),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_313),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_257),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_216),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_331),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_340),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_259),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_263),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_346),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_315),
.Y(n_495)
);

INVxp33_ASAP7_75t_SL g496 ( 
.A(n_246),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_323),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_354),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_324),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_346),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_354),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_356),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_328),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_356),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_269),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_264),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_265),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_349),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_216),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_351),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_246),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_307),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_271),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_272),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_375),
.Y(n_516)
);

CKINVDCx11_ASAP7_75t_R g517 ( 
.A(n_489),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_446),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_482),
.Y(n_520)
);

BUFx8_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_505),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_454),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_459),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_516),
.B(n_375),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_410),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_457),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_437),
.B(n_410),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_461),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_418),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_437),
.B(n_318),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_456),
.B(n_318),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_456),
.B(n_284),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_431),
.B(n_318),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_500),
.B(n_242),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_513),
.A2(n_380),
.B1(n_333),
.B2(n_394),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_421),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_468),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_468),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_472),
.B(n_284),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_505),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_471),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_444),
.B(n_242),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_419),
.Y(n_547)
);

NOR2x1_ASAP7_75t_L g548 ( 
.A(n_486),
.B(n_248),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_412),
.B(n_311),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_431),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_432),
.B(n_248),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_450),
.B(n_311),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_433),
.B(n_281),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_415),
.A2(n_273),
.B1(n_408),
.B2(n_407),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_480),
.A2(n_316),
.B1(n_408),
.B2(n_407),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_433),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_423),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_412),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_463),
.B(n_320),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_436),
.B(n_281),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_451),
.B(n_303),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_436),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_414),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_505),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_440),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_440),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_505),
.B(n_269),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_443),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_452),
.B(n_311),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_417),
.B(n_303),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_445),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_488),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_424),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_425),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_413),
.A2(n_348),
.B1(n_405),
.B2(n_249),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_445),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_492),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_493),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_426),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_496),
.B(n_321),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_430),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_469),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_464),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_507),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_506),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_464),
.B(n_337),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_414),
.Y(n_591)
);

OA21x2_ASAP7_75t_L g592 ( 
.A1(n_498),
.A2(n_337),
.B(n_214),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_417),
.B(n_212),
.Y(n_593)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_462),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_506),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_509),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_509),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_498),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_562),
.B(n_428),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_519),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_519),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_539),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_584),
.B(n_428),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_539),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_535),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_577),
.B(n_429),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_577),
.B(n_429),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_578),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_577),
.B(n_435),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_527),
.B(n_435),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_527),
.B(n_447),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_539),
.Y(n_612)
);

OR2x6_ASAP7_75t_L g613 ( 
.A(n_548),
.B(n_217),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_551),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_529),
.B(n_501),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_544),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_535),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_553),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_532),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_553),
.B(n_447),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_545),
.B(n_448),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_545),
.B(n_448),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_538),
.A2(n_370),
.B1(n_386),
.B2(n_237),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_559),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_539),
.Y(n_627)
);

NAND3xp33_ASAP7_75t_L g628 ( 
.A(n_546),
.B(n_467),
.C(n_465),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_529),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_565),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_565),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_568),
.B(n_453),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_554),
.B(n_501),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_568),
.B(n_453),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_548),
.B(n_455),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_532),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_547),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_569),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_569),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_554),
.B(n_502),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_571),
.B(n_455),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_573),
.B(n_466),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_573),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_547),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_575),
.Y(n_646)
);

AOI22x1_ASAP7_75t_L g647 ( 
.A1(n_536),
.A2(n_481),
.B1(n_512),
.B2(n_416),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_549),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_575),
.Y(n_649)
);

NAND2xp33_ASAP7_75t_L g650 ( 
.A(n_526),
.B(n_528),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_580),
.B(n_219),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_539),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_549),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_556),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_539),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_556),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_580),
.B(n_466),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_560),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_521),
.B(n_476),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_560),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_521),
.B(n_476),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_579),
.A2(n_441),
.B1(n_391),
.B2(n_300),
.Y(n_662)
);

BUFx10_ASAP7_75t_L g663 ( 
.A(n_566),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_583),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_540),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_583),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_552),
.A2(n_360),
.B1(n_363),
.B2(n_355),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_533),
.B(n_534),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_550),
.B(n_508),
.Y(n_669)
);

AND2x6_ASAP7_75t_L g670 ( 
.A(n_536),
.B(n_269),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_572),
.B(n_589),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_593),
.B(n_510),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_567),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_521),
.B(n_479),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_518),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_523),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_518),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_587),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_587),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_538),
.A2(n_300),
.B1(n_344),
.B2(n_249),
.Y(n_681)
);

XOR2xp5_ASAP7_75t_L g682 ( 
.A(n_558),
.B(n_427),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_587),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_585),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_520),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_544),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_585),
.B(n_479),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_585),
.B(n_487),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_585),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_574),
.B(n_487),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_567),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_524),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_587),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_586),
.B(n_514),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_524),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_536),
.B(n_221),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_525),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_525),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_536),
.B(n_222),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_530),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_567),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_530),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_572),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_567),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_531),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_531),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_521),
.B(n_495),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_578),
.B(n_495),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_598),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_578),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_589),
.B(n_502),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_578),
.B(n_552),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_578),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_543),
.B(n_515),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_567),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_598),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_598),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_578),
.B(n_497),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_595),
.B(n_504),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_522),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_561),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_555),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_522),
.Y(n_725)
);

BUFx4f_ASAP7_75t_L g726 ( 
.A(n_592),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_557),
.A2(n_579),
.B1(n_558),
.B2(n_348),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_544),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_555),
.B(n_497),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_594),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_561),
.B(n_499),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_555),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_SL g734 ( 
.A(n_591),
.B(n_499),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_522),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_595),
.B(n_504),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_563),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_563),
.B(n_227),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_591),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_563),
.Y(n_740)
);

AND3x2_ASAP7_75t_L g741 ( 
.A(n_590),
.B(n_235),
.C(n_234),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_L g742 ( 
.A(n_563),
.B(n_475),
.C(n_474),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_544),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_541),
.Y(n_744)
);

BUFx4f_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_590),
.A2(n_368),
.B1(n_384),
.B2(n_377),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_537),
.B(n_503),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_592),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_541),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_542),
.Y(n_751)
);

INVxp67_ASAP7_75t_L g752 ( 
.A(n_677),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_726),
.B(n_269),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_665),
.B(n_503),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_629),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_665),
.B(n_590),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_629),
.B(n_615),
.Y(n_757)
);

BUFx5_ASAP7_75t_L g758 ( 
.A(n_748),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_614),
.B(n_590),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_614),
.B(n_564),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_709),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_726),
.B(n_269),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_615),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_726),
.B(n_283),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_SL g765 ( 
.A(n_669),
.B(n_716),
.Y(n_765)
);

AND2x6_ASAP7_75t_SL g766 ( 
.A(n_694),
.B(n_398),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_745),
.B(n_283),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_610),
.B(n_594),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_745),
.B(n_283),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_748),
.A2(n_404),
.B1(n_409),
.B2(n_283),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_740),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_618),
.B(n_236),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_618),
.B(n_240),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_745),
.B(n_283),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_619),
.B(n_624),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_611),
.B(n_594),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_714),
.A2(n_542),
.B(n_597),
.Y(n_777)
);

OR2x2_ASAP7_75t_SL g778 ( 
.A(n_672),
.B(n_517),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_633),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_740),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_619),
.B(n_241),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_605),
.B(n_596),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_624),
.B(n_243),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_740),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_633),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_626),
.B(n_247),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_703),
.A2(n_434),
.B1(n_439),
.B2(n_473),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_709),
.Y(n_788)
);

INVxp67_ASAP7_75t_SL g789 ( 
.A(n_749),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_672),
.B(n_576),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_621),
.A2(n_597),
.B(n_596),
.C(n_485),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_626),
.B(n_630),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_671),
.B(n_581),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_L g794 ( 
.A(n_687),
.B(n_276),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_630),
.B(n_251),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_690),
.B(n_739),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_605),
.B(n_310),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_631),
.B(n_252),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_608),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_631),
.B(n_260),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_638),
.B(n_261),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_690),
.B(n_594),
.Y(n_803)
);

AND2x4_ASAP7_75t_L g804 ( 
.A(n_617),
.B(n_477),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_617),
.B(n_310),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_SL g806 ( 
.A(n_599),
.B(n_438),
.Y(n_806)
);

INVx8_ASAP7_75t_L g807 ( 
.A(n_613),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_711),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_711),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_703),
.B(n_310),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_718),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_719),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_582),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_739),
.B(n_588),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_688),
.B(n_310),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_713),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_638),
.B(n_266),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_639),
.B(n_278),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_713),
.A2(n_442),
.B1(n_458),
.B2(n_470),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_719),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_639),
.B(n_282),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_724),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_724),
.B(n_310),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_728),
.A2(n_295),
.B(n_379),
.C(n_378),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_632),
.B(n_208),
.Y(n_825)
);

INVx8_ASAP7_75t_L g826 ( 
.A(n_613),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_728),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_733),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_613),
.A2(n_341),
.B1(n_279),
.B2(n_291),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_733),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_641),
.B(n_294),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_634),
.B(n_208),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_737),
.B(n_314),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_641),
.B(n_319),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_732),
.B(n_478),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_737),
.B(n_326),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_723),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_712),
.Y(n_838)
);

BUFx12f_ASAP7_75t_SL g839 ( 
.A(n_613),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_708),
.B(n_329),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_644),
.B(n_347),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_749),
.A2(n_376),
.B1(n_350),
.B2(n_392),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_712),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_640),
.B(n_483),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_644),
.B(n_396),
.Y(n_845)
);

BUFx4_ASAP7_75t_L g846 ( 
.A(n_685),
.Y(n_846)
);

NOR2x1p5_ASAP7_75t_L g847 ( 
.A(n_730),
.B(n_344),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_642),
.B(n_209),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_720),
.B(n_397),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_640),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_646),
.B(n_649),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_604),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_620),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_646),
.B(n_403),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_699),
.B(n_296),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_721),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_723),
.B(n_484),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_649),
.B(n_297),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_699),
.B(n_304),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_604),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_306),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_699),
.B(n_308),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_643),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_657),
.B(n_312),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_620),
.Y(n_865)
);

NOR2x1_ASAP7_75t_L g866 ( 
.A(n_603),
.B(n_490),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_606),
.B(n_209),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_613),
.A2(n_322),
.B1(n_342),
.B2(n_339),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_636),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_721),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_L g871 ( 
.A(n_670),
.B(n_317),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_736),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_692),
.B(n_325),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_696),
.B(n_334),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_607),
.B(n_210),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_736),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_734),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_609),
.B(n_210),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_692),
.B(n_570),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_697),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_663),
.B(n_491),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_650),
.A2(n_365),
.B1(n_226),
.B2(n_228),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_697),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_636),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_706),
.B(n_570),
.Y(n_885)
);

INVxp33_ASAP7_75t_L g886 ( 
.A(n_682),
.Y(n_886)
);

AND2x2_ASAP7_75t_SL g887 ( 
.A(n_681),
.B(n_511),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_706),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_684),
.B(n_570),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_747),
.B(n_213),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_696),
.B(n_213),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_663),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_695),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_684),
.B(n_570),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_685),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_689),
.B(n_570),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_689),
.B(n_226),
.Y(n_897)
);

NAND2x1p5_ASAP7_75t_L g898 ( 
.A(n_731),
.B(n_511),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_695),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_628),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_663),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_616),
.B(n_570),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_698),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_637),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_686),
.B(n_570),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_637),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_731),
.B(n_228),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_679),
.B(n_232),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_668),
.B(n_232),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_679),
.B(n_238),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_670),
.A2(n_366),
.B1(n_405),
.B2(n_402),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_698),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_645),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_700),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_670),
.A2(n_366),
.B1(n_402),
.B2(n_399),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_668),
.B(n_238),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_668),
.B(n_239),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_663),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_645),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_668),
.B(n_239),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_680),
.B(n_343),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_604),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_668),
.B(n_343),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_780),
.Y(n_924)
);

NOR2x2_ASAP7_75t_L g925 ( 
.A(n_765),
.B(n_682),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_758),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_796),
.B(n_635),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_895),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_768),
.B(n_700),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_758),
.B(n_680),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_863),
.A2(n_738),
.B1(n_658),
.B2(n_664),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_768),
.A2(n_776),
.B1(n_803),
.B2(n_900),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_758),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_808),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_752),
.B(n_628),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_757),
.B(n_763),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_776),
.B(n_702),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_809),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_816),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_780),
.B(n_800),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_SL g941 ( 
.A1(n_886),
.A2(n_681),
.B1(n_727),
.B2(n_625),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_822),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_807),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_918),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_835),
.B(n_727),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_753),
.A2(n_738),
.B(n_693),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_758),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_827),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_852),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_758),
.B(n_683),
.Y(n_950)
);

AND3x1_ASAP7_75t_SL g951 ( 
.A(n_847),
.B(n_625),
.C(n_662),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_755),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_754),
.B(n_622),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_756),
.B(n_702),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_755),
.Y(n_955)
);

INVxp67_ASAP7_75t_L g956 ( 
.A(n_857),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_L g957 ( 
.A1(n_842),
.A2(n_647),
.B1(n_651),
.B2(n_667),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_790),
.B(n_623),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_828),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_789),
.B(n_705),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_758),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_830),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_842),
.A2(n_662),
.B1(n_670),
.B2(n_647),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_867),
.B(n_705),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_787),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_853),
.Y(n_966)
);

INVx1_ASAP7_75t_SL g967 ( 
.A(n_814),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_780),
.B(n_683),
.Y(n_968)
);

INVx6_ASAP7_75t_L g969 ( 
.A(n_757),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_753),
.A2(n_710),
.B(n_608),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_881),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_793),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_813),
.B(n_659),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_867),
.B(n_675),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_837),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_770),
.A2(n_742),
.B(n_651),
.C(n_746),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_865),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_780),
.B(n_693),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_875),
.B(n_675),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_803),
.B(n_782),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_893),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_899),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_852),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_869),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_884),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_903),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_912),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_914),
.Y(n_988)
);

INVx5_ASAP7_75t_L g989 ( 
.A(n_852),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_771),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_839),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_784),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_844),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_875),
.A2(n_658),
.B1(n_666),
.B2(n_664),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_878),
.B(n_678),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_825),
.B(n_661),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_878),
.B(n_678),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_825),
.A2(n_848),
.B1(n_832),
.B2(n_779),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_770),
.A2(n_742),
.B(n_750),
.C(n_744),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_880),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_883),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_760),
.B(n_832),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_918),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_782),
.B(n_729),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_888),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_848),
.B(n_666),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_904),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_852),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_775),
.B(n_648),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_792),
.B(n_648),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_906),
.Y(n_1011)
);

BUFx2_ASAP7_75t_L g1012 ( 
.A(n_877),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_913),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_919),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_838),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_860),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_819),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_887),
.A2(n_670),
.B1(n_750),
.B2(n_744),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_843),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_761),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_851),
.B(n_785),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_866),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_788),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_850),
.B(n_653),
.Y(n_1024)
);

OR2x2_ASAP7_75t_SL g1025 ( 
.A(n_766),
.B(n_438),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_856),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_870),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_807),
.Y(n_1028)
);

AND2x4_ASAP7_75t_L g1029 ( 
.A(n_872),
.B(n_674),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_876),
.B(n_653),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_840),
.A2(n_707),
.B1(n_670),
.B2(n_729),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_864),
.B(n_654),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_804),
.B(n_751),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_798),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_860),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_759),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_811),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_804),
.B(n_890),
.Y(n_1038)
);

NOR2x2_ASAP7_75t_L g1039 ( 
.A(n_887),
.B(n_369),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_807),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_812),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_820),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_772),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_860),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_911),
.A2(n_670),
.B1(n_751),
.B2(n_654),
.Y(n_1045)
);

CKINVDCx11_ASAP7_75t_R g1046 ( 
.A(n_846),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_840),
.A2(n_743),
.B1(n_729),
.B2(n_656),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_773),
.Y(n_1048)
);

AO22x1_ASAP7_75t_L g1049 ( 
.A1(n_890),
.A2(n_371),
.B1(n_395),
.B2(n_393),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_911),
.A2(n_656),
.B1(n_660),
.B2(n_601),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_858),
.B(n_660),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_860),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_778),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_R g1054 ( 
.A(n_806),
.B(n_345),
.Y(n_1054)
);

INVx1_ASAP7_75t_SL g1055 ( 
.A(n_892),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_800),
.B(n_743),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_901),
.B(n_352),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_891),
.B(n_897),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_826),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_907),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_922),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_781),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_922),
.B(n_743),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_891),
.B(n_352),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_873),
.B(n_602),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_849),
.A2(n_608),
.B1(n_710),
.B2(n_715),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_783),
.B(n_786),
.Y(n_1067)
);

AND2x6_ASAP7_75t_SL g1068 ( 
.A(n_909),
.B(n_353),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_897),
.B(n_353),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_L g1070 ( 
.A(n_826),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_922),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_795),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_916),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_917),
.Y(n_1074)
);

INVx3_ASAP7_75t_L g1075 ( 
.A(n_922),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_826),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_889),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_799),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_879),
.B(n_608),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_801),
.B(n_602),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_885),
.B(n_710),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_802),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_810),
.A2(n_600),
.B(n_601),
.C(n_725),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_849),
.A2(n_710),
.B1(n_715),
.B2(n_600),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_920),
.B(n_715),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_817),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_818),
.B(n_602),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_810),
.A2(n_722),
.B(n_735),
.C(n_725),
.Y(n_1088)
);

INVxp67_ASAP7_75t_SL g1089 ( 
.A(n_762),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_923),
.B(n_715),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_821),
.B(n_627),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_908),
.B(n_332),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_831),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_908),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_762),
.B(n_604),
.Y(n_1095)
);

INVx5_ASAP7_75t_L g1096 ( 
.A(n_764),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_834),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_764),
.A2(n_722),
.B1(n_735),
.B2(n_387),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_841),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_894),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_845),
.B(n_854),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_797),
.B(n_627),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_882),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_833),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_797),
.B(n_627),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_898),
.B(n_361),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_767),
.B(n_604),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_898),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_915),
.A2(n_383),
.B1(n_361),
.B2(n_367),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_910),
.Y(n_1110)
);

NOR3xp33_ASAP7_75t_SL g1111 ( 
.A(n_855),
.B(n_372),
.C(n_399),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_896),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_805),
.B(n_652),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_833),
.Y(n_1114)
);

AOI21x1_ASAP7_75t_L g1115 ( 
.A1(n_767),
.A2(n_652),
.B(n_717),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_769),
.A2(n_365),
.B1(n_387),
.B2(n_388),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_769),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_996),
.A2(n_915),
.B1(n_921),
.B2(n_910),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_949),
.A2(n_774),
.B(n_905),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1002),
.B(n_874),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_996),
.A2(n_774),
.B(n_815),
.C(n_805),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_962),
.Y(n_1122)
);

AO21x1_ASAP7_75t_L g1123 ( 
.A1(n_998),
.A2(n_815),
.B(n_836),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_967),
.B(n_829),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1038),
.B(n_868),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1036),
.B(n_777),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_962),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_932),
.B(n_836),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1043),
.B(n_791),
.Y(n_1129)
);

NAND2x1p5_ASAP7_75t_L g1130 ( 
.A(n_949),
.B(n_823),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_934),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_940),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1048),
.B(n_1062),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1072),
.B(n_1078),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_980),
.A2(n_921),
.B(n_874),
.C(n_794),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_963),
.A2(n_862),
.B1(n_861),
.B2(n_859),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1074),
.B(n_855),
.Y(n_1137)
);

AOI21xp33_ASAP7_75t_L g1138 ( 
.A1(n_957),
.A2(n_859),
.B(n_823),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1082),
.B(n_902),
.Y(n_1139)
);

NOR2x1_ASAP7_75t_SL g1140 ( 
.A(n_949),
.B(n_612),
.Y(n_1140)
);

O2A1O1Ixp5_ASAP7_75t_L g1141 ( 
.A1(n_1095),
.A2(n_824),
.B(n_652),
.C(n_655),
.Y(n_1141)
);

AOI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1092),
.A2(n_871),
.B(n_395),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_945),
.B(n_335),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1023),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_953),
.B(n_336),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_963),
.A2(n_383),
.B1(n_393),
.B2(n_389),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_949),
.A2(n_612),
.B(n_673),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1018),
.A2(n_382),
.B1(n_389),
.B2(n_373),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_953),
.B(n_971),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_989),
.A2(n_612),
.B(n_673),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1076),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1076),
.Y(n_1153)
);

NAND2xp33_ASAP7_75t_L g1154 ( 
.A(n_1096),
.B(n_612),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_989),
.A2(n_612),
.B(n_673),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_956),
.B(n_338),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_SL g1157 ( 
.A(n_1017),
.B(n_371),
.C(n_367),
.Y(n_1157)
);

AO21x1_ASAP7_75t_L g1158 ( 
.A1(n_1095),
.A2(n_1),
.B(n_2),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_941),
.A2(n_345),
.B1(n_364),
.B2(n_374),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_975),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_R g1161 ( 
.A(n_928),
.B(n_357),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_993),
.B(n_372),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_938),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_989),
.A2(n_701),
.B(n_676),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1023),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_952),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_952),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_955),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1086),
.B(n_655),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1076),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1018),
.A2(n_382),
.B1(n_373),
.B2(n_359),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_939),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_955),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_972),
.B(n_357),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_989),
.A2(n_701),
.B(n_676),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_1012),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_980),
.A2(n_717),
.B(n_704),
.C(n_691),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1107),
.A2(n_701),
.B(n_676),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_927),
.B(n_358),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_940),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1035),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_SL g1182 ( 
.A1(n_1085),
.A2(n_655),
.B(n_717),
.C(n_704),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1107),
.A2(n_673),
.B(n_701),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1096),
.A2(n_358),
.B1(n_359),
.B2(n_362),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1076),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1092),
.A2(n_704),
.B(n_691),
.C(n_364),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1096),
.A2(n_362),
.B1(n_374),
.B2(n_385),
.Y(n_1187)
);

INVx5_ASAP7_75t_SL g1188 ( 
.A(n_936),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_927),
.B(n_385),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_936),
.B(n_388),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1035),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_970),
.A2(n_673),
.B(n_701),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_1073),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_958),
.B(n_691),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_991),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1067),
.A2(n_676),
.B(n_158),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1101),
.A2(n_676),
.B(n_156),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_944),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_929),
.A2(n_154),
.B(n_198),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1096),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_937),
.A2(n_145),
.B(n_195),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1058),
.A2(n_741),
.B1(n_18),
.B2(n_20),
.Y(n_1202)
);

INVxp67_ASAP7_75t_L g1203 ( 
.A(n_1057),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1028),
.B(n_193),
.Y(n_1204)
);

CKINVDCx11_ASAP7_75t_R g1205 ( 
.A(n_1046),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1034),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_965),
.B(n_14),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_L g1208 ( 
.A(n_944),
.B(n_191),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_958),
.B(n_20),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1029),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1003),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1069),
.B(n_21),
.Y(n_1212)
);

INVx3_ASAP7_75t_SL g1213 ( 
.A(n_925),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1035),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_969),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_973),
.A2(n_184),
.B1(n_179),
.B2(n_177),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_942),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1029),
.B(n_171),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1093),
.A2(n_23),
.B(n_24),
.C(n_25),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1094),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1089),
.A2(n_168),
.B(n_163),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1003),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1032),
.A2(n_162),
.B(n_160),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1103),
.B(n_1021),
.Y(n_1224)
);

CKINVDCx14_ASAP7_75t_R g1225 ( 
.A(n_1046),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1068),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1097),
.A2(n_29),
.B(n_31),
.C(n_33),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1099),
.B(n_138),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_935),
.B(n_134),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1035),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1110),
.A2(n_37),
.B(n_40),
.C(n_42),
.Y(n_1231)
);

OAI22x1_ASAP7_75t_L g1232 ( 
.A1(n_1022),
.A2(n_1019),
.B1(n_1027),
.B2(n_1026),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_964),
.B(n_124),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_924),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1085),
.A2(n_122),
.B(n_112),
.C(n_109),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1060),
.B(n_37),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_969),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1006),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_948),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_974),
.B(n_108),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_1053),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_969),
.B(n_45),
.Y(n_1242)
);

AOI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1090),
.A2(n_102),
.B(n_96),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1055),
.B(n_45),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1033),
.B(n_95),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1065),
.A2(n_83),
.B(n_50),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_R g1247 ( 
.A(n_943),
.B(n_68),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1108),
.B(n_979),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_954),
.A2(n_49),
.B(n_51),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_995),
.B(n_49),
.Y(n_1250)
);

BUFx4_ASAP7_75t_SL g1251 ( 
.A(n_1028),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1025),
.Y(n_1252)
);

O2A1O1Ixp5_ASAP7_75t_L g1253 ( 
.A1(n_997),
.A2(n_53),
.B(n_55),
.C(n_56),
.Y(n_1253)
);

BUFx2_ASAP7_75t_L g1254 ( 
.A(n_925),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1040),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1090),
.A2(n_1115),
.B(n_978),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_999),
.A2(n_53),
.B(n_59),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1008),
.B(n_60),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1040),
.B(n_1059),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1104),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.Y(n_1260)
);

AO32x2_ASAP7_75t_L g1261 ( 
.A1(n_1098),
.A2(n_61),
.A3(n_67),
.B1(n_1116),
.B2(n_1071),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1030),
.A2(n_1015),
.B(n_1001),
.C(n_1005),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1051),
.A2(n_947),
.B(n_926),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1008),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_926),
.A2(n_947),
.B(n_961),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1000),
.A2(n_959),
.B(n_1024),
.C(n_1004),
.Y(n_1266)
);

BUFx12f_ASAP7_75t_L g1267 ( 
.A(n_1059),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1108),
.B(n_943),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1117),
.A2(n_1045),
.B1(n_976),
.B2(n_933),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_933),
.A2(n_961),
.B(n_930),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1070),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_981),
.Y(n_1272)
);

AND2x2_ASAP7_75t_SL g1273 ( 
.A(n_1070),
.B(n_1109),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_930),
.A2(n_950),
.B(n_1010),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1064),
.A2(n_951),
.B1(n_1114),
.B2(n_1106),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1004),
.A2(n_990),
.B(n_992),
.C(n_986),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1111),
.B(n_931),
.Y(n_1277)
);

AND3x1_ASAP7_75t_SL g1278 ( 
.A(n_951),
.B(n_1039),
.C(n_1049),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1071),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_SL g1280 ( 
.A(n_1117),
.B(n_924),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1054),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_982),
.B(n_987),
.Y(n_1282)
);

AO22x1_ASAP7_75t_L g1283 ( 
.A1(n_1117),
.A2(n_988),
.B1(n_1014),
.B2(n_1013),
.Y(n_1283)
);

AO21x1_ASAP7_75t_L g1284 ( 
.A1(n_1136),
.A2(n_1009),
.B(n_946),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1154),
.A2(n_1117),
.B(n_1091),
.Y(n_1285)
);

OA21x2_ASAP7_75t_L g1286 ( 
.A1(n_1121),
.A2(n_1080),
.B(n_1087),
.Y(n_1286)
);

AOI221xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1257),
.A2(n_1109),
.B1(n_976),
.B2(n_999),
.C(n_960),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1123),
.A2(n_994),
.B(n_1105),
.Y(n_1288)
);

AOI221x1_ASAP7_75t_L g1289 ( 
.A1(n_1257),
.A2(n_1112),
.B1(n_1113),
.B2(n_1102),
.C(n_1100),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1254),
.B(n_1041),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1138),
.A2(n_1056),
.B(n_1063),
.C(n_968),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1133),
.B(n_1077),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1138),
.A2(n_1083),
.B(n_1088),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1141),
.A2(n_1274),
.B(n_1240),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1152),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1160),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1152),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1126),
.A2(n_950),
.B(n_1056),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1126),
.A2(n_1081),
.B(n_1079),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1133),
.B(n_1077),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1271),
.B(n_1037),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1134),
.B(n_1100),
.Y(n_1302)
);

AO32x2_ASAP7_75t_L g1303 ( 
.A1(n_1269),
.A2(n_1050),
.A3(n_1045),
.B1(n_1054),
.B2(n_1031),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1134),
.B(n_1120),
.Y(n_1304)
);

INVx3_ASAP7_75t_L g1305 ( 
.A(n_1152),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1136),
.A2(n_1081),
.B(n_1079),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1269),
.A2(n_1061),
.A3(n_1044),
.B(n_1034),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1224),
.B(n_1042),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1182),
.A2(n_1186),
.B(n_1192),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1139),
.B(n_966),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1158),
.A2(n_1044),
.B(n_1061),
.Y(n_1311)
);

NAND3x1_ASAP7_75t_L g1312 ( 
.A(n_1209),
.B(n_1016),
.C(n_1075),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1139),
.B(n_966),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1150),
.B(n_977),
.Y(n_1314)
);

O2A1O1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1146),
.A2(n_968),
.B(n_978),
.C(n_1063),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1167),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1179),
.B(n_977),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1118),
.A2(n_1273),
.B1(n_1275),
.B2(n_1128),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1189),
.B(n_1143),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1263),
.A2(n_1112),
.B(n_984),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1256),
.A2(n_1011),
.B(n_984),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1270),
.A2(n_1265),
.B(n_1183),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1233),
.A2(n_985),
.A3(n_1007),
.B(n_1011),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1213),
.B(n_1156),
.Y(n_1324)
);

INVxp67_ASAP7_75t_SL g1325 ( 
.A(n_1173),
.Y(n_1325)
);

AND2x2_ASAP7_75t_SL g1326 ( 
.A(n_1260),
.B(n_1050),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1225),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1137),
.B(n_985),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1119),
.A2(n_1066),
.B(n_1084),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1128),
.B(n_1007),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_1161),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1233),
.A2(n_1047),
.B(n_1016),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1194),
.B(n_1075),
.Y(n_1333)
);

NOR2xp67_ASAP7_75t_L g1334 ( 
.A(n_1203),
.B(n_1124),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1122),
.B(n_983),
.Y(n_1335)
);

NAND3xp33_ASAP7_75t_SL g1336 ( 
.A(n_1159),
.B(n_1247),
.C(n_1207),
.Y(n_1336)
);

AO32x2_ASAP7_75t_L g1337 ( 
.A1(n_1200),
.A2(n_983),
.A3(n_1052),
.B1(n_1147),
.B2(n_1149),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1250),
.A2(n_1129),
.B1(n_1172),
.B2(n_1239),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1176),
.B(n_1052),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1202),
.A2(n_1220),
.B(n_1212),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1240),
.A2(n_1135),
.B(n_1125),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1232),
.A2(n_1250),
.A3(n_1197),
.B(n_1196),
.Y(n_1342)
);

OAI22x1_ASAP7_75t_L g1343 ( 
.A1(n_1277),
.A2(n_1236),
.B1(n_1210),
.B2(n_1190),
.Y(n_1343)
);

INVx1_ASAP7_75t_SL g1344 ( 
.A(n_1166),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1140),
.A2(n_1129),
.B(n_1283),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1248),
.A2(n_1228),
.B(n_1181),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1131),
.B(n_1163),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1235),
.A2(n_1178),
.B(n_1142),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1228),
.A2(n_1181),
.B(n_1266),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1181),
.A2(n_1262),
.B(n_1164),
.Y(n_1350)
);

BUFx4_ASAP7_75t_SL g1351 ( 
.A(n_1198),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1217),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1253),
.A2(n_1246),
.B(n_1201),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1177),
.A2(n_1243),
.B(n_1175),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1151),
.Y(n_1355)
);

AOI221x1_ASAP7_75t_L g1356 ( 
.A1(n_1142),
.A2(n_1200),
.B1(n_1249),
.B2(n_1227),
.C(n_1219),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1181),
.A2(n_1169),
.B(n_1229),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_SL g1358 ( 
.A1(n_1221),
.A2(n_1276),
.B(n_1199),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1169),
.A2(n_1130),
.B(n_1132),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1218),
.A2(n_1147),
.B1(n_1282),
.B2(n_1242),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1259),
.B(n_1268),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1193),
.B(n_1168),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1245),
.A2(n_1223),
.B(n_1216),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1144),
.B(n_1165),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1272),
.A2(n_1282),
.B1(n_1204),
.B2(n_1171),
.Y(n_1365)
);

AOI221xp5_ASAP7_75t_L g1366 ( 
.A1(n_1149),
.A2(n_1171),
.B1(n_1238),
.B2(n_1244),
.C(n_1174),
.Y(n_1366)
);

AO31x2_ASAP7_75t_L g1367 ( 
.A1(n_1231),
.A2(n_1187),
.A3(n_1184),
.B(n_1145),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_SL g1368 ( 
.A1(n_1204),
.A2(n_1259),
.B(n_1261),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1130),
.A2(n_1132),
.B(n_1180),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1153),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1153),
.Y(n_1371)
);

CKINVDCx8_ASAP7_75t_R g1372 ( 
.A(n_1241),
.Y(n_1372)
);

AND3x4_ASAP7_75t_L g1373 ( 
.A(n_1157),
.B(n_1255),
.C(n_1211),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1206),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1180),
.A2(n_1234),
.B(n_1264),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1188),
.B(n_1237),
.Y(n_1376)
);

AOI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1278),
.A2(n_1281),
.B1(n_1188),
.B2(n_1195),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1234),
.A2(n_1279),
.B(n_1264),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1222),
.Y(n_1379)
);

NAND2x1_ASAP7_75t_L g1380 ( 
.A(n_1280),
.B(n_1279),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1208),
.A2(n_1184),
.B(n_1187),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1258),
.A2(n_1230),
.B(n_1191),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1215),
.B(n_1188),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1191),
.A2(n_1230),
.B(n_1258),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1162),
.A2(n_1170),
.B(n_1261),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1251),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1185),
.B(n_1267),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1185),
.A2(n_1214),
.B(n_1261),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1214),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1185),
.Y(n_1390)
);

AOI221x1_ASAP7_75t_L g1391 ( 
.A1(n_1214),
.A2(n_1257),
.B1(n_1209),
.B2(n_1142),
.C(n_1138),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1252),
.B(n_1226),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_1181),
.B(n_1170),
.Y(n_1393)
);

AOI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1250),
.A2(n_1128),
.B(n_1233),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1123),
.A2(n_1269),
.A3(n_1136),
.B(n_1186),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1131),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1002),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1133),
.B(n_1002),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1263),
.A2(n_1256),
.B(n_1270),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1131),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1121),
.A2(n_1138),
.B(n_1136),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1263),
.A2(n_1256),
.B(n_1270),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1133),
.B(n_1002),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1160),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1002),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1121),
.A2(n_1138),
.B(n_1136),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1002),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1131),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1160),
.Y(n_1409)
);

NAND2x1_ASAP7_75t_L g1410 ( 
.A(n_1280),
.B(n_1008),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1121),
.A2(n_1138),
.B(n_1136),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1283),
.A2(n_1256),
.B(n_1136),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1224),
.A2(n_765),
.B1(n_996),
.B2(n_814),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1263),
.A2(n_1256),
.B(n_1270),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1121),
.A2(n_1138),
.B(n_1136),
.Y(n_1415)
);

NAND2x1p5_ASAP7_75t_L g1416 ( 
.A(n_1181),
.B(n_1170),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1127),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1160),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1209),
.A2(n_996),
.B(n_998),
.C(n_1146),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1131),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1002),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1263),
.A2(n_1256),
.B(n_1270),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1121),
.A2(n_1138),
.B(n_1136),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1205),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1160),
.Y(n_1425)
);

BUFx4_ASAP7_75t_SL g1426 ( 
.A(n_1271),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1143),
.B(n_945),
.Y(n_1427)
);

AOI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1002),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1131),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1143),
.B(n_945),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1224),
.B(n_814),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1127),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1133),
.B(n_1002),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1152),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1181),
.B(n_1170),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1209),
.A2(n_996),
.B(n_998),
.C(n_1146),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1152),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1131),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1002),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1127),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1271),
.B(n_1259),
.Y(n_1441)
);

NOR2xp67_ASAP7_75t_L g1442 ( 
.A(n_1203),
.B(n_928),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1214),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1143),
.B(n_945),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1133),
.B(n_1002),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1133),
.B(n_1002),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1133),
.B(n_1002),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1123),
.A2(n_1269),
.A3(n_1136),
.B(n_1186),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1443),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1319),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1344),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1351),
.Y(n_1452)
);

AO21x2_ASAP7_75t_L g1453 ( 
.A1(n_1401),
.A2(n_1411),
.B(n_1406),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1345),
.A2(n_1412),
.B(n_1349),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1366),
.A2(n_1318),
.B1(n_1326),
.B2(n_1336),
.Y(n_1455)
);

AO31x2_ASAP7_75t_L g1456 ( 
.A1(n_1391),
.A2(n_1284),
.A3(n_1289),
.B(n_1318),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1413),
.A2(n_1430),
.B1(n_1427),
.B2(n_1444),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1401),
.A2(n_1411),
.B(n_1406),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_SL g1459 ( 
.A1(n_1311),
.A2(n_1381),
.B(n_1382),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1360),
.A2(n_1431),
.B1(n_1381),
.B2(n_1447),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1446),
.A2(n_1317),
.B1(n_1423),
.B2(n_1415),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1422),
.A2(n_1322),
.B(n_1355),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1340),
.A2(n_1356),
.B(n_1308),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1344),
.Y(n_1465)
);

AOI221xp5_ASAP7_75t_L g1466 ( 
.A1(n_1340),
.A2(n_1423),
.B1(n_1415),
.B2(n_1343),
.C(n_1338),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1369),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1341),
.A2(n_1405),
.B(n_1397),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1354),
.A2(n_1320),
.B(n_1359),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1394),
.A2(n_1329),
.B(n_1350),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1341),
.A2(n_1306),
.B(n_1293),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1347),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1299),
.A2(n_1293),
.B(n_1298),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1426),
.Y(n_1474)
);

INVx4_ASAP7_75t_L g1475 ( 
.A(n_1443),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1287),
.A2(n_1421),
.B(n_1407),
.Y(n_1476)
);

O2A1O1Ixp33_ASAP7_75t_SL g1477 ( 
.A1(n_1398),
.A2(n_1445),
.B(n_1403),
.C(n_1433),
.Y(n_1477)
);

AO22x2_ASAP7_75t_L g1478 ( 
.A1(n_1338),
.A2(n_1365),
.B1(n_1385),
.B2(n_1358),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1398),
.B(n_1403),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1428),
.A2(n_1439),
.B(n_1285),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1417),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1346),
.A2(n_1388),
.B(n_1357),
.Y(n_1482)
);

AO31x2_ASAP7_75t_L g1483 ( 
.A1(n_1365),
.A2(n_1330),
.A3(n_1333),
.B(n_1313),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1393),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1348),
.A2(n_1309),
.B(n_1291),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1432),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1433),
.A2(n_1445),
.B(n_1304),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_L g1488 ( 
.A1(n_1304),
.A2(n_1339),
.B(n_1328),
.C(n_1290),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1294),
.A2(n_1384),
.B(n_1286),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1334),
.A2(n_1331),
.B1(n_1377),
.B2(n_1296),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1314),
.A2(n_1363),
.B1(n_1302),
.B2(n_1300),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1347),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1443),
.Y(n_1493)
);

OAI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1296),
.A2(n_1379),
.B1(n_1442),
.B2(n_1409),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1294),
.A2(n_1286),
.B(n_1330),
.Y(n_1495)
);

OA21x2_ASAP7_75t_L g1496 ( 
.A1(n_1287),
.A2(n_1333),
.B(n_1310),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1348),
.A2(n_1309),
.B(n_1332),
.Y(n_1497)
);

INVx8_ASAP7_75t_L g1498 ( 
.A(n_1443),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1379),
.A2(n_1404),
.B1(n_1314),
.B2(n_1418),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1332),
.A2(n_1363),
.B(n_1315),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1425),
.A2(n_1292),
.B1(n_1300),
.B2(n_1325),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1316),
.B(n_1324),
.Y(n_1502)
);

OAI221xp5_ASAP7_75t_L g1503 ( 
.A1(n_1362),
.A2(n_1383),
.B1(n_1372),
.B2(n_1392),
.C(n_1292),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1352),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1361),
.B(n_1376),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1297),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1441),
.Y(n_1507)
);

BUFx4f_ASAP7_75t_L g1508 ( 
.A(n_1373),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1310),
.A2(n_1313),
.B(n_1335),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1312),
.A2(n_1368),
.B(n_1353),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1393),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1353),
.A2(n_1288),
.B(n_1375),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1440),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1288),
.A2(n_1335),
.B(n_1410),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1396),
.A2(n_1420),
.B1(n_1400),
.B2(n_1408),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1424),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1416),
.Y(n_1517)
);

AND2x4_ASAP7_75t_SL g1518 ( 
.A(n_1361),
.B(n_1301),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1378),
.A2(n_1380),
.B(n_1364),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1301),
.Y(n_1520)
);

AO31x2_ASAP7_75t_L g1521 ( 
.A1(n_1395),
.A2(n_1448),
.A3(n_1307),
.B(n_1323),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1429),
.B(n_1438),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1364),
.A2(n_1374),
.B(n_1416),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1389),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1435),
.A2(n_1387),
.B(n_1437),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1435),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1390),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1307),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_SL g1529 ( 
.A1(n_1392),
.A2(n_1367),
.B(n_1337),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1295),
.A2(n_1370),
.B(n_1305),
.C(n_1437),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1295),
.A2(n_1371),
.B1(n_1370),
.B2(n_1305),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1303),
.A2(n_1342),
.B(n_1395),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1342),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1371),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1395),
.A2(n_1448),
.B(n_1337),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1297),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1303),
.A2(n_1434),
.B1(n_1327),
.B2(n_1337),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1367),
.B(n_1434),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1434),
.A2(n_1436),
.B1(n_1419),
.B2(n_1413),
.Y(n_1539)
);

INVx3_ASAP7_75t_L g1540 ( 
.A(n_1386),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1541)
);

A2O1A1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1257),
.C(n_996),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1427),
.B(n_1430),
.Y(n_1543)
);

CKINVDCx16_ASAP7_75t_R g1544 ( 
.A(n_1331),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_SL g1545 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1257),
.C(n_1366),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1386),
.Y(n_1546)
);

AOI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1345),
.A2(n_1412),
.B(n_1349),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1347),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1146),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1386),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1413),
.A2(n_765),
.B1(n_998),
.B2(n_965),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1401),
.A2(n_1411),
.B(n_1406),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1257),
.C(n_996),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1427),
.B(n_1430),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_765),
.C(n_996),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1316),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1347),
.Y(n_1562)
);

AOI21xp33_ASAP7_75t_L g1563 ( 
.A1(n_1419),
.A2(n_765),
.B(n_1146),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1347),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1443),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1397),
.A2(n_1407),
.B(n_1405),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1568)
);

BUFx10_ASAP7_75t_L g1569 ( 
.A(n_1386),
.Y(n_1569)
);

INVx3_ASAP7_75t_L g1570 ( 
.A(n_1369),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1347),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1321),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1443),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1419),
.B(n_1436),
.Y(n_1574)
);

CKINVDCx16_ASAP7_75t_R g1575 ( 
.A(n_1331),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1319),
.B(n_1427),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1347),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_SL g1578 ( 
.A1(n_1319),
.A2(n_765),
.B1(n_996),
.B2(n_941),
.Y(n_1578)
);

AO32x2_ASAP7_75t_L g1579 ( 
.A1(n_1318),
.A2(n_1338),
.A3(n_1365),
.B1(n_1200),
.B2(n_941),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1361),
.B(n_1382),
.Y(n_1580)
);

INVx4_ASAP7_75t_L g1581 ( 
.A(n_1443),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1347),
.Y(n_1582)
);

OAI21x1_ASAP7_75t_L g1583 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1583)
);

AOI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1345),
.A2(n_1412),
.B(n_1349),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1399),
.A2(n_1414),
.B(n_1402),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1404),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1347),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1369),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1419),
.B(n_1436),
.Y(n_1591)
);

AOI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1366),
.A2(n_1209),
.B1(n_941),
.B2(n_996),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1146),
.Y(n_1593)
);

AOI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1419),
.A2(n_765),
.B(n_1146),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_SL g1595 ( 
.A1(n_1345),
.A2(n_1158),
.B(n_1257),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1401),
.A2(n_1411),
.B(n_1406),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1319),
.B(n_1427),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1321),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1347),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1446),
.B(n_1447),
.Y(n_1600)
);

OA21x2_ASAP7_75t_L g1601 ( 
.A1(n_1401),
.A2(n_1411),
.B(n_1406),
.Y(n_1601)
);

O2A1O1Ixp5_ASAP7_75t_L g1602 ( 
.A1(n_1549),
.A2(n_1593),
.B(n_1542),
.C(n_1554),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1542),
.A2(n_1554),
.B(n_1591),
.C(n_1574),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1580),
.B(n_1518),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1543),
.B(n_1555),
.Y(n_1605)
);

O2A1O1Ixp5_ASAP7_75t_L g1606 ( 
.A1(n_1574),
.A2(n_1591),
.B(n_1468),
.C(n_1563),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1505),
.B(n_1576),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1597),
.B(n_1457),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1457),
.B(n_1578),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1450),
.B(n_1502),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1545),
.A2(n_1567),
.B(n_1487),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1587),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1527),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1592),
.A2(n_1455),
.B1(n_1461),
.B2(n_1503),
.Y(n_1614)
);

AOI21xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1557),
.A2(n_1600),
.B(n_1589),
.Y(n_1615)
);

O2A1O1Ixp33_ASAP7_75t_L g1616 ( 
.A1(n_1594),
.A2(n_1592),
.B(n_1545),
.C(n_1551),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1455),
.A2(n_1461),
.B1(n_1464),
.B2(n_1479),
.Y(n_1617)
);

OA22x2_ASAP7_75t_L g1618 ( 
.A1(n_1539),
.A2(n_1529),
.B1(n_1565),
.B2(n_1472),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1502),
.B(n_1451),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1462),
.A2(n_1508),
.B1(n_1490),
.B2(n_1494),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1462),
.A2(n_1508),
.B1(n_1499),
.B2(n_1466),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1546),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1492),
.B(n_1548),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1465),
.B(n_1520),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1562),
.B(n_1571),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1449),
.B(n_1573),
.Y(n_1627)
);

AOI21xp5_ASAP7_75t_L g1628 ( 
.A1(n_1477),
.A2(n_1471),
.B(n_1473),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1577),
.B(n_1582),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1527),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1507),
.B(n_1588),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1599),
.B(n_1488),
.Y(n_1632)
);

O2A1O1Ixp33_ASAP7_75t_L g1633 ( 
.A1(n_1595),
.A2(n_1501),
.B(n_1459),
.C(n_1561),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1470),
.A2(n_1495),
.B(n_1480),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1515),
.A2(n_1537),
.B1(n_1522),
.B2(n_1491),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1522),
.Y(n_1636)
);

AOI21x1_ASAP7_75t_SL g1637 ( 
.A1(n_1579),
.A2(n_1478),
.B(n_1544),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1481),
.B(n_1486),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1528),
.Y(n_1639)
);

AOI21x1_ASAP7_75t_SL g1640 ( 
.A1(n_1579),
.A2(n_1478),
.B(n_1575),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1513),
.B(n_1524),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1513),
.B(n_1515),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_R g1643 ( 
.A(n_1546),
.B(n_1550),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1534),
.B(n_1453),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1509),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1536),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1537),
.B(n_1506),
.Y(n_1647)
);

NOR2xp67_ASAP7_75t_L g1648 ( 
.A(n_1540),
.B(n_1452),
.Y(n_1648)
);

AOI221x1_ASAP7_75t_SL g1649 ( 
.A1(n_1531),
.A2(n_1596),
.B1(n_1458),
.B2(n_1456),
.C(n_1552),
.Y(n_1649)
);

AOI21x1_ASAP7_75t_SL g1650 ( 
.A1(n_1498),
.A2(n_1510),
.B(n_1547),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_SL g1651 ( 
.A1(n_1498),
.A2(n_1510),
.B(n_1454),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1532),
.A2(n_1512),
.B(n_1489),
.Y(n_1652)
);

OA21x2_ASAP7_75t_L g1653 ( 
.A1(n_1512),
.A2(n_1489),
.B(n_1469),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1491),
.A2(n_1523),
.B1(n_1493),
.B2(n_1511),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1475),
.A2(n_1581),
.B(n_1566),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1509),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1550),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1475),
.A2(n_1581),
.B(n_1566),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1483),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1493),
.A2(n_1484),
.B1(n_1511),
.B2(n_1517),
.Y(n_1660)
);

O2A1O1Ixp5_ASAP7_75t_L g1661 ( 
.A1(n_1584),
.A2(n_1533),
.B(n_1572),
.C(n_1598),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1509),
.B(n_1458),
.Y(n_1662)
);

O2A1O1Ixp5_ASAP7_75t_L g1663 ( 
.A1(n_1533),
.A2(n_1570),
.B(n_1467),
.C(n_1590),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1469),
.A2(n_1463),
.B(n_1460),
.Y(n_1664)
);

OA21x2_ASAP7_75t_L g1665 ( 
.A1(n_1463),
.A2(n_1568),
.B(n_1460),
.Y(n_1665)
);

AOI21x1_ASAP7_75t_SL g1666 ( 
.A1(n_1456),
.A2(n_1514),
.B(n_1530),
.Y(n_1666)
);

O2A1O1Ixp5_ASAP7_75t_L g1667 ( 
.A1(n_1533),
.A2(n_1570),
.B(n_1467),
.C(n_1590),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_L g1668 ( 
.A1(n_1552),
.A2(n_1601),
.B(n_1474),
.C(n_1540),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1526),
.B(n_1525),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1525),
.B(n_1540),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1526),
.A2(n_1601),
.B1(n_1552),
.B2(n_1566),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1569),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1526),
.B(n_1483),
.Y(n_1673)
);

OA21x2_ASAP7_75t_L g1674 ( 
.A1(n_1541),
.A2(n_1553),
.B(n_1585),
.Y(n_1674)
);

AND2x4_ASAP7_75t_L g1675 ( 
.A(n_1590),
.B(n_1467),
.Y(n_1675)
);

O2A1O1Ixp5_ASAP7_75t_L g1676 ( 
.A1(n_1570),
.A2(n_1456),
.B(n_1500),
.C(n_1485),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1496),
.A2(n_1476),
.B1(n_1516),
.B2(n_1535),
.Y(n_1677)
);

AOI21x1_ASAP7_75t_SL g1678 ( 
.A1(n_1569),
.A2(n_1521),
.B(n_1485),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1519),
.B(n_1483),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1483),
.B(n_1496),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1521),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1496),
.B(n_1535),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1521),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1535),
.B(n_1497),
.Y(n_1685)
);

INVx6_ASAP7_75t_L g1686 ( 
.A(n_1569),
.Y(n_1686)
);

NOR2xp67_ASAP7_75t_R g1687 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1558),
.A2(n_1559),
.B1(n_1560),
.B2(n_1564),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1583),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1556),
.B(n_1586),
.Y(n_1690)
);

OAI22xp5_ASAP7_75t_SL g1691 ( 
.A1(n_1578),
.A2(n_1592),
.B1(n_941),
.B2(n_1455),
.Y(n_1691)
);

NOR2xp67_ASAP7_75t_L g1692 ( 
.A(n_1503),
.B(n_1576),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1576),
.B(n_1597),
.Y(n_1693)
);

O2A1O1Ixp5_ASAP7_75t_L g1694 ( 
.A1(n_1549),
.A2(n_1593),
.B(n_1554),
.C(n_1542),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1567),
.A2(n_1470),
.B(n_1468),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1543),
.B(n_1555),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1556),
.B(n_1586),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1592),
.A2(n_1419),
.B1(n_1436),
.B2(n_1413),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1543),
.B(n_1555),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1546),
.Y(n_1700)
);

AND2x2_ASAP7_75t_SL g1701 ( 
.A(n_1574),
.B(n_1591),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1567),
.A2(n_1470),
.B(n_1468),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1543),
.B(n_1555),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1592),
.A2(n_1419),
.B1(n_1436),
.B2(n_1413),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1546),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1504),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1574),
.B(n_1591),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1625),
.B(n_1673),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1670),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1625),
.B(n_1644),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1662),
.B(n_1659),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1611),
.A2(n_1707),
.B(n_1701),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1642),
.Y(n_1713)
);

AOI21x1_ASAP7_75t_L g1714 ( 
.A1(n_1688),
.A2(n_1677),
.B(n_1628),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1639),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1659),
.B(n_1680),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1663),
.A2(n_1667),
.B(n_1651),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1636),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1625),
.B(n_1644),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1675),
.B(n_1679),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1701),
.B(n_1707),
.Y(n_1721)
);

INVxp67_ASAP7_75t_R g1722 ( 
.A(n_1610),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1690),
.B(n_1697),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1645),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1656),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1685),
.B(n_1681),
.Y(n_1726)
);

OAI21x1_ASAP7_75t_L g1727 ( 
.A1(n_1663),
.A2(n_1667),
.B(n_1650),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1681),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1602),
.A2(n_1694),
.B(n_1606),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1619),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1683),
.B(n_1682),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1706),
.B(n_1608),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1675),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1624),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1638),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1615),
.B(n_1607),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1647),
.B(n_1618),
.Y(n_1738)
);

INVx2_ASAP7_75t_SL g1739 ( 
.A(n_1686),
.Y(n_1739)
);

AOI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1689),
.A2(n_1614),
.B(n_1617),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1618),
.B(n_1604),
.Y(n_1741)
);

INVx8_ASAP7_75t_L g1742 ( 
.A(n_1627),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1605),
.B(n_1696),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1668),
.B(n_1684),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1602),
.A2(n_1694),
.B(n_1704),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1603),
.B(n_1641),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1691),
.A2(n_1698),
.B1(n_1621),
.B2(n_1620),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1699),
.B(n_1703),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1623),
.Y(n_1749)
);

BUFx5_ASAP7_75t_L g1750 ( 
.A(n_1684),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1626),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1629),
.Y(n_1752)
);

BUFx3_ASAP7_75t_L g1753 ( 
.A(n_1613),
.Y(n_1753)
);

OAI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1676),
.A2(n_1661),
.B(n_1666),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1609),
.B(n_1702),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1632),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1612),
.Y(n_1757)
);

OAI21x1_ASAP7_75t_L g1758 ( 
.A1(n_1653),
.A2(n_1678),
.B(n_1664),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1649),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1652),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1652),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1634),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1692),
.B(n_1631),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_1735),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1755),
.B(n_1709),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1762),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1711),
.B(n_1702),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1755),
.B(n_1702),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1724),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1724),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

AOI222xp33_ASAP7_75t_L g1772 ( 
.A1(n_1747),
.A2(n_1635),
.B1(n_1616),
.B2(n_1672),
.C1(n_1648),
.C2(n_1654),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1711),
.B(n_1695),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1742),
.Y(n_1774)
);

AO21x2_ASAP7_75t_L g1775 ( 
.A1(n_1714),
.A2(n_1633),
.B(n_1687),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1760),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1726),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1761),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1761),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1709),
.B(n_1634),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1756),
.B(n_1653),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1759),
.B(n_1664),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1759),
.B(n_1664),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1731),
.B(n_1674),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1716),
.B(n_1660),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1728),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1716),
.B(n_1665),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1750),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1777),
.B(n_1719),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1769),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1769),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1769),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1785),
.B(n_1732),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1777),
.Y(n_1794)
);

OA21x2_ASAP7_75t_L g1795 ( 
.A1(n_1776),
.A2(n_1758),
.B(n_1717),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1776),
.Y(n_1796)
);

AOI31xp33_ASAP7_75t_L g1797 ( 
.A1(n_1772),
.A2(n_1712),
.A3(n_1745),
.B(n_1721),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1765),
.B(n_1710),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1772),
.A2(n_1721),
.B(n_1729),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1770),
.Y(n_1800)
);

OAI33xp33_ASAP7_75t_L g1801 ( 
.A1(n_1782),
.A2(n_1783),
.A3(n_1785),
.B1(n_1781),
.B2(n_1787),
.B3(n_1773),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1778),
.Y(n_1802)
);

AOI31xp33_ASAP7_75t_L g1803 ( 
.A1(n_1772),
.A2(n_1737),
.A3(n_1763),
.B(n_1738),
.Y(n_1803)
);

OAI211xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1781),
.A2(n_1723),
.B(n_1757),
.C(n_1730),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1774),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1777),
.A2(n_1744),
.B1(n_1738),
.B2(n_1746),
.C(n_1733),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1781),
.B(n_1719),
.Y(n_1807)
);

AOI33xp33_ASAP7_75t_L g1808 ( 
.A1(n_1768),
.A2(n_1746),
.A3(n_1749),
.B1(n_1751),
.B2(n_1752),
.B3(n_1748),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1771),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1764),
.A2(n_1722),
.B1(n_1741),
.B2(n_1740),
.Y(n_1810)
);

INVx5_ASAP7_75t_L g1811 ( 
.A(n_1788),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1775),
.A2(n_1658),
.B(n_1655),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1767),
.A2(n_1740),
.B1(n_1739),
.B2(n_1718),
.C(n_1744),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1767),
.B(n_1733),
.Y(n_1814)
);

OAI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1767),
.A2(n_1739),
.B1(n_1744),
.B2(n_1686),
.C(n_1713),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1765),
.B(n_1780),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1764),
.A2(n_1741),
.B1(n_1710),
.B2(n_1720),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1765),
.B(n_1722),
.Y(n_1818)
);

AOI322xp5_ASAP7_75t_L g1819 ( 
.A1(n_1768),
.A2(n_1748),
.A3(n_1743),
.B1(n_1708),
.B2(n_1640),
.C1(n_1637),
.C2(n_1715),
.Y(n_1819)
);

OR2x6_ASAP7_75t_L g1820 ( 
.A(n_1774),
.B(n_1742),
.Y(n_1820)
);

NOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1783),
.B(n_1753),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1773),
.A2(n_1744),
.B1(n_1686),
.B2(n_1734),
.C(n_1753),
.Y(n_1822)
);

BUFx3_ASAP7_75t_L g1823 ( 
.A(n_1774),
.Y(n_1823)
);

NAND4xp25_ASAP7_75t_L g1824 ( 
.A(n_1768),
.B(n_1736),
.C(n_1646),
.D(n_1630),
.Y(n_1824)
);

AND2x6_ASAP7_75t_SL g1825 ( 
.A(n_1820),
.B(n_1643),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1821),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1790),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1811),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1820),
.Y(n_1829)
);

INVx2_ASAP7_75t_SL g1830 ( 
.A(n_1811),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1816),
.B(n_1765),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1808),
.B(n_1786),
.Y(n_1832)
);

BUFx3_ASAP7_75t_L g1833 ( 
.A(n_1805),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1796),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1794),
.Y(n_1835)
);

AOI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1812),
.A2(n_1779),
.B(n_1766),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1790),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1791),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1791),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1792),
.Y(n_1840)
);

INVx4_ASAP7_75t_SL g1841 ( 
.A(n_1820),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1792),
.Y(n_1842)
);

OAI21x1_ASAP7_75t_L g1843 ( 
.A1(n_1795),
.A2(n_1727),
.B(n_1754),
.Y(n_1843)
);

INVx1_ASAP7_75t_SL g1844 ( 
.A(n_1789),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1800),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1793),
.B(n_1786),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1816),
.B(n_1780),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1803),
.B(n_1774),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1814),
.B(n_1784),
.Y(n_1849)
);

BUFx2_ASAP7_75t_L g1850 ( 
.A(n_1820),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1811),
.Y(n_1851)
);

OR2x6_ASAP7_75t_L g1852 ( 
.A(n_1810),
.B(n_1774),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1798),
.B(n_1780),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1827),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1841),
.B(n_1818),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1827),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1841),
.B(n_1818),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1851),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1841),
.B(n_1798),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1834),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1829),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1837),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1835),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1832),
.B(n_1799),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1837),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1838),
.Y(n_1866)
);

OA21x2_ASAP7_75t_L g1867 ( 
.A1(n_1843),
.A2(n_1779),
.B(n_1802),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1832),
.B(n_1814),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1838),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1841),
.B(n_1807),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1839),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1834),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1848),
.A2(n_1804),
.B1(n_1801),
.B2(n_1824),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1841),
.B(n_1807),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1829),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1844),
.B(n_1789),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1841),
.B(n_1811),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1850),
.B(n_1811),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1844),
.B(n_1797),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1850),
.B(n_1780),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1846),
.B(n_1819),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1846),
.B(n_1817),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1839),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1849),
.B(n_1806),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_1852),
.B(n_1813),
.C(n_1815),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1831),
.B(n_1805),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1852),
.B(n_1784),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1833),
.B(n_1809),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1828),
.B(n_1823),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1852),
.B(n_1784),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1840),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_SL g1892 ( 
.A(n_1826),
.B(n_1822),
.C(n_1643),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1840),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1842),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1833),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1831),
.B(n_1823),
.Y(n_1896)
);

AO22x1_ASAP7_75t_L g1897 ( 
.A1(n_1879),
.A2(n_1826),
.B1(n_1833),
.B2(n_1851),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1864),
.A2(n_1852),
.B(n_1836),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1854),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1854),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1873),
.B(n_1853),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1856),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1868),
.B(n_1852),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1856),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1892),
.B(n_1622),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1875),
.B(n_1853),
.Y(n_1906)
);

HB1xp67_ASAP7_75t_L g1907 ( 
.A(n_1863),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1859),
.B(n_1852),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1895),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1861),
.B(n_1853),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1862),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_1889),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1862),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1865),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1865),
.Y(n_1915)
);

BUFx2_ASAP7_75t_SL g1916 ( 
.A(n_1877),
.Y(n_1916)
);

NOR2xp33_ASAP7_75t_L g1917 ( 
.A(n_1882),
.B(n_1622),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1876),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1868),
.B(n_1842),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1860),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1860),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1881),
.B(n_1831),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1866),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1859),
.B(n_1855),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1888),
.B(n_1847),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1872),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1867),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1855),
.B(n_1847),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1866),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1884),
.B(n_1847),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1884),
.B(n_1845),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1857),
.B(n_1828),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1857),
.B(n_1828),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1918),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1916),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1916),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1912),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1912),
.Y(n_1938)
);

OAI21xp33_ASAP7_75t_L g1939 ( 
.A1(n_1901),
.A2(n_1885),
.B(n_1874),
.Y(n_1939)
);

INVx1_ASAP7_75t_SL g1940 ( 
.A(n_1924),
.Y(n_1940)
);

INVxp67_ASAP7_75t_SL g1941 ( 
.A(n_1907),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1924),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1899),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1932),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1932),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1930),
.B(n_1922),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1917),
.B(n_1657),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1928),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1899),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1928),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1933),
.B(n_1889),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1931),
.B(n_1919),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1933),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1909),
.B(n_1896),
.Y(n_1954)
);

INVx2_ASAP7_75t_SL g1955 ( 
.A(n_1908),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1908),
.Y(n_1956)
);

INVxp67_ASAP7_75t_L g1957 ( 
.A(n_1905),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1900),
.Y(n_1958)
);

CKINVDCx16_ASAP7_75t_R g1959 ( 
.A(n_1903),
.Y(n_1959)
);

NAND3xp33_ASAP7_75t_SL g1960 ( 
.A(n_1898),
.B(n_1874),
.C(n_1870),
.Y(n_1960)
);

OR2x2_ASAP7_75t_L g1961 ( 
.A(n_1919),
.B(n_1876),
.Y(n_1961)
);

AOI222xp33_ASAP7_75t_L g1962 ( 
.A1(n_1939),
.A2(n_1960),
.B1(n_1941),
.B2(n_1957),
.C1(n_1934),
.C2(n_1898),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1934),
.B(n_1929),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1940),
.B(n_1942),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1938),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1946),
.B(n_1906),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1938),
.Y(n_1967)
);

O2A1O1Ixp33_ASAP7_75t_L g1968 ( 
.A1(n_1935),
.A2(n_1936),
.B(n_1952),
.C(n_1937),
.Y(n_1968)
);

AO21x1_ASAP7_75t_L g1969 ( 
.A1(n_1937),
.A2(n_1902),
.B(n_1900),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1953),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1953),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1943),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1951),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1955),
.A2(n_1870),
.B1(n_1897),
.B2(n_1910),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1943),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1951),
.B(n_1886),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1949),
.Y(n_1977)
);

OAI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1956),
.A2(n_1903),
.B(n_1925),
.Y(n_1978)
);

AND2x4_ASAP7_75t_SL g1979 ( 
.A(n_1955),
.B(n_1877),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1947),
.B(n_1954),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1959),
.B(n_1889),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1944),
.A2(n_1897),
.B1(n_1878),
.B2(n_1886),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1979),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1970),
.Y(n_1984)
);

NOR2xp33_ASAP7_75t_L g1985 ( 
.A(n_1980),
.B(n_1946),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1965),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1971),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1967),
.B(n_1945),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1973),
.B(n_1948),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1969),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1964),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1964),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1972),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1962),
.B(n_1952),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1968),
.B(n_1948),
.Y(n_1995)
);

AOI322xp5_ASAP7_75t_L g1996 ( 
.A1(n_1994),
.A2(n_1981),
.A3(n_1978),
.B1(n_1982),
.B2(n_1974),
.C1(n_1963),
.C2(n_1975),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1983),
.B(n_1962),
.Y(n_1997)
);

NAND3xp33_ASAP7_75t_L g1998 ( 
.A(n_1994),
.B(n_1968),
.C(n_1963),
.Y(n_1998)
);

AOI21x1_ASAP7_75t_L g1999 ( 
.A1(n_1990),
.A2(n_1977),
.B(n_1958),
.Y(n_1999)
);

AOI222xp33_ASAP7_75t_L g2000 ( 
.A1(n_1995),
.A2(n_1950),
.B1(n_1949),
.B2(n_1958),
.C1(n_1976),
.C2(n_1915),
.Y(n_2000)
);

OAI211xp5_ASAP7_75t_L g2001 ( 
.A1(n_1985),
.A2(n_1988),
.B(n_1983),
.C(n_1987),
.Y(n_2001)
);

NOR2xp67_ASAP7_75t_L g2002 ( 
.A(n_1991),
.B(n_1961),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1985),
.A2(n_1966),
.B(n_1961),
.Y(n_2003)
);

OAI21xp33_ASAP7_75t_L g2004 ( 
.A1(n_1986),
.A2(n_1950),
.B(n_1904),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1989),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_L g2006 ( 
.A(n_1992),
.B(n_1657),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1984),
.A2(n_1920),
.B1(n_1926),
.B2(n_1921),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_2002),
.B(n_1993),
.Y(n_2008)
);

NAND4xp25_ASAP7_75t_L g2009 ( 
.A(n_1996),
.B(n_1929),
.C(n_1914),
.D(n_1913),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1997),
.Y(n_2010)
);

AOI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_1998),
.A2(n_1904),
.B1(n_1915),
.B2(n_1923),
.C(n_1914),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_2001),
.B(n_1700),
.Y(n_2012)
);

AOI211xp5_ASAP7_75t_SL g2013 ( 
.A1(n_2004),
.A2(n_1902),
.B(n_1911),
.C(n_1913),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_2003),
.B(n_1896),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_2006),
.A2(n_2005),
.B1(n_2000),
.B2(n_2007),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1999),
.Y(n_2016)
);

NOR3xp33_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_1705),
.C(n_1911),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_2008),
.B(n_1878),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2014),
.B(n_1923),
.Y(n_2019)
);

NOR2x1_ASAP7_75t_L g2020 ( 
.A(n_2016),
.B(n_1858),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2015),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2009),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2011),
.Y(n_2023)
);

HB1xp67_ASAP7_75t_L g2024 ( 
.A(n_2012),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2013),
.Y(n_2025)
);

NAND2xp33_ASAP7_75t_SL g2026 ( 
.A(n_2025),
.B(n_1858),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_2018),
.Y(n_2027)
);

AOI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_2021),
.A2(n_1858),
.B1(n_1926),
.B2(n_1921),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_R g2029 ( 
.A(n_2022),
.B(n_1825),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_2018),
.Y(n_2030)
);

NOR2x1_ASAP7_75t_L g2031 ( 
.A(n_2020),
.B(n_2023),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2030),
.Y(n_2032)
);

NOR4xp25_ASAP7_75t_L g2033 ( 
.A(n_2027),
.B(n_2019),
.C(n_2024),
.D(n_2017),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_L g2034 ( 
.A(n_2031),
.B(n_1920),
.Y(n_2034)
);

NAND3xp33_ASAP7_75t_SL g2035 ( 
.A(n_2033),
.B(n_2029),
.C(n_2026),
.Y(n_2035)
);

AOI322xp5_ASAP7_75t_L g2036 ( 
.A1(n_2035),
.A2(n_2032),
.A3(n_2034),
.B1(n_2028),
.B2(n_1927),
.C1(n_1880),
.C2(n_1830),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2036),
.B(n_1872),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_2036),
.Y(n_2038)
);

AOI22xp33_ASAP7_75t_SL g2039 ( 
.A1(n_2038),
.A2(n_1927),
.B1(n_1851),
.B2(n_1830),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_2037),
.B(n_1887),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2040),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2039),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_2042),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2043),
.B(n_2041),
.Y(n_2044)
);

AOI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_2044),
.A2(n_1927),
.B1(n_1851),
.B2(n_1830),
.Y(n_2045)
);

AOI322xp5_ASAP7_75t_L g2046 ( 
.A1(n_2045),
.A2(n_1891),
.A3(n_1869),
.B1(n_1883),
.B2(n_1893),
.C1(n_1871),
.C2(n_1894),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_2046),
.A2(n_1880),
.B1(n_1883),
.B2(n_1869),
.Y(n_2047)
);

AOI211xp5_ASAP7_75t_L g2048 ( 
.A1(n_2047),
.A2(n_1890),
.B(n_1887),
.C(n_1613),
.Y(n_2048)
);


endmodule