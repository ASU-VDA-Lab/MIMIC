module real_jpeg_28336_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_2),
.B(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_2),
.B(n_10),
.Y(n_15)
);

OAI221xp5_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_8),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_7)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_24),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_13),
.CON(n_12),
.SN(n_12)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_23),
.Y(n_29)
);

NOR3xp33_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_21),
.C(n_30),
.Y(n_6)
);

OAI22xp33_ASAP7_75t_L g21 ( 
.A1(n_8),
.A2(n_15),
.B1(n_22),
.B2(n_28),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_10),
.A2(n_11),
.B1(n_17),
.B2(n_19),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_11),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_11),
.Y(n_10)
);

CKINVDCx5p33_ASAP7_75t_R g11 ( 
.A(n_12),
.Y(n_11)
);

BUFx24_ASAP7_75t_SL g34 ( 
.A(n_12),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_18),
.Y(n_17)
);

OR2x2_ASAP7_75t_SL g20 ( 
.A(n_14),
.B(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);


endmodule