module fake_jpeg_19419_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_25),
.B1(n_19),
.B2(n_33),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_16),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_49),
.B(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_25),
.B1(n_19),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_25),
.B1(n_33),
.B2(n_28),
.Y(n_51)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_22),
.Y(n_73)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_34),
.B1(n_16),
.B2(n_29),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_68),
.B1(n_29),
.B2(n_32),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_32),
.B(n_17),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_26),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_35),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_71),
.B(n_74),
.Y(n_131)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_32),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_75),
.A2(n_86),
.B1(n_100),
.B2(n_30),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_55),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_76),
.B(n_84),
.Y(n_114)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_81),
.B(n_92),
.Y(n_117)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_40),
.B1(n_39),
.B2(n_31),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_102),
.B1(n_111),
.B2(n_52),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_22),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_89),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_39),
.B1(n_40),
.B2(n_31),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_95),
.Y(n_123)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_63),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_90),
.B(n_94),
.Y(n_133)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_59),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_30),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_108),
.C(n_23),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_31),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_98),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_60),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_52),
.A2(n_26),
.B1(n_12),
.B2(n_15),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_53),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_106),
.B1(n_107),
.B2(n_21),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_51),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_12),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_12),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_67),
.B(n_53),
.Y(n_108)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_52),
.B1(n_58),
.B2(n_50),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_113),
.A2(n_118),
.B1(n_132),
.B2(n_134),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_116),
.B1(n_86),
.B2(n_125),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_26),
.B1(n_23),
.B2(n_15),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_116),
.A2(n_125),
.B1(n_100),
.B2(n_76),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_89),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_23),
.B1(n_14),
.B2(n_13),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_127),
.B(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_85),
.A2(n_24),
.B1(n_21),
.B2(n_18),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_88),
.A2(n_24),
.B1(n_18),
.B2(n_2),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_69),
.B1(n_110),
.B2(n_78),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_18),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_146),
.B1(n_151),
.B2(n_159),
.Y(n_186)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_155),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_157),
.B(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_115),
.A2(n_81),
.B1(n_75),
.B2(n_71),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_111),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_152),
.Y(n_190)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_149),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_97),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_101),
.C(n_93),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_168),
.C(n_120),
.Y(n_176)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_101),
.B(n_93),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_136),
.A2(n_79),
.B1(n_80),
.B2(n_104),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_95),
.B1(n_108),
.B2(n_94),
.Y(n_159)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_161),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_90),
.A3(n_99),
.B1(n_91),
.B2(n_87),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_69),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_139),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_90),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_14),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_165),
.B(n_173),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_166),
.A2(n_167),
.B1(n_174),
.B2(n_133),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_77),
.B1(n_72),
.B2(n_82),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_87),
.C(n_109),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_172),
.B1(n_120),
.B2(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

AND2x4_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_0),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_113),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_114),
.B(n_1),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_138),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_133),
.B1(n_118),
.B2(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_201),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_153),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_206),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_112),
.C(n_119),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_203),
.C(n_174),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_168),
.Y(n_183)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_191),
.B1(n_151),
.B2(n_169),
.Y(n_219)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_188),
.Y(n_222)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_134),
.B1(n_141),
.B2(n_126),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_194),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_129),
.B1(n_126),
.B2(n_121),
.Y(n_196)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_171),
.B(n_129),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_171),
.B(n_145),
.Y(n_211)
);

BUFx24_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g228 ( 
.A(n_200),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_142),
.B(n_139),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_156),
.B(n_159),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_121),
.C(n_5),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_4),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_204),
.B(n_10),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_195),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_224),
.C(n_231),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_211),
.A2(n_216),
.B(n_199),
.Y(n_255)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_196),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_145),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_220),
.Y(n_250)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_227),
.B1(n_191),
.B2(n_221),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_201),
.Y(n_223)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_223),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_150),
.C(n_5),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_4),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_225),
.B(n_226),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_177),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_6),
.C(n_7),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_6),
.C(n_7),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_203),
.C(n_182),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_202),
.B(n_180),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_243),
.B(n_248),
.C(n_228),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_232),
.A2(n_212),
.B1(n_217),
.B2(n_186),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_241),
.A2(n_249),
.B1(n_234),
.B2(n_228),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_246),
.B1(n_256),
.B2(n_234),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_233),
.A2(n_184),
.B(n_197),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_184),
.B1(n_196),
.B2(n_175),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_247),
.B(n_254),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_196),
.B(n_175),
.C(n_193),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_190),
.B1(n_178),
.B2(n_181),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_216),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_211),
.B(n_193),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_230),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_245),
.B1(n_248),
.B2(n_228),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_225),
.A2(n_190),
.B1(n_199),
.B2(n_198),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_189),
.C(n_179),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_244),
.C(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_253),
.Y(n_260)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_215),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_213),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_264),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_220),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_268),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_271),
.C(n_275),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_274),
.B(n_243),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_223),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_235),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_270),
.Y(n_278)
);

OAI21x1_ASAP7_75t_L g270 ( 
.A1(n_236),
.A2(n_213),
.B(n_222),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_222),
.C(n_230),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_246),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_240),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_231),
.C(n_208),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_255),
.B(n_256),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_218),
.B1(n_215),
.B2(n_226),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_274),
.B(n_283),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_260),
.B1(n_248),
.B2(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_266),
.C(n_265),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_291),
.C(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_285),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_268),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_242),
.C(n_252),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_248),
.C(n_192),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_267),
.B(n_277),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_261),
.C(n_8),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_287),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_261),
.B(n_8),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_278),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_293),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_308),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_291),
.B1(n_292),
.B2(n_280),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_278),
.B1(n_288),
.B2(n_294),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_300),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NOR2x1p5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_305),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_318),
.A2(n_299),
.B(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_297),
.C(n_280),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_301),
.B(n_306),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_322),
.A2(n_323),
.B(n_320),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_315),
.A2(n_307),
.B(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_309),
.C(n_314),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_325),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_326),
.B1(n_318),
.B2(n_321),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI221xp5_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_296),
.B1(n_286),
.B2(n_10),
.C(n_9),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_7),
.B(n_10),
.Y(n_331)
);


endmodule