module fake_ibex_1710_n_4658 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4658);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4658;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_3548;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_873;
wire n_962;
wire n_4632;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_3838;
wire n_957;
wire n_4514;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4353;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4343;
wire n_4648;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_4142;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3411;
wire n_3025;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_963;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_875;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4445;
wire n_876;
wire n_3211;
wire n_3479;
wire n_1840;
wire n_2837;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_3392;
wire n_1937;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_4447;
wire n_4491;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2846;
wire n_2685;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_4312;
wire n_4567;
wire n_917;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_4014;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1960;
wire n_1723;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3910;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3769;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_971;
wire n_4444;
wire n_1350;
wire n_3627;
wire n_906;
wire n_4499;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_3199;
wire n_1616;
wire n_2723;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_3217;
wire n_2511;
wire n_2782;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_4505;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_4615;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3963;
wire n_3800;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4549;
wire n_4573;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4523;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_4571;
wire n_959;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4501;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_4403;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_965;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_3082;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4485;
wire n_4608;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2910;
wire n_2552;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_4500;
wire n_4559;
wire n_998;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1400;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_2842;
wire n_2711;
wire n_3477;
wire n_3070;
wire n_3646;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_3557;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1185;
wire n_1683;
wire n_4256;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_3252;
wire n_2696;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_961;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_2127;
wire n_3735;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1601;
wire n_1294;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3673;
wire n_3476;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3269;
wire n_3029;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_4007;
wire n_3960;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1962;
wire n_1225;
wire n_2346;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3912;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_4638;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_3899;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_4637;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_3746;
wire n_2758;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2984;
wire n_2732;
wire n_3162;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2251;
wire n_2012;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_3229;
wire n_2225;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1989;
wire n_1740;
wire n_3604;
wire n_1838;
wire n_3649;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4162;
wire n_4111;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_4611;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_3368;
wire n_3561;
wire n_956;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_4562;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3972;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1366;
wire n_1518;
wire n_4380;
wire n_4350;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3173;
wire n_2653;
wire n_2872;
wire n_3102;
wire n_4281;
wire n_4345;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_4045;
wire n_854;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1912;
wire n_1297;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_3296;
wire n_1911;
wire n_2293;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_980;
wire n_849;
wire n_1193;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_1074;
wire n_3225;
wire n_3380;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_4412;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_4560;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1027;
wire n_1516;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2855;
wire n_2618;
wire n_2357;
wire n_4448;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_4544;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2961;
wire n_2770;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_4589;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_2619;
wire n_3873;
wire n_3738;
wire n_4506;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4251;
wire n_4106;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_856;
wire n_3193;
wire n_4534;
wire n_3635;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1678;
wire n_1091;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2673;
wire n_2676;
wire n_921;
wire n_2430;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

INVx1_ASAP7_75t_L g840 ( 
.A(n_495),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_136),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_742),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_213),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_702),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_239),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_639),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_392),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_381),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_492),
.Y(n_849)
);

HB1xp67_ASAP7_75t_L g850 ( 
.A(n_771),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_517),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_545),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_339),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_134),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_397),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_807),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_685),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_373),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_511),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_776),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_191),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_331),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_171),
.Y(n_863)
);

BUFx2_ASAP7_75t_SL g864 ( 
.A(n_328),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_567),
.Y(n_865)
);

BUFx10_ASAP7_75t_L g866 ( 
.A(n_767),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_233),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_640),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_360),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_791),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_668),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_323),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_300),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_772),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_469),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_421),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_351),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_482),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_790),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_269),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_806),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_68),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_260),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_297),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_710),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_239),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_787),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_67),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_551),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_663),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_94),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_537),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_761),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_521),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_682),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_700),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_321),
.Y(n_897)
);

BUFx5_ASAP7_75t_L g898 ( 
.A(n_491),
.Y(n_898)
);

BUFx10_ASAP7_75t_L g899 ( 
.A(n_608),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_460),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_787),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_732),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_673),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_778),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_292),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_570),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_609),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_281),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_760),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_48),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_802),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_669),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_538),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_210),
.Y(n_914)
);

BUFx10_ASAP7_75t_L g915 ( 
.A(n_109),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_369),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_656),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_620),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_794),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_305),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_1),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_676),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_578),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_453),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_574),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_20),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_67),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_313),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_614),
.Y(n_929)
);

BUFx5_ASAP7_75t_L g930 ( 
.A(n_659),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_625),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_98),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_106),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_747),
.Y(n_934)
);

BUFx10_ASAP7_75t_L g935 ( 
.A(n_45),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_660),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_793),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_316),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_636),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_703),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_498),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_257),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_463),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_758),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_247),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_648),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_406),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_315),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_279),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_759),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_53),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_643),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_105),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_769),
.Y(n_954)
);

CKINVDCx16_ASAP7_75t_R g955 ( 
.A(n_743),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_298),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_574),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_107),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_259),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_69),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_679),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_464),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_171),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_477),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_258),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_459),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_789),
.Y(n_967)
);

CKINVDCx14_ASAP7_75t_R g968 ( 
.A(n_673),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_204),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_784),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_288),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_713),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_792),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_309),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_395),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_462),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_786),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_475),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_768),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_226),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_424),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_74),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_464),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_10),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_484),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_810),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_677),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_667),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_525),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_587),
.Y(n_990)
);

CKINVDCx16_ASAP7_75t_R g991 ( 
.A(n_356),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_406),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_773),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_796),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_178),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_353),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_457),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_781),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_616),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_258),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_29),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_618),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_5),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_808),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_764),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_680),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_775),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_810),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_704),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_119),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_486),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_161),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_501),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_283),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_770),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_803),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_473),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_167),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_714),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_40),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_618),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_283),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_762),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_352),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_483),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_418),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_815),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_336),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_400),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_398),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_455),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_653),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_379),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_586),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_420),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_658),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_262),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_608),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_28),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_637),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_776),
.Y(n_1041)
);

CKINVDCx20_ASAP7_75t_R g1042 ( 
.A(n_721),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_26),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_486),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_233),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_648),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_643),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_302),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_729),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_674),
.Y(n_1050)
);

CKINVDCx14_ASAP7_75t_R g1051 ( 
.A(n_512),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_301),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_516),
.Y(n_1053)
);

CKINVDCx16_ASAP7_75t_R g1054 ( 
.A(n_354),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_804),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_758),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_10),
.Y(n_1057)
);

CKINVDCx16_ASAP7_75t_R g1058 ( 
.A(n_808),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_161),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_314),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_299),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_576),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_442),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_619),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_139),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_582),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_325),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_242),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_37),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_129),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_751),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_756),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_666),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_577),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_393),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_221),
.Y(n_1076)
);

CKINVDCx16_ASAP7_75t_R g1077 ( 
.A(n_101),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_347),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_401),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_779),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_332),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_153),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_362),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_544),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_250),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_44),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_149),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_604),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_45),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_209),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_540),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_88),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_465),
.Y(n_1093)
);

CKINVDCx14_ASAP7_75t_R g1094 ( 
.A(n_491),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_510),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_201),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_324),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_410),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_125),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_204),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_809),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_694),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_720),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_372),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_746),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_405),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_513),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_54),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_800),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_375),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_609),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_413),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_425),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_532),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_386),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_829),
.Y(n_1116)
);

CKINVDCx16_ASAP7_75t_R g1117 ( 
.A(n_224),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_405),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_694),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_436),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_318),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_97),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_777),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_732),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_178),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_268),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_205),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_345),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_131),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_280),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_262),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_76),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_692),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_780),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_223),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_374),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_457),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_782),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_676),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_251),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_756),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_117),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_241),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_795),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_693),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_563),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_521),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_91),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_97),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_122),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_270),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_824),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_88),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_739),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_411),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_444),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_626),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_182),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_527),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_517),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_427),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_265),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_81),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_32),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_477),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_269),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_584),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_371),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_781),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_549),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_208),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_811),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_166),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_693),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_783),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_765),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_549),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_340),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_801),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_6),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_590),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_809),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_598),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_699),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_223),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_589),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_741),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_503),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_461),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_783),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_140),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_658),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_814),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_785),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_672),
.Y(n_1195)
);

CKINVDCx16_ASAP7_75t_R g1196 ( 
.A(n_749),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_524),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_435),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_218),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_710),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_182),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_825),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_6),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_670),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_383),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_201),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_345),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_632),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_8),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_393),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_379),
.Y(n_1211)
);

BUFx3_ASAP7_75t_L g1212 ( 
.A(n_475),
.Y(n_1212)
);

CKINVDCx20_ASAP7_75t_R g1213 ( 
.A(n_307),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_199),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_519),
.Y(n_1215)
);

BUFx2_ASAP7_75t_SL g1216 ( 
.A(n_704),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_798),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_350),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_739),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_349),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_109),
.Y(n_1221)
);

CKINVDCx20_ASAP7_75t_R g1222 ( 
.A(n_587),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_36),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_82),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_599),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_653),
.Y(n_1226)
);

BUFx5_ASAP7_75t_L g1227 ( 
.A(n_202),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_391),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_173),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_763),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_774),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_605),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_578),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_480),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_802),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_714),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_211),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_814),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_172),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_791),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_199),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_206),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_330),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_427),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_15),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_425),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_168),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_22),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_760),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_525),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_151),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_249),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_308),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_217),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_514),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_65),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_231),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_203),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_106),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_806),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_157),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_314),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_746),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_114),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_553),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_543),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_520),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_496),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_408),
.Y(n_1269)
);

BUFx2_ASAP7_75t_SL g1270 ( 
.A(n_750),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_212),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_489),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_77),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_498),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_108),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_432),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_288),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_168),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_669),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_478),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_805),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_151),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_623),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_363),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_703),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_169),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_660),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_516),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_564),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_784),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_373),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_455),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_227),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_471),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_424),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_143),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_686),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_595),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_336),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_361),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_281),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_125),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_375),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_640),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_801),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_435),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_210),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_786),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_409),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_588),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_73),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_589),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_636),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_679),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_214),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_695),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_506),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_724),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_90),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_528),
.Y(n_1320)
);

CKINVDCx16_ASAP7_75t_R g1321 ( 
.A(n_788),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_797),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_130),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_626),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_259),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_504),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_417),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_47),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_747),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_263),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_675),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_26),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_308),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_447),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_114),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_159),
.Y(n_1336)
);

CKINVDCx14_ASAP7_75t_R g1337 ( 
.A(n_729),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_554),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_755),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_263),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_222),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_799),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_431),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_117),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_471),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_485),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_649),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_766),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_99),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_622),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_533),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_535),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_356),
.Y(n_1353)
);

BUFx2_ASAP7_75t_SL g1354 ( 
.A(n_54),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_757),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_357),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_462),
.Y(n_1357)
);

CKINVDCx16_ASAP7_75t_R g1358 ( 
.A(n_315),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_612),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_153),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_850),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_946),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_859),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_946),
.Y(n_1364)
);

BUFx8_ASAP7_75t_SL g1365 ( 
.A(n_862),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_946),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1306),
.B(n_0),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_936),
.B(n_0),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_894),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_898),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_898),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_982),
.B(n_2),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_936),
.B(n_1),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_898),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_859),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_898),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_898),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1301),
.B(n_2),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1116),
.B(n_3),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_894),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_898),
.Y(n_1381)
);

BUFx2_ASAP7_75t_L g1382 ( 
.A(n_997),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1301),
.B(n_3),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_854),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_898),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1038),
.B(n_4),
.Y(n_1386)
);

BUFx8_ASAP7_75t_SL g1387 ( 
.A(n_862),
.Y(n_1387)
);

BUFx8_ASAP7_75t_SL g1388 ( 
.A(n_876),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_854),
.B(n_4),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_930),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1172),
.B(n_5),
.Y(n_1391)
);

BUFx8_ASAP7_75t_SL g1392 ( 
.A(n_876),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1174),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_859),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_869),
.B(n_7),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1204),
.B(n_7),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_866),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1313),
.B(n_8),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_869),
.Y(n_1399)
);

INVx5_ASAP7_75t_L g1400 ( 
.A(n_894),
.Y(n_1400)
);

INVx5_ASAP7_75t_L g1401 ( 
.A(n_894),
.Y(n_1401)
);

BUFx12f_ASAP7_75t_L g1402 ( 
.A(n_866),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_930),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_968),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1051),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1094),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_866),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_890),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_964),
.B(n_11),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_976),
.B(n_9),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_930),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_954),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_914),
.B(n_9),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_955),
.B(n_11),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_L g1415 ( 
.A(n_954),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_930),
.Y(n_1416)
);

INVx5_ASAP7_75t_L g1417 ( 
.A(n_954),
.Y(n_1417)
);

INVx6_ASAP7_75t_L g1418 ( 
.A(n_886),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_930),
.Y(n_1419)
);

BUFx6f_ASAP7_75t_L g1420 ( 
.A(n_954),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_890),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_886),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_886),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_991),
.B(n_12),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_998),
.B(n_1059),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1028),
.B(n_12),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_899),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1155),
.B(n_13),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_983),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_983),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_930),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1179),
.B(n_14),
.Y(n_1432)
);

BUFx6f_ASAP7_75t_L g1433 ( 
.A(n_983),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_983),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1337),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_998),
.Y(n_1436)
);

BUFx12f_ASAP7_75t_L g1437 ( 
.A(n_899),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_930),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1059),
.B(n_13),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1227),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1070),
.B(n_14),
.Y(n_1441)
);

BUFx8_ASAP7_75t_L g1442 ( 
.A(n_1227),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1054),
.B(n_16),
.Y(n_1443)
);

INVx5_ASAP7_75t_L g1444 ( 
.A(n_1036),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1058),
.B(n_16),
.Y(n_1445)
);

NOR2x1_ASAP7_75t_L g1446 ( 
.A(n_1070),
.B(n_15),
.Y(n_1446)
);

INVx5_ASAP7_75t_L g1447 ( 
.A(n_1036),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1227),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1036),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1036),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1227),
.Y(n_1451)
);

INVx5_ASAP7_75t_L g1452 ( 
.A(n_1045),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1077),
.B(n_18),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1045),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1099),
.B(n_17),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1099),
.B(n_17),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_961),
.B(n_18),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_840),
.B(n_19),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1203),
.B(n_19),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1227),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1203),
.B(n_20),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_870),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1173),
.B(n_21),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1212),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1117),
.B(n_22),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1196),
.B(n_21),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1045),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1212),
.B(n_23),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1045),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1261),
.B(n_1286),
.Y(n_1470)
);

BUFx12f_ASAP7_75t_L g1471 ( 
.A(n_899),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1321),
.B(n_1358),
.Y(n_1472)
);

BUFx8_ASAP7_75t_L g1473 ( 
.A(n_1227),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1227),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1261),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1286),
.Y(n_1476)
);

BUFx12f_ASAP7_75t_L g1477 ( 
.A(n_915),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1317),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_915),
.B(n_935),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1317),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_870),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1121),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_SL g1483 ( 
.A(n_1329),
.B(n_838),
.Y(n_1483)
);

INVx5_ASAP7_75t_L g1484 ( 
.A(n_1121),
.Y(n_1484)
);

INVx5_ASAP7_75t_L g1485 ( 
.A(n_1121),
.Y(n_1485)
);

AND2x6_ASAP7_75t_L g1486 ( 
.A(n_1329),
.B(n_839),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_871),
.B(n_24),
.Y(n_1487)
);

BUFx8_ASAP7_75t_SL g1488 ( 
.A(n_895),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1472),
.A2(n_873),
.B1(n_874),
.B2(n_871),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1382),
.B(n_915),
.Y(n_1490)
);

AO22x2_ASAP7_75t_L g1491 ( 
.A1(n_1413),
.A2(n_1414),
.B1(n_1426),
.B2(n_1424),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1393),
.B(n_935),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1404),
.B(n_1406),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1462),
.A2(n_874),
.B1(n_875),
.B2(n_873),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1373),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1361),
.B(n_935),
.Y(n_1496)
);

AO22x2_ASAP7_75t_L g1497 ( 
.A1(n_1466),
.A2(n_864),
.B1(n_1270),
.B2(n_1216),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1481),
.A2(n_877),
.B1(n_878),
.B2(n_875),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1369),
.Y(n_1499)
);

OAI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1410),
.A2(n_878),
.B1(n_879),
.B2(n_877),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1435),
.B(n_1348),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1443),
.A2(n_882),
.B1(n_883),
.B2(n_879),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1479),
.A2(n_883),
.B1(n_887),
.B2(n_882),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1373),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_1365),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1418),
.B(n_1348),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1367),
.A2(n_888),
.B1(n_891),
.B2(n_887),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1418),
.B(n_1348),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1379),
.A2(n_891),
.B1(n_1316),
.B2(n_888),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1375),
.B(n_842),
.Y(n_1510)
);

AND2x2_ASAP7_75t_SL g1511 ( 
.A(n_1378),
.B(n_845),
.Y(n_1511)
);

OAI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1445),
.A2(n_1318),
.B1(n_1319),
.B2(n_1316),
.Y(n_1512)
);

AO22x2_ASAP7_75t_L g1513 ( 
.A1(n_1378),
.A2(n_1354),
.B1(n_900),
.B2(n_969),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1375),
.B(n_1333),
.Y(n_1514)
);

OAI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1453),
.A2(n_1319),
.B1(n_1320),
.B2(n_1318),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1383),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1386),
.A2(n_1324),
.B1(n_1326),
.B2(n_1320),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1391),
.A2(n_1326),
.B1(n_1328),
.B2(n_1324),
.Y(n_1518)
);

AO22x2_ASAP7_75t_L g1519 ( 
.A1(n_1383),
.A2(n_989),
.B1(n_1013),
.B2(n_847),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1396),
.A2(n_1331),
.B1(n_1328),
.B2(n_848),
.Y(n_1520)
);

INVxp33_ASAP7_75t_L g1521 ( 
.A(n_1387),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1394),
.B(n_1333),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1394),
.B(n_1331),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1407),
.B(n_1423),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1384),
.Y(n_1525)
);

AO22x2_ASAP7_75t_L g1526 ( 
.A1(n_1389),
.A2(n_1049),
.B1(n_1100),
.B2(n_1015),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1405),
.A2(n_849),
.B1(n_851),
.B2(n_844),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1389),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1407),
.Y(n_1529)
);

BUFx6f_ASAP7_75t_L g1530 ( 
.A(n_1369),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1395),
.Y(n_1531)
);

AO22x2_ASAP7_75t_L g1532 ( 
.A1(n_1395),
.A2(n_1277),
.B1(n_1300),
.B2(n_1246),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1423),
.B(n_1351),
.Y(n_1533)
);

OAI22xp33_ASAP7_75t_R g1534 ( 
.A1(n_1388),
.A2(n_843),
.B1(n_846),
.B2(n_841),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1427),
.B(n_1347),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1427),
.B(n_1347),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1439),
.A2(n_855),
.B1(n_856),
.B2(n_853),
.Y(n_1537)
);

AOI22x1_ASAP7_75t_L g1538 ( 
.A1(n_1371),
.A2(n_907),
.B1(n_909),
.B2(n_845),
.Y(n_1538)
);

OA22x2_ASAP7_75t_L g1539 ( 
.A1(n_1372),
.A2(n_1432),
.B1(n_1409),
.B2(n_1465),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1366),
.B(n_852),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1439),
.Y(n_1541)
);

OA22x2_ASAP7_75t_L g1542 ( 
.A1(n_1487),
.A2(n_917),
.B1(n_925),
.B2(n_896),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1408),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1421),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1363),
.B(n_1397),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1402),
.B(n_907),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1422),
.B(n_909),
.Y(n_1547)
);

OAI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1368),
.A2(n_860),
.B1(n_863),
.B2(n_857),
.Y(n_1548)
);

AO22x2_ASAP7_75t_L g1549 ( 
.A1(n_1441),
.A2(n_1359),
.B1(n_1357),
.B2(n_861),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1441),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1368),
.A2(n_865),
.B1(n_868),
.B2(n_867),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1475),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1455),
.A2(n_897),
.B1(n_901),
.B2(n_893),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1437),
.B(n_923),
.Y(n_1554)
);

AO22x2_ASAP7_75t_L g1555 ( 
.A1(n_1455),
.A2(n_1352),
.B1(n_1356),
.B2(n_1349),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1442),
.B(n_1344),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1458),
.A2(n_1355),
.B1(n_928),
.B2(n_990),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1471),
.B(n_923),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1477),
.A2(n_928),
.B1(n_990),
.B2(n_895),
.Y(n_1559)
);

AO22x2_ASAP7_75t_L g1560 ( 
.A1(n_1456),
.A2(n_872),
.B1(n_880),
.B2(n_858),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1392),
.A2(n_1000),
.B1(n_1001),
.B2(n_992),
.Y(n_1561)
);

AO22x2_ASAP7_75t_L g1562 ( 
.A1(n_1456),
.A2(n_1343),
.B1(n_1340),
.B2(n_884),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1425),
.B(n_932),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1478),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1459),
.A2(n_905),
.B1(n_911),
.B2(n_904),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1459),
.A2(n_916),
.B1(n_919),
.B2(n_913),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1458),
.A2(n_1355),
.B1(n_1000),
.B2(n_1001),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1398),
.A2(n_921),
.B1(n_922),
.B2(n_920),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1461),
.A2(n_927),
.B1(n_931),
.B2(n_924),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1399),
.B(n_1334),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1366),
.B(n_933),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1428),
.A2(n_940),
.B1(n_942),
.B2(n_938),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1461),
.A2(n_947),
.B1(n_949),
.B2(n_944),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1480),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1488),
.A2(n_1011),
.B1(n_1039),
.B2(n_992),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1362),
.B(n_932),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1442),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1399),
.Y(n_1578)
);

AO22x2_ASAP7_75t_L g1579 ( 
.A1(n_1468),
.A2(n_1425),
.B1(n_1470),
.B2(n_1364),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1436),
.B(n_950),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1436),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1468),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1364),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1470),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1464),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1362),
.B(n_999),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1362),
.A2(n_1039),
.B1(n_1042),
.B2(n_1011),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1483),
.A2(n_1065),
.B1(n_1068),
.B2(n_1042),
.Y(n_1588)
);

OA22x2_ASAP7_75t_L g1589 ( 
.A1(n_1464),
.A2(n_979),
.B1(n_993),
.B2(n_970),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1370),
.A2(n_956),
.B1(n_959),
.B2(n_951),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_SL g1591 ( 
.A1(n_1457),
.A2(n_962),
.B1(n_963),
.B2(n_960),
.Y(n_1591)
);

AOI22x1_ASAP7_75t_L g1592 ( 
.A1(n_1374),
.A2(n_1008),
.B1(n_1023),
.B2(n_999),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1473),
.A2(n_966),
.B1(n_972),
.B2(n_965),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1463),
.A2(n_1068),
.B1(n_1069),
.B2(n_1065),
.Y(n_1594)
);

AO22x2_ASAP7_75t_L g1595 ( 
.A1(n_1476),
.A2(n_885),
.B1(n_889),
.B2(n_881),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1370),
.A2(n_978),
.B1(n_980),
.B2(n_975),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1446),
.A2(n_1071),
.B1(n_1092),
.B2(n_1069),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1476),
.B(n_981),
.Y(n_1598)
);

OAI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1483),
.A2(n_1092),
.B1(n_1102),
.B2(n_1071),
.Y(n_1599)
);

CKINVDCx16_ASAP7_75t_R g1600 ( 
.A(n_1486),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1473),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1381),
.B(n_1008),
.Y(n_1602)
);

OA22x2_ASAP7_75t_L g1603 ( 
.A1(n_1381),
.A2(n_1010),
.B1(n_1030),
.B2(n_996),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1446),
.B(n_1023),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1385),
.B(n_1474),
.Y(n_1605)
);

NAND3x1_ASAP7_75t_L g1606 ( 
.A(n_1385),
.B(n_1113),
.C(n_1102),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1438),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1438),
.A2(n_1118),
.B1(n_1119),
.B2(n_1113),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1460),
.B(n_1327),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1460),
.B(n_1336),
.Y(n_1610)
);

NAND3x1_ASAP7_75t_L g1611 ( 
.A(n_1474),
.B(n_1119),
.C(n_1118),
.Y(n_1611)
);

AO22x2_ASAP7_75t_L g1612 ( 
.A1(n_1376),
.A2(n_1332),
.B1(n_1330),
.B2(n_902),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1377),
.B(n_1027),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1390),
.B(n_1338),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1403),
.A2(n_1185),
.B1(n_1192),
.B2(n_1163),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1486),
.A2(n_986),
.B1(n_987),
.B2(n_985),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1400),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1486),
.A2(n_1002),
.B1(n_1003),
.B2(n_994),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1486),
.A2(n_1005),
.B1(n_1006),
.B2(n_1004),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1411),
.A2(n_1185),
.B1(n_1192),
.B2(n_1163),
.Y(n_1620)
);

AND2x2_ASAP7_75t_SL g1621 ( 
.A(n_1416),
.B(n_1027),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1419),
.B(n_1339),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1400),
.Y(n_1623)
);

NOR2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1431),
.B(n_903),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1440),
.A2(n_1213),
.B1(n_1222),
.B2(n_1197),
.Y(n_1625)
);

OAI22xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1448),
.A2(n_1012),
.B1(n_1014),
.B2(n_1009),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1451),
.A2(n_1213),
.B1(n_1222),
.B2(n_1197),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1400),
.A2(n_1020),
.B1(n_1026),
.B2(n_1018),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1401),
.A2(n_1034),
.B1(n_1037),
.B2(n_1033),
.Y(n_1629)
);

AOI22xp5_ASAP7_75t_L g1630 ( 
.A1(n_1401),
.A2(n_1043),
.B1(n_1044),
.B2(n_1041),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1401),
.B(n_1327),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_SL g1632 ( 
.A(n_1369),
.Y(n_1632)
);

NAND3x1_ASAP7_75t_L g1633 ( 
.A(n_1417),
.B(n_1263),
.C(n_1252),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1417),
.B(n_1335),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1417),
.B(n_1335),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1380),
.Y(n_1636)
);

AO22x2_ASAP7_75t_L g1637 ( 
.A1(n_1444),
.A2(n_1325),
.B1(n_906),
.B2(n_908),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1444),
.A2(n_1047),
.B1(n_1048),
.B2(n_1046),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1485),
.B(n_1063),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1444),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1447),
.B(n_1050),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1447),
.B(n_1063),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1447),
.A2(n_1263),
.B1(n_1252),
.B2(n_910),
.Y(n_1643)
);

OAI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1449),
.A2(n_912),
.B1(n_918),
.B2(n_892),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1485),
.B(n_1323),
.Y(n_1645)
);

OAI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1449),
.A2(n_929),
.B1(n_934),
.B2(n_926),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1449),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1452),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1452),
.B(n_1082),
.Y(n_1649)
);

AOI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1452),
.A2(n_1053),
.B1(n_1055),
.B2(n_1052),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1469),
.B(n_1484),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1469),
.A2(n_1060),
.B1(n_1061),
.B2(n_1056),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1469),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1484),
.B(n_1082),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1484),
.B(n_1064),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1485),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1380),
.Y(n_1657)
);

OAI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1380),
.A2(n_939),
.B1(n_941),
.B2(n_937),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1412),
.A2(n_1073),
.B1(n_1075),
.B2(n_1066),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1412),
.Y(n_1660)
);

OAI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1412),
.A2(n_1079),
.B1(n_1080),
.B2(n_1078),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1415),
.B(n_943),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1415),
.B(n_945),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1415),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1420),
.B(n_1146),
.Y(n_1665)
);

OAI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1420),
.A2(n_952),
.B1(n_953),
.B2(n_948),
.Y(n_1666)
);

AOI22xp5_ASAP7_75t_L g1667 ( 
.A1(n_1420),
.A2(n_1083),
.B1(n_1084),
.B2(n_1081),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1429),
.B(n_1310),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1429),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1429),
.B(n_1085),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1430),
.B(n_1323),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1430),
.B(n_1433),
.Y(n_1672)
);

AOI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1430),
.A2(n_1089),
.B1(n_1090),
.B2(n_1086),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1433),
.B(n_957),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1433),
.Y(n_1675)
);

OAI22xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1434),
.A2(n_1095),
.B1(n_1096),
.B2(n_1093),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1434),
.A2(n_1101),
.B1(n_1104),
.B2(n_1098),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1434),
.B(n_1146),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1450),
.B(n_1105),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1450),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1450),
.Y(n_1681)
);

AO22x2_ASAP7_75t_L g1682 ( 
.A1(n_1454),
.A2(n_1315),
.B1(n_1322),
.B2(n_1311),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1454),
.B(n_1176),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1454),
.Y(n_1684)
);

OAI22xp33_ASAP7_75t_SL g1685 ( 
.A1(n_1467),
.A2(n_1108),
.B1(n_1109),
.B2(n_1106),
.Y(n_1685)
);

AO22x2_ASAP7_75t_L g1686 ( 
.A1(n_1467),
.A2(n_967),
.B1(n_971),
.B2(n_958),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1467),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1482),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1482),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1482),
.B(n_1176),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1404),
.B(n_1111),
.Y(n_1691)
);

AO22x2_ASAP7_75t_L g1692 ( 
.A1(n_1413),
.A2(n_974),
.B1(n_977),
.B2(n_973),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1382),
.A2(n_1120),
.B1(n_1122),
.B2(n_1115),
.Y(n_1693)
);

OAI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1466),
.A2(n_1124),
.B1(n_1125),
.B2(n_1123),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1384),
.Y(n_1695)
);

AO22x2_ASAP7_75t_L g1696 ( 
.A1(n_1413),
.A2(n_988),
.B1(n_995),
.B2(n_984),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1462),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1382),
.A2(n_1129),
.B1(n_1130),
.B2(n_1127),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1382),
.A2(n_1135),
.B1(n_1136),
.B2(n_1132),
.Y(n_1699)
);

OA22x2_ASAP7_75t_L g1700 ( 
.A1(n_1361),
.A2(n_1162),
.B1(n_1171),
.B2(n_1144),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1373),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1382),
.B(n_1137),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1472),
.A2(n_1140),
.B1(n_1141),
.B2(n_1139),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1529),
.B(n_1142),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1584),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1601),
.B(n_1007),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1514),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1522),
.Y(n_1708)
);

XNOR2x2_ASAP7_75t_L g1709 ( 
.A(n_1519),
.B(n_1016),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_SL g1710 ( 
.A(n_1616),
.B(n_1618),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1697),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1535),
.Y(n_1712)
);

OR2x6_ASAP7_75t_L g1713 ( 
.A(n_1633),
.B(n_1019),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1536),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1523),
.B(n_1145),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1505),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1612),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1524),
.B(n_1147),
.Y(n_1718)
);

OAI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1607),
.A2(n_1021),
.B(n_1017),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1702),
.Y(n_1720)
);

NAND2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1545),
.B(n_1022),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1612),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1510),
.B(n_1149),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1563),
.Y(n_1724)
);

CKINVDCx16_ASAP7_75t_R g1725 ( 
.A(n_1577),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1662),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1493),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1663),
.Y(n_1728)
);

XOR2xp5_ASAP7_75t_L g1729 ( 
.A(n_1561),
.B(n_1360),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1674),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1575),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1619),
.B(n_1121),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1496),
.B(n_1151),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1631),
.Y(n_1734)
);

BUFx5_ASAP7_75t_L g1735 ( 
.A(n_1605),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1634),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1495),
.A2(n_1025),
.B(n_1024),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1635),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1639),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1642),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1645),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1490),
.B(n_1492),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1649),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1552),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1654),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1579),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1579),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1501),
.B(n_1157),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1576),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1586),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1613),
.Y(n_1751)
);

AOI21x1_ASAP7_75t_L g1752 ( 
.A1(n_1583),
.A2(n_1031),
.B(n_1029),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1564),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1504),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1494),
.B(n_1158),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1516),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1701),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1574),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1602),
.Y(n_1759)
);

XOR2x2_ASAP7_75t_L g1760 ( 
.A(n_1625),
.B(n_23),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1559),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1498),
.B(n_1160),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1506),
.B(n_1161),
.Y(n_1763)
);

CKINVDCx16_ASAP7_75t_R g1764 ( 
.A(n_1608),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1683),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1609),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1508),
.B(n_1165),
.Y(n_1767)
);

XNOR2xp5_ASAP7_75t_L g1768 ( 
.A(n_1606),
.B(n_1167),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1540),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1533),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1682),
.Y(n_1771)
);

XOR2xp5_ASAP7_75t_L g1772 ( 
.A(n_1521),
.B(n_1346),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1682),
.Y(n_1773)
);

XNOR2x2_ASAP7_75t_L g1774 ( 
.A(n_1519),
.B(n_1032),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1686),
.Y(n_1775)
);

XNOR2xp5_ASAP7_75t_L g1776 ( 
.A(n_1611),
.B(n_1168),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1665),
.Y(n_1777)
);

XNOR2x2_ASAP7_75t_L g1778 ( 
.A(n_1526),
.B(n_1532),
.Y(n_1778)
);

CKINVDCx20_ASAP7_75t_R g1779 ( 
.A(n_1594),
.Y(n_1779)
);

XOR2xp5_ASAP7_75t_L g1780 ( 
.A(n_1491),
.B(n_1169),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1686),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1528),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1531),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1541),
.Y(n_1784)
);

BUFx5_ASAP7_75t_L g1785 ( 
.A(n_1648),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1546),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1550),
.Y(n_1787)
);

XOR2xp5_ASAP7_75t_L g1788 ( 
.A(n_1491),
.B(n_1299),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1513),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1582),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1668),
.Y(n_1791)
);

CKINVDCx5p33_ASAP7_75t_R g1792 ( 
.A(n_1703),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1671),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1597),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1691),
.B(n_1170),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1507),
.B(n_1175),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1557),
.B(n_1305),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1571),
.B(n_1177),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1610),
.A2(n_1040),
.B(n_1035),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1678),
.Y(n_1800)
);

CKINVDCx20_ASAP7_75t_R g1801 ( 
.A(n_1693),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1690),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1509),
.B(n_1178),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1549),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1549),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1511),
.B(n_1180),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1555),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1555),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1560),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1517),
.B(n_1181),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1560),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1562),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1657),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1570),
.B(n_1580),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1518),
.B(n_1183),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1698),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1562),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1503),
.B(n_1520),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1624),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1595),
.Y(n_1820)
);

BUFx2_ASAP7_75t_L g1821 ( 
.A(n_1513),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1567),
.B(n_1615),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1525),
.Y(n_1823)
);

XOR2xp5_ASAP7_75t_L g1824 ( 
.A(n_1587),
.B(n_1342),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1595),
.Y(n_1825)
);

XOR2xp5_ASAP7_75t_L g1826 ( 
.A(n_1588),
.B(n_1599),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1620),
.B(n_1345),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1543),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1544),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1695),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1699),
.B(n_1184),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1497),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1497),
.Y(n_1833)
);

INVx4_ASAP7_75t_SL g1834 ( 
.A(n_1632),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1547),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1538),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1692),
.B(n_1696),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1592),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1614),
.A2(n_1062),
.B(n_1057),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1578),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1539),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1621),
.Y(n_1842)
);

INVxp67_ASAP7_75t_SL g1843 ( 
.A(n_1500),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1627),
.B(n_1295),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1692),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1696),
.B(n_1186),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1600),
.B(n_1128),
.Y(n_1847)
);

NOR3xp33_ASAP7_75t_L g1848 ( 
.A(n_1643),
.B(n_1189),
.C(n_1188),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1581),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1585),
.Y(n_1850)
);

NAND2xp33_ASAP7_75t_SL g1851 ( 
.A(n_1556),
.B(n_1307),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1554),
.B(n_1190),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1603),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1558),
.B(n_1191),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1617),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1637),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1637),
.Y(n_1857)
);

OR2x6_ASAP7_75t_L g1858 ( 
.A(n_1526),
.B(n_1304),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1604),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1573),
.B(n_1128),
.Y(n_1860)
);

CKINVDCx20_ASAP7_75t_R g1861 ( 
.A(n_1593),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1604),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1527),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1589),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1670),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1679),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1658),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1598),
.B(n_1193),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1666),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1542),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1537),
.B(n_1194),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1622),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1644),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1489),
.B(n_1312),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1646),
.Y(n_1875)
);

BUFx3_ASAP7_75t_L g1876 ( 
.A(n_1623),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1661),
.Y(n_1877)
);

OR2x2_ASAP7_75t_L g1878 ( 
.A(n_1502),
.B(n_1314),
.Y(n_1878)
);

XNOR2x2_ASAP7_75t_L g1879 ( 
.A(n_1532),
.B(n_1067),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1676),
.Y(n_1880)
);

NOR2xp67_ASAP7_75t_L g1881 ( 
.A(n_1659),
.B(n_25),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1685),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1590),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1640),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1700),
.Y(n_1885)
);

NOR2xp67_ASAP7_75t_L g1886 ( 
.A(n_1667),
.B(n_25),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1553),
.B(n_1072),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1641),
.A2(n_1076),
.B(n_1074),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1565),
.B(n_1195),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1655),
.Y(n_1890)
);

XOR2x2_ASAP7_75t_L g1891 ( 
.A(n_1512),
.B(n_24),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1596),
.A2(n_1088),
.B(n_1087),
.Y(n_1892)
);

INVxp33_ASAP7_75t_L g1893 ( 
.A(n_1673),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1677),
.A2(n_1097),
.B(n_1091),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1647),
.Y(n_1895)
);

XOR2xp5_ASAP7_75t_L g1896 ( 
.A(n_1566),
.B(n_1298),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1569),
.B(n_1628),
.Y(n_1897)
);

NOR2xp67_ASAP7_75t_L g1898 ( 
.A(n_1629),
.B(n_28),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1653),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1656),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1626),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1548),
.Y(n_1902)
);

BUFx6f_ASAP7_75t_L g1903 ( 
.A(n_1651),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1551),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1591),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1687),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1499),
.Y(n_1907)
);

CKINVDCx20_ASAP7_75t_R g1908 ( 
.A(n_1630),
.Y(n_1908)
);

INVxp67_ASAP7_75t_L g1909 ( 
.A(n_1638),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1694),
.Y(n_1910)
);

XOR2x2_ASAP7_75t_L g1911 ( 
.A(n_1568),
.B(n_27),
.Y(n_1911)
);

XNOR2xp5_ASAP7_75t_L g1912 ( 
.A(n_1515),
.B(n_1199),
.Y(n_1912)
);

INVxp67_ASAP7_75t_SL g1913 ( 
.A(n_1650),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1572),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1652),
.Y(n_1915)
);

HB1xp67_ASAP7_75t_L g1916 ( 
.A(n_1534),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1636),
.B(n_1200),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1672),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1664),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1684),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1689),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1660),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1669),
.A2(n_1680),
.B(n_1675),
.Y(n_1923)
);

XNOR2xp5_ASAP7_75t_L g1924 ( 
.A(n_1681),
.B(n_1202),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1499),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1530),
.B(n_1205),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_L g1927 ( 
.A(n_1530),
.B(n_29),
.Y(n_1927)
);

XOR2xp5_ASAP7_75t_L g1928 ( 
.A(n_1688),
.B(n_1353),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1688),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1529),
.B(n_1206),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1584),
.Y(n_1931)
);

XNOR2x2_ASAP7_75t_L g1932 ( 
.A(n_1519),
.B(n_1103),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1584),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1662),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1584),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1584),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1584),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1584),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1616),
.B(n_1128),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1529),
.B(n_1207),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1584),
.Y(n_1941)
);

NAND2x1p5_ASAP7_75t_L g1942 ( 
.A(n_1601),
.B(n_1107),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1584),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1584),
.Y(n_1944)
);

AND2x6_ASAP7_75t_L g1945 ( 
.A(n_1600),
.B(n_1292),
.Y(n_1945)
);

AOI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1495),
.A2(n_1112),
.B(n_1110),
.Y(n_1946)
);

BUFx5_ASAP7_75t_L g1947 ( 
.A(n_1605),
.Y(n_1947)
);

AND2x2_ASAP7_75t_SL g1948 ( 
.A(n_1545),
.B(n_1302),
.Y(n_1948)
);

BUFx6f_ASAP7_75t_L g1949 ( 
.A(n_1683),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1584),
.Y(n_1950)
);

INVxp33_ASAP7_75t_SL g1951 ( 
.A(n_1545),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1584),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1584),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1584),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1702),
.B(n_1208),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1702),
.B(n_1210),
.Y(n_1956)
);

INVx4_ASAP7_75t_SL g1957 ( 
.A(n_1601),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1662),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1584),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1584),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1584),
.Y(n_1961)
);

INVx1_ASAP7_75t_SL g1962 ( 
.A(n_1702),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1584),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1514),
.B(n_1211),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1662),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1584),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1584),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1529),
.B(n_1214),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1584),
.Y(n_1969)
);

CKINVDCx20_ASAP7_75t_R g1970 ( 
.A(n_1577),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1662),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1702),
.B(n_1218),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1529),
.B(n_1219),
.Y(n_1973)
);

INVx4_ASAP7_75t_SL g1974 ( 
.A(n_1601),
.Y(n_1974)
);

NOR2xp67_ASAP7_75t_L g1975 ( 
.A(n_1545),
.B(n_30),
.Y(n_1975)
);

NAND2x1p5_ASAP7_75t_L g1976 ( 
.A(n_1601),
.B(n_1114),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1584),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_1577),
.Y(n_1978)
);

BUFx5_ASAP7_75t_L g1979 ( 
.A(n_1605),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1584),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1584),
.Y(n_1981)
);

INVxp33_ASAP7_75t_L g1982 ( 
.A(n_1625),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1702),
.B(n_1220),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1584),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1584),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1529),
.B(n_1221),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1529),
.B(n_1224),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1584),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1584),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1514),
.B(n_1228),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1584),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1662),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1702),
.B(n_1229),
.Y(n_1993)
);

CKINVDCx20_ASAP7_75t_R g1994 ( 
.A(n_1577),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1584),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1770),
.B(n_1230),
.Y(n_1996)
);

INVxp67_ASAP7_75t_SL g1997 ( 
.A(n_1771),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1947),
.Y(n_1998)
);

HB1xp67_ASAP7_75t_L g1999 ( 
.A(n_1727),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1947),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1957),
.B(n_1126),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1947),
.Y(n_2002)
);

OAI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1836),
.A2(n_1133),
.B(n_1131),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1947),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1962),
.B(n_1231),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1947),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1970),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1720),
.B(n_1232),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1979),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1742),
.B(n_1909),
.Y(n_2010)
);

CKINVDCx6p67_ASAP7_75t_R g2011 ( 
.A(n_1725),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1979),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_1979),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1979),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1979),
.B(n_1233),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1711),
.B(n_1234),
.Y(n_2016)
);

BUFx12f_ASAP7_75t_L g2017 ( 
.A(n_1716),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1769),
.B(n_1236),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1846),
.B(n_1237),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1735),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1955),
.B(n_1239),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1735),
.B(n_1243),
.Y(n_2022)
);

AND2x2_ASAP7_75t_SL g2023 ( 
.A(n_1764),
.B(n_1134),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1735),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1956),
.B(n_1244),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1735),
.B(n_1245),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1915),
.B(n_1248),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1872),
.B(n_1249),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1972),
.B(n_1250),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1907),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1706),
.B(n_1251),
.Y(n_2031)
);

OR2x2_ASAP7_75t_SL g2032 ( 
.A(n_1916),
.B(n_1138),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_1706),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1983),
.B(n_1253),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1707),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1744),
.Y(n_2036)
);

AND2x4_ASAP7_75t_L g2037 ( 
.A(n_1957),
.B(n_1148),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1993),
.B(n_1733),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1708),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1835),
.B(n_1254),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1712),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1753),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1773),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1837),
.B(n_1255),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1714),
.Y(n_2045)
);

AND2x4_ASAP7_75t_SL g2046 ( 
.A(n_1978),
.B(n_1152),
.Y(n_2046)
);

INVx2_ASAP7_75t_SL g2047 ( 
.A(n_1942),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1754),
.B(n_1756),
.Y(n_2048)
);

INVxp67_ASAP7_75t_L g2049 ( 
.A(n_1928),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1730),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1828),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1757),
.B(n_1258),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1841),
.B(n_1259),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1796),
.B(n_1260),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1782),
.B(n_1262),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1934),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1783),
.B(n_1265),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1855),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1784),
.B(n_1267),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1994),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1884),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1758),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1813),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1958),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1803),
.B(n_1268),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1810),
.B(n_1271),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1787),
.B(n_1272),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1840),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1815),
.B(n_1273),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1965),
.Y(n_2070)
);

BUFx5_ASAP7_75t_L g2071 ( 
.A(n_1945),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1790),
.B(n_1274),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1797),
.B(n_1275),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1799),
.B(n_1276),
.Y(n_2074)
);

AND2x4_ASAP7_75t_L g2075 ( 
.A(n_1974),
.B(n_1853),
.Y(n_2075)
);

INVxp33_ASAP7_75t_L g2076 ( 
.A(n_1824),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1849),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1971),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_1976),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1822),
.B(n_1278),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1850),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1748),
.B(n_1279),
.Y(n_2082)
);

HB1xp67_ASAP7_75t_L g2083 ( 
.A(n_1775),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1873),
.B(n_1281),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1875),
.B(n_1867),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1895),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_1974),
.B(n_1153),
.Y(n_2087)
);

OAI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_1838),
.A2(n_1752),
.B(n_1737),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_1883),
.B(n_1284),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1899),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1827),
.B(n_1282),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_1844),
.B(n_1287),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1992),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1900),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1786),
.B(n_1291),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1705),
.Y(n_2096)
);

INVx2_ASAP7_75t_SL g2097 ( 
.A(n_1721),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1785),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1785),
.Y(n_2099)
);

NAND2x1p5_ASAP7_75t_L g2100 ( 
.A(n_1746),
.B(n_1747),
.Y(n_2100)
);

INVx2_ASAP7_75t_SL g2101 ( 
.A(n_1917),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1931),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1813),
.Y(n_2103)
);

BUFx4f_ASAP7_75t_L g2104 ( 
.A(n_1945),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1755),
.B(n_1293),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1933),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1907),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_1859),
.B(n_1294),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_1813),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_1781),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1935),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1762),
.B(n_1296),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1831),
.B(n_1308),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_1818),
.B(n_1309),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1869),
.B(n_1341),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1936),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1856),
.B(n_1350),
.Y(n_2117)
);

BUFx3_ASAP7_75t_L g2118 ( 
.A(n_1876),
.Y(n_2118)
);

AND2x4_ASAP7_75t_L g2119 ( 
.A(n_1870),
.B(n_1154),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1946),
.B(n_1156),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1785),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1785),
.Y(n_2122)
);

AND2x2_ASAP7_75t_SL g2123 ( 
.A(n_1821),
.B(n_1159),
.Y(n_2123)
);

INVx1_ASAP7_75t_SL g2124 ( 
.A(n_1717),
.Y(n_2124)
);

NOR2xp67_ASAP7_75t_R g2125 ( 
.A(n_1857),
.B(n_1164),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1871),
.B(n_1166),
.Y(n_2126)
);

OAI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1839),
.A2(n_1187),
.B(n_1182),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_1713),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1918),
.Y(n_2129)
);

BUFx3_ASAP7_75t_L g2130 ( 
.A(n_1903),
.Y(n_2130)
);

HB1xp67_ASAP7_75t_L g2131 ( 
.A(n_1858),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_SL g2132 ( 
.A(n_1722),
.B(n_1128),
.Y(n_2132)
);

BUFx2_ASAP7_75t_SL g2133 ( 
.A(n_1945),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1903),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1814),
.B(n_1143),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1937),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_1858),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1719),
.B(n_1198),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_1845),
.B(n_1201),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1938),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1710),
.B(n_1215),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1834),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1941),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1864),
.B(n_1217),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_1804),
.B(n_1223),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1791),
.B(n_1225),
.Y(n_2146)
);

INVx1_ASAP7_75t_SL g2147 ( 
.A(n_1945),
.Y(n_2147)
);

HB1xp67_ASAP7_75t_L g2148 ( 
.A(n_1834),
.Y(n_2148)
);

BUFx8_ASAP7_75t_SL g2149 ( 
.A(n_1713),
.Y(n_2149)
);

BUFx3_ASAP7_75t_L g2150 ( 
.A(n_1903),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1943),
.Y(n_2151)
);

BUFx6f_ASAP7_75t_L g2152 ( 
.A(n_1907),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_1862),
.B(n_1269),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1944),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1829),
.Y(n_2155)
);

BUFx6f_ASAP7_75t_L g2156 ( 
.A(n_1765),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1950),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1952),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1889),
.B(n_1226),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1830),
.Y(n_2160)
);

NOR2xp33_ASAP7_75t_L g2161 ( 
.A(n_1913),
.B(n_1283),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_1823),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_1765),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1843),
.B(n_1235),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_1948),
.B(n_1238),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1777),
.Y(n_2166)
);

OAI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_1892),
.A2(n_1888),
.B(n_1732),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1759),
.B(n_1240),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1893),
.B(n_1303),
.Y(n_2169)
);

INVxp67_ASAP7_75t_SL g2170 ( 
.A(n_1726),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1953),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1766),
.B(n_1241),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_1852),
.B(n_1242),
.Y(n_2173)
);

INVx1_ASAP7_75t_SL g2174 ( 
.A(n_1789),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1854),
.B(n_1247),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_1912),
.B(n_1256),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1765),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_1778),
.Y(n_2178)
);

HB1xp67_ASAP7_75t_L g2179 ( 
.A(n_1728),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1823),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1949),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1887),
.B(n_1264),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1887),
.B(n_1266),
.Y(n_2183)
);

INVxp67_ASAP7_75t_SL g2184 ( 
.A(n_1826),
.Y(n_2184)
);

OAI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_1939),
.A2(n_1894),
.B(n_1890),
.Y(n_2185)
);

BUFx2_ASAP7_75t_L g2186 ( 
.A(n_1709),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1949),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1995),
.B(n_1280),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1806),
.B(n_1285),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1949),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_1951),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_1878),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1954),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1991),
.B(n_1288),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_1874),
.B(n_1289),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1959),
.B(n_1143),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1960),
.B(n_1143),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1961),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1963),
.B(n_1143),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_1982),
.B(n_1848),
.Y(n_2200)
);

AND2x2_ASAP7_75t_SL g2201 ( 
.A(n_1897),
.B(n_1150),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1966),
.Y(n_2202)
);

AND2x4_ASAP7_75t_L g2203 ( 
.A(n_1805),
.B(n_1807),
.Y(n_2203)
);

NOR2xp67_ASAP7_75t_R g2204 ( 
.A(n_1820),
.B(n_1825),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_1763),
.B(n_1150),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1767),
.B(n_1150),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1808),
.B(n_1150),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1967),
.B(n_1209),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_SL g2209 ( 
.A(n_1809),
.B(n_1209),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1897),
.B(n_1209),
.Y(n_2210)
);

AND2x6_ASAP7_75t_L g2211 ( 
.A(n_1811),
.B(n_1209),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_1924),
.Y(n_2212)
);

INVxp67_ASAP7_75t_L g2213 ( 
.A(n_1964),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_1774),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1793),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1969),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_1780),
.B(n_1257),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1812),
.B(n_1257),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1800),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1802),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_1788),
.B(n_1257),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_1718),
.B(n_1257),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1977),
.B(n_1290),
.Y(n_2223)
);

NOR2xp33_ASAP7_75t_L g2224 ( 
.A(n_1795),
.B(n_1290),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1817),
.B(n_1290),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1980),
.B(n_1290),
.Y(n_2226)
);

BUFx2_ASAP7_75t_L g2227 ( 
.A(n_1932),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_1879),
.Y(n_2228)
);

AND2x2_ASAP7_75t_SL g2229 ( 
.A(n_1832),
.B(n_1297),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1734),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1981),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_1736),
.Y(n_2232)
);

BUFx3_ASAP7_75t_L g2233 ( 
.A(n_1877),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_SL g2234 ( 
.A(n_1901),
.B(n_1905),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_1990),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1984),
.B(n_1297),
.Y(n_2236)
);

AND2x2_ASAP7_75t_SL g2237 ( 
.A(n_1833),
.B(n_1297),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_1985),
.B(n_1297),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1988),
.Y(n_2239)
);

BUFx2_ASAP7_75t_L g2240 ( 
.A(n_1863),
.Y(n_2240)
);

INVxp33_ASAP7_75t_L g2241 ( 
.A(n_1896),
.Y(n_2241)
);

NOR2xp67_ASAP7_75t_R g2242 ( 
.A(n_1902),
.B(n_27),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1738),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_1751),
.B(n_837),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1989),
.Y(n_2245)
);

AND2x6_ASAP7_75t_L g2246 ( 
.A(n_1880),
.B(n_30),
.Y(n_2246)
);

INVx3_ASAP7_75t_L g2247 ( 
.A(n_1739),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_1740),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1904),
.B(n_31),
.Y(n_2249)
);

AND2x4_ASAP7_75t_L g2250 ( 
.A(n_1910),
.B(n_31),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1749),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_1816),
.B(n_1914),
.Y(n_2252)
);

INVx1_ASAP7_75t_SL g2253 ( 
.A(n_1882),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_1881),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1704),
.B(n_823),
.Y(n_2255)
);

OAI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_1865),
.A2(n_32),
.B(n_33),
.Y(n_2256)
);

OAI21xp5_ASAP7_75t_L g2257 ( 
.A1(n_1866),
.A2(n_33),
.B(n_34),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_1930),
.B(n_1940),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1842),
.B(n_825),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1741),
.Y(n_2260)
);

INVxp67_ASAP7_75t_SL g2261 ( 
.A(n_1886),
.Y(n_2261)
);

NAND2x1p5_ASAP7_75t_L g2262 ( 
.A(n_1847),
.B(n_34),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1743),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1968),
.B(n_827),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_1745),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_1750),
.B(n_827),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1724),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_1792),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_1715),
.B(n_35),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_1819),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1723),
.B(n_828),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1860),
.Y(n_2272)
);

BUFx3_ASAP7_75t_L g2273 ( 
.A(n_1885),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1975),
.B(n_1898),
.Y(n_2274)
);

AND2x2_ASAP7_75t_SL g2275 ( 
.A(n_1760),
.B(n_35),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1919),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1798),
.B(n_829),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1973),
.B(n_830),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_1986),
.B(n_1987),
.Y(n_2279)
);

INVx4_ASAP7_75t_L g2280 ( 
.A(n_1891),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1768),
.B(n_830),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1926),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_1776),
.B(n_831),
.Y(n_2283)
);

INVx3_ASAP7_75t_L g2284 ( 
.A(n_1906),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1920),
.Y(n_2285)
);

HB1xp67_ASAP7_75t_L g2286 ( 
.A(n_1729),
.Y(n_2286)
);

NAND2x1p5_ASAP7_75t_L g2287 ( 
.A(n_1927),
.B(n_36),
.Y(n_2287)
);

OAI21xp5_ASAP7_75t_L g2288 ( 
.A1(n_1923),
.A2(n_37),
.B(n_38),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_1801),
.B(n_1911),
.Y(n_2289)
);

BUFx3_ASAP7_75t_L g2290 ( 
.A(n_1772),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_1908),
.B(n_1861),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1921),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_1868),
.B(n_833),
.Y(n_2293)
);

OAI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_1922),
.A2(n_38),
.B(n_39),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_1925),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_1779),
.Y(n_2296)
);

AND2x6_ASAP7_75t_L g2297 ( 
.A(n_1929),
.B(n_39),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1851),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_1794),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1761),
.Y(n_2300)
);

INVx3_ASAP7_75t_SL g2301 ( 
.A(n_1731),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1770),
.B(n_835),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_1907),
.Y(n_2303)
);

BUFx3_ASAP7_75t_L g2304 ( 
.A(n_1970),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1947),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1947),
.Y(n_2306)
);

OAI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_1836),
.A2(n_40),
.B(n_41),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_1947),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_1770),
.B(n_836),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1947),
.B(n_836),
.Y(n_2310)
);

INVx3_ASAP7_75t_L g2311 ( 
.A(n_1947),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_1770),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1947),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_1947),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_1942),
.Y(n_2315)
);

OAI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_1836),
.A2(n_41),
.B(n_42),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_1947),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_1770),
.B(n_42),
.Y(n_2318)
);

INVx4_ASAP7_75t_L g2319 ( 
.A(n_1834),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1947),
.Y(n_2320)
);

BUFx3_ASAP7_75t_L g2321 ( 
.A(n_1970),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1947),
.B(n_818),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1947),
.B(n_818),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_L g2324 ( 
.A(n_1770),
.B(n_43),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_1947),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1947),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_1770),
.B(n_819),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_1770),
.B(n_819),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_1770),
.B(n_43),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1947),
.Y(n_2330)
);

INVx1_ASAP7_75t_SL g2331 ( 
.A(n_1727),
.Y(n_2331)
);

OAI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_1836),
.A2(n_44),
.B(n_46),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_1770),
.B(n_822),
.Y(n_2333)
);

INVx3_ASAP7_75t_SL g2334 ( 
.A(n_1834),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1947),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1947),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_1947),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1770),
.B(n_822),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2331),
.B(n_46),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_2311),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2047),
.B(n_47),
.Y(n_2341)
);

NOR2xp67_ASAP7_75t_L g2342 ( 
.A(n_2319),
.B(n_48),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2129),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2077),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_2030),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2048),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2048),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2030),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2081),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2315),
.B(n_49),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_1999),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2170),
.B(n_49),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2331),
.B(n_50),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_1999),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2068),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2114),
.B(n_50),
.Y(n_2356)
);

INVx2_ASAP7_75t_L g2357 ( 
.A(n_2062),
.Y(n_2357)
);

BUFx4f_ASAP7_75t_L g2358 ( 
.A(n_2011),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2192),
.B(n_51),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2312),
.B(n_51),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2170),
.B(n_52),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2155),
.Y(n_2362)
);

BUFx2_ASAP7_75t_SL g2363 ( 
.A(n_2071),
.Y(n_2363)
);

AND2x4_ASAP7_75t_L g2364 ( 
.A(n_2079),
.B(n_52),
.Y(n_2364)
);

BUFx6f_ASAP7_75t_L g2365 ( 
.A(n_2030),
.Y(n_2365)
);

CKINVDCx8_ASAP7_75t_R g2366 ( 
.A(n_2133),
.Y(n_2366)
);

OR2x6_ASAP7_75t_L g2367 ( 
.A(n_2017),
.B(n_53),
.Y(n_2367)
);

BUFx2_ASAP7_75t_L g2368 ( 
.A(n_2312),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2179),
.B(n_55),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2160),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2096),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2179),
.B(n_55),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_2149),
.Y(n_2373)
);

OR2x6_ASAP7_75t_L g2374 ( 
.A(n_2079),
.B(n_56),
.Y(n_2374)
);

AND2x2_ASAP7_75t_L g2375 ( 
.A(n_2192),
.B(n_56),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2091),
.B(n_57),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2080),
.B(n_57),
.Y(n_2377)
);

INVxp67_ASAP7_75t_SL g2378 ( 
.A(n_2006),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2102),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2195),
.B(n_2235),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2276),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2235),
.B(n_2050),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2191),
.B(n_58),
.Y(n_2383)
);

NAND2x1p5_ASAP7_75t_L g2384 ( 
.A(n_2319),
.B(n_59),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2285),
.Y(n_2385)
);

INVx6_ASAP7_75t_L g2386 ( 
.A(n_2007),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2292),
.Y(n_2387)
);

AND2x2_ASAP7_75t_L g2388 ( 
.A(n_2092),
.B(n_58),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2073),
.B(n_2113),
.Y(n_2389)
);

NOR2xp33_ASAP7_75t_SL g2390 ( 
.A(n_2104),
.B(n_59),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2010),
.B(n_817),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2106),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2054),
.B(n_60),
.Y(n_2393)
);

BUFx4f_ASAP7_75t_L g2394 ( 
.A(n_2334),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2111),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2116),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_SL g2397 ( 
.A(n_2104),
.B(n_60),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2056),
.B(n_61),
.Y(n_2398)
);

BUFx3_ASAP7_75t_L g2399 ( 
.A(n_2334),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_2033),
.Y(n_2400)
);

OR2x2_ASAP7_75t_L g2401 ( 
.A(n_2184),
.B(n_2240),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2060),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_SL g2403 ( 
.A(n_2229),
.B(n_2237),
.Y(n_2403)
);

OR2x6_ASAP7_75t_L g2404 ( 
.A(n_2304),
.B(n_61),
.Y(n_2404)
);

AND2x4_ASAP7_75t_L g2405 ( 
.A(n_2203),
.B(n_2006),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2064),
.B(n_62),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2070),
.B(n_62),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2136),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2078),
.Y(n_2409)
);

BUFx8_ASAP7_75t_L g2410 ( 
.A(n_2321),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2140),
.Y(n_2411)
);

AND2x4_ASAP7_75t_L g2412 ( 
.A(n_2203),
.B(n_63),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2233),
.B(n_63),
.Y(n_2413)
);

AND2x4_ASAP7_75t_L g2414 ( 
.A(n_2213),
.B(n_2131),
.Y(n_2414)
);

BUFx12f_ASAP7_75t_L g2415 ( 
.A(n_2097),
.Y(n_2415)
);

AND2x4_ASAP7_75t_L g2416 ( 
.A(n_2213),
.B(n_64),
.Y(n_2416)
);

NAND2x1p5_ASAP7_75t_L g2417 ( 
.A(n_2118),
.B(n_65),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2093),
.Y(n_2418)
);

NAND2xp33_ASAP7_75t_L g2419 ( 
.A(n_2107),
.B(n_64),
.Y(n_2419)
);

OR2x2_ASAP7_75t_L g2420 ( 
.A(n_2184),
.B(n_66),
.Y(n_2420)
);

OR2x2_ASAP7_75t_L g2421 ( 
.A(n_2049),
.B(n_66),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2161),
.B(n_68),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2253),
.B(n_69),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2065),
.B(n_70),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2253),
.B(n_70),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_2311),
.Y(n_2426)
);

AND2x4_ASAP7_75t_L g2427 ( 
.A(n_2131),
.B(n_71),
.Y(n_2427)
);

INVx5_ASAP7_75t_L g2428 ( 
.A(n_2211),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_2107),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2066),
.B(n_71),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2164),
.B(n_72),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2038),
.B(n_2084),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2143),
.Y(n_2433)
);

OR2x6_ASAP7_75t_L g2434 ( 
.A(n_2137),
.B(n_72),
.Y(n_2434)
);

INVxp67_ASAP7_75t_SL g2435 ( 
.A(n_2137),
.Y(n_2435)
);

AND2x4_ASAP7_75t_L g2436 ( 
.A(n_2128),
.B(n_73),
.Y(n_2436)
);

BUFx4f_ASAP7_75t_L g2437 ( 
.A(n_2201),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_2107),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2013),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2151),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_2063),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2154),
.Y(n_2442)
);

BUFx6f_ASAP7_75t_L g2443 ( 
.A(n_2152),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_SL g2444 ( 
.A(n_2123),
.B(n_2147),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2069),
.B(n_74),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2157),
.Y(n_2446)
);

INVx1_ASAP7_75t_SL g2447 ( 
.A(n_2046),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2158),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2325),
.Y(n_2449)
);

AND2x4_ASAP7_75t_L g2450 ( 
.A(n_2013),
.B(n_75),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_2027),
.B(n_815),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2075),
.B(n_75),
.Y(n_2452)
);

BUFx6f_ASAP7_75t_L g2453 ( 
.A(n_2152),
.Y(n_2453)
);

AND2x4_ASAP7_75t_L g2454 ( 
.A(n_2075),
.B(n_76),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2084),
.B(n_77),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2171),
.Y(n_2456)
);

NAND2x1p5_ASAP7_75t_L g2457 ( 
.A(n_2103),
.B(n_79),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2193),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2198),
.Y(n_2459)
);

BUFx6f_ASAP7_75t_L g2460 ( 
.A(n_2152),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2105),
.B(n_2112),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2018),
.B(n_78),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_2028),
.B(n_78),
.Y(n_2463)
);

OR2x6_ASAP7_75t_L g2464 ( 
.A(n_2142),
.B(n_2148),
.Y(n_2464)
);

OR2x2_ASAP7_75t_L g2465 ( 
.A(n_2049),
.B(n_79),
.Y(n_2465)
);

AND2x4_ASAP7_75t_L g2466 ( 
.A(n_2232),
.B(n_80),
.Y(n_2466)
);

NAND2x1p5_ASAP7_75t_L g2467 ( 
.A(n_2147),
.B(n_81),
.Y(n_2467)
);

BUFx4f_ASAP7_75t_L g2468 ( 
.A(n_2246),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2176),
.B(n_80),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2202),
.Y(n_2470)
);

OR2x6_ASAP7_75t_L g2471 ( 
.A(n_2142),
.B(n_82),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_2148),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2028),
.B(n_83),
.Y(n_2473)
);

INVx5_ASAP7_75t_L g2474 ( 
.A(n_2211),
.Y(n_2474)
);

BUFx2_ASAP7_75t_L g2475 ( 
.A(n_2005),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2115),
.B(n_83),
.Y(n_2476)
);

INVx2_ASAP7_75t_SL g2477 ( 
.A(n_2001),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2244),
.Y(n_2478)
);

NAND2x1_ASAP7_75t_SL g2479 ( 
.A(n_2214),
.B(n_84),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2115),
.B(n_84),
.Y(n_2480)
);

BUFx2_ASAP7_75t_L g2481 ( 
.A(n_1996),
.Y(n_2481)
);

INVx3_ASAP7_75t_L g2482 ( 
.A(n_2325),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2266),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2216),
.Y(n_2484)
);

AND2x2_ASAP7_75t_L g2485 ( 
.A(n_2019),
.B(n_85),
.Y(n_2485)
);

AND2x4_ASAP7_75t_L g2486 ( 
.A(n_2232),
.B(n_85),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2231),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2266),
.Y(n_2488)
);

AND2x6_ASAP7_75t_L g2489 ( 
.A(n_2250),
.B(n_86),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2210),
.B(n_86),
.Y(n_2490)
);

OR2x6_ASAP7_75t_L g2491 ( 
.A(n_2250),
.B(n_2280),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2165),
.B(n_87),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2239),
.B(n_2245),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2247),
.B(n_87),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2021),
.B(n_89),
.Y(n_2495)
);

INVxp67_ASAP7_75t_L g2496 ( 
.A(n_2008),
.Y(n_2496)
);

AND2x4_ASAP7_75t_L g2497 ( 
.A(n_2247),
.B(n_89),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2303),
.Y(n_2498)
);

NOR2xp33_ASAP7_75t_L g2499 ( 
.A(n_2252),
.B(n_90),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2126),
.B(n_91),
.Y(n_2500)
);

AND2x6_ASAP7_75t_L g2501 ( 
.A(n_2207),
.B(n_92),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2159),
.B(n_92),
.Y(n_2502)
);

BUFx3_ASAP7_75t_L g2503 ( 
.A(n_2290),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2301),
.Y(n_2504)
);

AND2x4_ASAP7_75t_L g2505 ( 
.A(n_2265),
.B(n_93),
.Y(n_2505)
);

BUFx5_ASAP7_75t_L g2506 ( 
.A(n_2211),
.Y(n_2506)
);

BUFx6f_ASAP7_75t_L g2507 ( 
.A(n_2303),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2265),
.B(n_2215),
.Y(n_2508)
);

NAND2x1_ASAP7_75t_L g2509 ( 
.A(n_2303),
.B(n_93),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2043),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2043),
.Y(n_2511)
);

NOR2x1_ASAP7_75t_L g2512 ( 
.A(n_2256),
.B(n_2257),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2036),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2127),
.B(n_94),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2156),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2156),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2127),
.B(n_95),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2219),
.B(n_95),
.Y(n_2518)
);

BUFx6f_ASAP7_75t_L g2519 ( 
.A(n_2156),
.Y(n_2519)
);

INVx4_ASAP7_75t_L g2520 ( 
.A(n_2163),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2163),
.Y(n_2521)
);

AND2x4_ASAP7_75t_L g2522 ( 
.A(n_2220),
.B(n_2035),
.Y(n_2522)
);

NOR2xp33_ASAP7_75t_L g2523 ( 
.A(n_2044),
.B(n_2200),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2251),
.Y(n_2524)
);

AND2x4_ASAP7_75t_L g2525 ( 
.A(n_2039),
.B(n_96),
.Y(n_2525)
);

INVx1_ASAP7_75t_L g2526 ( 
.A(n_2041),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_SL g2527 ( 
.A(n_2071),
.B(n_96),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2025),
.B(n_98),
.Y(n_2528)
);

AO21x2_ASAP7_75t_L g2529 ( 
.A1(n_2088),
.A2(n_2316),
.B(n_2307),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2042),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_2029),
.B(n_826),
.Y(n_2531)
);

INVx4_ASAP7_75t_L g2532 ( 
.A(n_2163),
.Y(n_2532)
);

OR2x6_ASAP7_75t_L g2533 ( 
.A(n_2280),
.B(n_99),
.Y(n_2533)
);

NAND2x1_ASAP7_75t_SL g2534 ( 
.A(n_2214),
.B(n_100),
.Y(n_2534)
);

AND2x2_ASAP7_75t_L g2535 ( 
.A(n_2034),
.B(n_100),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2169),
.B(n_101),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2139),
.B(n_102),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2045),
.B(n_102),
.Y(n_2538)
);

BUFx12f_ASAP7_75t_L g2539 ( 
.A(n_2023),
.Y(n_2539)
);

OR2x2_ASAP7_75t_L g2540 ( 
.A(n_2291),
.B(n_103),
.Y(n_2540)
);

NAND2x1p5_ASAP7_75t_L g2541 ( 
.A(n_2109),
.B(n_2177),
.Y(n_2541)
);

OR2x2_ASAP7_75t_L g2542 ( 
.A(n_2212),
.B(n_2074),
.Y(n_2542)
);

AND2x2_ASAP7_75t_SL g2543 ( 
.A(n_2275),
.B(n_103),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2139),
.B(n_104),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_SL g2545 ( 
.A(n_2071),
.B(n_104),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2086),
.Y(n_2546)
);

OR2x6_ASAP7_75t_L g2547 ( 
.A(n_2101),
.B(n_2286),
.Y(n_2547)
);

AND2x2_ASAP7_75t_SL g2548 ( 
.A(n_2289),
.B(n_105),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2001),
.Y(n_2549)
);

BUFx6f_ASAP7_75t_L g2550 ( 
.A(n_2177),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2230),
.B(n_107),
.Y(n_2551)
);

INVx3_ASAP7_75t_L g2552 ( 
.A(n_2177),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2243),
.B(n_108),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2090),
.Y(n_2554)
);

INVx1_ASAP7_75t_SL g2555 ( 
.A(n_2302),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_L g2556 ( 
.A(n_2082),
.B(n_2031),
.Y(n_2556)
);

INVx5_ASAP7_75t_L g2557 ( 
.A(n_2211),
.Y(n_2557)
);

AND2x4_ASAP7_75t_L g2558 ( 
.A(n_2260),
.B(n_110),
.Y(n_2558)
);

AND2x6_ASAP7_75t_L g2559 ( 
.A(n_2207),
.B(n_110),
.Y(n_2559)
);

NAND2x1p5_ASAP7_75t_L g2560 ( 
.A(n_2162),
.B(n_112),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2310),
.Y(n_2561)
);

AND2x6_ASAP7_75t_L g2562 ( 
.A(n_2225),
.B(n_111),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2016),
.B(n_111),
.Y(n_2563)
);

AND2x4_ASAP7_75t_L g2564 ( 
.A(n_2263),
.B(n_112),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2182),
.B(n_113),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2037),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2166),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2183),
.B(n_113),
.Y(n_2568)
);

INVx6_ASAP7_75t_SL g2569 ( 
.A(n_2037),
.Y(n_2569)
);

AND2x6_ASAP7_75t_L g2570 ( 
.A(n_2225),
.B(n_115),
.Y(n_2570)
);

INVx3_ASAP7_75t_L g2571 ( 
.A(n_1998),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2145),
.B(n_115),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2145),
.B(n_116),
.Y(n_2573)
);

NOR2xp33_ASAP7_75t_SL g2574 ( 
.A(n_2071),
.B(n_116),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2189),
.B(n_2175),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2000),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2130),
.Y(n_2577)
);

INVxp67_ASAP7_75t_L g2578 ( 
.A(n_2040),
.Y(n_2578)
);

OR2x6_ASAP7_75t_L g2579 ( 
.A(n_2286),
.B(n_118),
.Y(n_2579)
);

INVx6_ASAP7_75t_L g2580 ( 
.A(n_2248),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2173),
.B(n_118),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2052),
.B(n_2055),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_SL g2583 ( 
.A(n_2071),
.B(n_119),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2052),
.B(n_120),
.Y(n_2584)
);

AND2x4_ASAP7_75t_L g2585 ( 
.A(n_2273),
.B(n_120),
.Y(n_2585)
);

HB1xp67_ASAP7_75t_L g2586 ( 
.A(n_2310),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2055),
.B(n_121),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2267),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2297),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2074),
.B(n_121),
.Y(n_2590)
);

AND2x4_ASAP7_75t_L g2591 ( 
.A(n_2298),
.B(n_122),
.Y(n_2591)
);

NOR2xp67_ASAP7_75t_L g2592 ( 
.A(n_2228),
.B(n_123),
.Y(n_2592)
);

BUFx2_ASAP7_75t_L g2593 ( 
.A(n_2297),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2057),
.B(n_123),
.Y(n_2594)
);

BUFx3_ASAP7_75t_L g2595 ( 
.A(n_2134),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2301),
.Y(n_2596)
);

INVx6_ASAP7_75t_L g2597 ( 
.A(n_2248),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2057),
.B(n_124),
.Y(n_2598)
);

AND2x4_ASAP7_75t_L g2599 ( 
.A(n_2002),
.B(n_124),
.Y(n_2599)
);

BUFx12f_ASAP7_75t_L g2600 ( 
.A(n_2032),
.Y(n_2600)
);

AND2x2_ASAP7_75t_SL g2601 ( 
.A(n_2186),
.B(n_126),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2281),
.B(n_126),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2083),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2283),
.B(n_127),
.Y(n_2604)
);

AND2x2_ASAP7_75t_L g2605 ( 
.A(n_2217),
.B(n_2221),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2299),
.B(n_127),
.Y(n_2606)
);

NAND2x1p5_ASAP7_75t_L g2607 ( 
.A(n_2024),
.B(n_2004),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2094),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2089),
.B(n_128),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_SL g2610 ( 
.A(n_2071),
.B(n_128),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2059),
.B(n_2067),
.Y(n_2611)
);

OR2x2_ASAP7_75t_L g2612 ( 
.A(n_2299),
.B(n_129),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2322),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2248),
.Y(n_2614)
);

INVx2_ASAP7_75t_SL g2615 ( 
.A(n_2087),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2059),
.B(n_130),
.Y(n_2616)
);

BUFx12f_ASAP7_75t_L g2617 ( 
.A(n_2087),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2083),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2309),
.B(n_131),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_2268),
.Y(n_2620)
);

BUFx4f_ASAP7_75t_L g2621 ( 
.A(n_2246),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2174),
.B(n_820),
.Y(n_2622)
);

INVx4_ASAP7_75t_L g2623 ( 
.A(n_2297),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_2009),
.B(n_132),
.Y(n_2624)
);

OR2x6_ASAP7_75t_L g2625 ( 
.A(n_2256),
.B(n_132),
.Y(n_2625)
);

BUFx6f_ASAP7_75t_L g2626 ( 
.A(n_2150),
.Y(n_2626)
);

AO21x2_ASAP7_75t_L g2627 ( 
.A1(n_2088),
.A2(n_133),
.B(n_134),
.Y(n_2627)
);

OR2x6_ASAP7_75t_L g2628 ( 
.A(n_2257),
.B(n_133),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_2296),
.Y(n_2629)
);

NOR2x1_ASAP7_75t_L g2630 ( 
.A(n_2294),
.B(n_135),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2015),
.B(n_135),
.Y(n_2631)
);

INVx3_ASAP7_75t_L g2632 ( 
.A(n_2306),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2110),
.Y(n_2633)
);

INVx4_ASAP7_75t_L g2634 ( 
.A(n_2297),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2067),
.B(n_136),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2110),
.Y(n_2636)
);

INVx5_ASAP7_75t_L g2637 ( 
.A(n_2211),
.Y(n_2637)
);

AND2x4_ASAP7_75t_L g2638 ( 
.A(n_2012),
.B(n_137),
.Y(n_2638)
);

NOR2xp33_ASAP7_75t_L g2639 ( 
.A(n_2174),
.B(n_828),
.Y(n_2639)
);

OR2x6_ASAP7_75t_L g2640 ( 
.A(n_2300),
.B(n_137),
.Y(n_2640)
);

AND2x4_ASAP7_75t_L g2641 ( 
.A(n_2014),
.B(n_138),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2258),
.B(n_832),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_1997),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2072),
.B(n_2146),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_1997),
.Y(n_2645)
);

HB1xp67_ASAP7_75t_L g2646 ( 
.A(n_2322),
.Y(n_2646)
);

AND2x2_ASAP7_75t_L g2647 ( 
.A(n_2318),
.B(n_138),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2296),
.B(n_2146),
.Y(n_2648)
);

NOR2x1_ASAP7_75t_SL g2649 ( 
.A(n_2323),
.B(n_139),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2100),
.Y(n_2650)
);

BUFx6f_ASAP7_75t_L g2651 ( 
.A(n_2314),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2072),
.B(n_140),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2305),
.B(n_141),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2279),
.B(n_141),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_SL g2655 ( 
.A(n_2246),
.B(n_142),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2317),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2308),
.B(n_142),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2058),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_2297),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2246),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2327),
.B(n_143),
.Y(n_2661)
);

OR2x6_ASAP7_75t_L g2662 ( 
.A(n_2100),
.B(n_144),
.Y(n_2662)
);

OR2x6_ASAP7_75t_L g2663 ( 
.A(n_2227),
.B(n_144),
.Y(n_2663)
);

BUFx2_ASAP7_75t_L g2664 ( 
.A(n_2328),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2333),
.Y(n_2665)
);

AND2x4_ASAP7_75t_L g2666 ( 
.A(n_2313),
.B(n_145),
.Y(n_2666)
);

AND2x6_ASAP7_75t_L g2667 ( 
.A(n_2326),
.B(n_2336),
.Y(n_2667)
);

CKINVDCx20_ASAP7_75t_R g2668 ( 
.A(n_2338),
.Y(n_2668)
);

NAND2xp5_ASAP7_75t_L g2669 ( 
.A(n_2053),
.B(n_145),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2053),
.B(n_146),
.Y(n_2670)
);

AND2x4_ASAP7_75t_L g2671 ( 
.A(n_2320),
.B(n_146),
.Y(n_2671)
);

NAND2x1p5_ASAP7_75t_L g2672 ( 
.A(n_2330),
.B(n_148),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2196),
.Y(n_2673)
);

NOR2xp33_ASAP7_75t_L g2674 ( 
.A(n_2254),
.B(n_817),
.Y(n_2674)
);

HB1xp67_ASAP7_75t_L g2675 ( 
.A(n_2323),
.Y(n_2675)
);

AND2x4_ASAP7_75t_L g2676 ( 
.A(n_2335),
.B(n_147),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2119),
.B(n_2144),
.Y(n_2677)
);

AND2x4_ASAP7_75t_L g2678 ( 
.A(n_2274),
.B(n_147),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2196),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2085),
.B(n_148),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2061),
.Y(n_2681)
);

BUFx2_ASAP7_75t_L g2682 ( 
.A(n_2337),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2051),
.Y(n_2683)
);

INVx1_ASAP7_75t_SL g2684 ( 
.A(n_2022),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2119),
.B(n_149),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2085),
.B(n_150),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2138),
.B(n_150),
.Y(n_2687)
);

INVx4_ASAP7_75t_L g2688 ( 
.A(n_2020),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2138),
.B(n_2234),
.Y(n_2689)
);

BUFx6f_ASAP7_75t_L g2690 ( 
.A(n_2295),
.Y(n_2690)
);

INVx3_ASAP7_75t_L g2691 ( 
.A(n_2181),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_L g2692 ( 
.A(n_2144),
.B(n_152),
.Y(n_2692)
);

OR2x6_ASAP7_75t_L g2693 ( 
.A(n_2262),
.B(n_152),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2254),
.B(n_831),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2274),
.B(n_154),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2141),
.B(n_154),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2222),
.Y(n_2697)
);

BUFx5_ASAP7_75t_L g2698 ( 
.A(n_2249),
.Y(n_2698)
);

BUFx6f_ASAP7_75t_L g2699 ( 
.A(n_2295),
.Y(n_2699)
);

NOR2xp33_ASAP7_75t_SL g2700 ( 
.A(n_2228),
.B(n_2241),
.Y(n_2700)
);

BUFx8_ASAP7_75t_L g2701 ( 
.A(n_2270),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2187),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2141),
.B(n_155),
.Y(n_2703)
);

AND2x4_ASAP7_75t_L g2704 ( 
.A(n_2282),
.B(n_155),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2197),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_2197),
.Y(n_2706)
);

AND2x4_ASAP7_75t_L g2707 ( 
.A(n_2117),
.B(n_156),
.Y(n_2707)
);

INVx3_ASAP7_75t_L g2708 ( 
.A(n_2190),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2284),
.Y(n_2709)
);

NOR2xp33_ASAP7_75t_L g2710 ( 
.A(n_2095),
.B(n_2108),
.Y(n_2710)
);

INVx6_ASAP7_75t_L g2711 ( 
.A(n_2272),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2324),
.B(n_156),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2199),
.Y(n_2713)
);

INVx5_ASAP7_75t_L g2714 ( 
.A(n_2295),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2167),
.B(n_157),
.Y(n_2715)
);

INVx5_ASAP7_75t_L g2716 ( 
.A(n_2284),
.Y(n_2716)
);

NOR2xp33_ASAP7_75t_L g2717 ( 
.A(n_2261),
.B(n_837),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2076),
.B(n_158),
.Y(n_2718)
);

INVx4_ASAP7_75t_L g2719 ( 
.A(n_2287),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2098),
.Y(n_2720)
);

BUFx6f_ASAP7_75t_L g2721 ( 
.A(n_2099),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2199),
.Y(n_2722)
);

INVx3_ASAP7_75t_L g2723 ( 
.A(n_2121),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2167),
.B(n_158),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2168),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2168),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2329),
.B(n_159),
.Y(n_2727)
);

NAND2x1_ASAP7_75t_L g2728 ( 
.A(n_2122),
.B(n_160),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2287),
.Y(n_2729)
);

AND2x4_ASAP7_75t_L g2730 ( 
.A(n_2261),
.B(n_160),
.Y(n_2730)
);

NOR2xp33_ASAP7_75t_SL g2731 ( 
.A(n_2178),
.B(n_162),
.Y(n_2731)
);

NOR2xp67_ASAP7_75t_L g2732 ( 
.A(n_2178),
.B(n_162),
.Y(n_2732)
);

AND2x6_ASAP7_75t_L g2733 ( 
.A(n_2124),
.B(n_163),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2172),
.Y(n_2734)
);

NOR2xp33_ASAP7_75t_L g2735 ( 
.A(n_2022),
.B(n_812),
.Y(n_2735)
);

BUFx3_ASAP7_75t_L g2736 ( 
.A(n_2180),
.Y(n_2736)
);

INVx5_ASAP7_75t_L g2737 ( 
.A(n_2272),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2262),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2208),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2208),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2172),
.Y(n_2741)
);

INVx6_ASAP7_75t_L g2742 ( 
.A(n_2272),
.Y(n_2742)
);

BUFx12f_ASAP7_75t_L g2743 ( 
.A(n_2293),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2188),
.B(n_163),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2223),
.Y(n_2745)
);

INVx3_ASAP7_75t_L g2746 ( 
.A(n_2124),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2188),
.Y(n_2747)
);

INVx4_ASAP7_75t_L g2748 ( 
.A(n_2255),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_SL g2749 ( 
.A(n_2307),
.B(n_164),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2194),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2153),
.B(n_164),
.Y(n_2751)
);

BUFx2_ASAP7_75t_L g2752 ( 
.A(n_2015),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2026),
.B(n_165),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_2026),
.Y(n_2754)
);

AND2x4_ASAP7_75t_L g2755 ( 
.A(n_2264),
.B(n_165),
.Y(n_2755)
);

NOR2xp67_ASAP7_75t_L g2756 ( 
.A(n_2259),
.B(n_166),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2223),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2226),
.Y(n_2758)
);

INVx4_ASAP7_75t_L g2759 ( 
.A(n_2205),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2194),
.Y(n_2760)
);

INVx3_ASAP7_75t_L g2761 ( 
.A(n_2206),
.Y(n_2761)
);

AND2x4_ASAP7_75t_L g2762 ( 
.A(n_2185),
.B(n_167),
.Y(n_2762)
);

BUFx6f_ASAP7_75t_L g2763 ( 
.A(n_2135),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2226),
.Y(n_2764)
);

OR2x6_ASAP7_75t_L g2765 ( 
.A(n_2294),
.B(n_2316),
.Y(n_2765)
);

AND2x4_ASAP7_75t_L g2766 ( 
.A(n_2185),
.B(n_169),
.Y(n_2766)
);

INVx4_ASAP7_75t_L g2767 ( 
.A(n_2125),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2120),
.B(n_2003),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2259),
.B(n_2120),
.Y(n_2769)
);

INVx6_ASAP7_75t_L g2770 ( 
.A(n_2242),
.Y(n_2770)
);

AND2x6_ASAP7_75t_L g2771 ( 
.A(n_2204),
.B(n_170),
.Y(n_2771)
);

AND2x4_ASAP7_75t_L g2772 ( 
.A(n_2278),
.B(n_170),
.Y(n_2772)
);

BUFx6f_ASAP7_75t_L g2773 ( 
.A(n_2236),
.Y(n_2773)
);

BUFx12f_ASAP7_75t_L g2774 ( 
.A(n_2242),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2003),
.B(n_172),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2288),
.Y(n_2776)
);

OR2x2_ASAP7_75t_L g2777 ( 
.A(n_2271),
.B(n_173),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2271),
.B(n_174),
.Y(n_2778)
);

AND2x2_ASAP7_75t_SL g2779 ( 
.A(n_2277),
.B(n_174),
.Y(n_2779)
);

BUFx6f_ASAP7_75t_L g2780 ( 
.A(n_2236),
.Y(n_2780)
);

INVx3_ASAP7_75t_L g2781 ( 
.A(n_2238),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2269),
.B(n_175),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2238),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2332),
.B(n_175),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2278),
.Y(n_2785)
);

AND2x4_ASAP7_75t_L g2786 ( 
.A(n_2277),
.B(n_176),
.Y(n_2786)
);

NAND2x1p5_ASAP7_75t_L g2787 ( 
.A(n_2209),
.B(n_177),
.Y(n_2787)
);

INVxp67_ASAP7_75t_L g2788 ( 
.A(n_2125),
.Y(n_2788)
);

BUFx2_ASAP7_75t_L g2789 ( 
.A(n_2288),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2204),
.Y(n_2790)
);

BUFx10_ASAP7_75t_L g2791 ( 
.A(n_2224),
.Y(n_2791)
);

CKINVDCx20_ASAP7_75t_R g2792 ( 
.A(n_2332),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2132),
.Y(n_2793)
);

NAND2x1p5_ASAP7_75t_L g2794 ( 
.A(n_2218),
.B(n_177),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2170),
.B(n_176),
.Y(n_2795)
);

INVx2_ASAP7_75t_SL g2796 ( 
.A(n_2334),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2047),
.B(n_179),
.Y(n_2797)
);

INVxp67_ASAP7_75t_SL g2798 ( 
.A(n_1999),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2048),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2129),
.Y(n_2800)
);

BUFx2_ASAP7_75t_L g2801 ( 
.A(n_1999),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2129),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2170),
.B(n_179),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2129),
.Y(n_2804)
);

BUFx6f_ASAP7_75t_L g2805 ( 
.A(n_2030),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2170),
.B(n_180),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2334),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2331),
.B(n_180),
.Y(n_2808)
);

AND2x4_ASAP7_75t_L g2809 ( 
.A(n_2047),
.B(n_181),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2048),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2334),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2129),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2030),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2048),
.Y(n_2814)
);

BUFx6f_ASAP7_75t_L g2815 ( 
.A(n_2030),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2170),
.B(n_181),
.Y(n_2816)
);

OR2x6_ASAP7_75t_L g2817 ( 
.A(n_2017),
.B(n_183),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2170),
.B(n_183),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2170),
.B(n_184),
.Y(n_2819)
);

BUFx6f_ASAP7_75t_L g2820 ( 
.A(n_2030),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2179),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2170),
.B(n_184),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2030),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2331),
.B(n_185),
.Y(n_2824)
);

NOR2xp33_ASAP7_75t_SL g2825 ( 
.A(n_2104),
.B(n_185),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2179),
.Y(n_2826)
);

CKINVDCx8_ASAP7_75t_R g2827 ( 
.A(n_2133),
.Y(n_2827)
);

CKINVDCx5p33_ASAP7_75t_R g2828 ( 
.A(n_2011),
.Y(n_2828)
);

BUFx2_ASAP7_75t_L g2829 ( 
.A(n_1999),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_1999),
.Y(n_2830)
);

CKINVDCx11_ASAP7_75t_R g2831 ( 
.A(n_2334),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2170),
.B(n_186),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_2334),
.Y(n_2833)
);

NOR2x1_ASAP7_75t_L g2834 ( 
.A(n_2319),
.B(n_186),
.Y(n_2834)
);

NAND2x1_ASAP7_75t_L g2835 ( 
.A(n_2030),
.B(n_187),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2331),
.B(n_187),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2331),
.B(n_188),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2331),
.B(n_188),
.Y(n_2838)
);

AND2x4_ASAP7_75t_L g2839 ( 
.A(n_2047),
.B(n_189),
.Y(n_2839)
);

INVxp67_ASAP7_75t_L g2840 ( 
.A(n_2312),
.Y(n_2840)
);

HB1xp67_ASAP7_75t_L g2841 ( 
.A(n_2331),
.Y(n_2841)
);

AND2x4_ASAP7_75t_L g2842 ( 
.A(n_2047),
.B(n_189),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2170),
.B(n_190),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2129),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2192),
.B(n_826),
.Y(n_2845)
);

INVx6_ASAP7_75t_L g2846 ( 
.A(n_2319),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2048),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2129),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2170),
.B(n_190),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2129),
.Y(n_2850)
);

HB1xp67_ASAP7_75t_L g2851 ( 
.A(n_2331),
.Y(n_2851)
);

INVxp67_ASAP7_75t_L g2852 ( 
.A(n_2312),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2331),
.B(n_191),
.Y(n_2853)
);

AND2x4_ASAP7_75t_L g2854 ( 
.A(n_2047),
.B(n_192),
.Y(n_2854)
);

CKINVDCx20_ASAP7_75t_R g2855 ( 
.A(n_2011),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2170),
.B(n_192),
.Y(n_2856)
);

AND2x4_ASAP7_75t_L g2857 ( 
.A(n_2047),
.B(n_193),
.Y(n_2857)
);

INVx3_ASAP7_75t_SL g2858 ( 
.A(n_2828),
.Y(n_2858)
);

BUFx8_ASAP7_75t_L g2859 ( 
.A(n_2539),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2346),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2701),
.Y(n_2861)
);

BUFx3_ASAP7_75t_L g2862 ( 
.A(n_2394),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2346),
.Y(n_2863)
);

BUFx6f_ASAP7_75t_L g2864 ( 
.A(n_2345),
.Y(n_2864)
);

CKINVDCx20_ASAP7_75t_R g2865 ( 
.A(n_2831),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2347),
.Y(n_2866)
);

CKINVDCx6p67_ASAP7_75t_R g2867 ( 
.A(n_2367),
.Y(n_2867)
);

BUFx3_ASAP7_75t_L g2868 ( 
.A(n_2394),
.Y(n_2868)
);

BUFx2_ASAP7_75t_L g2869 ( 
.A(n_2701),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2399),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2347),
.Y(n_2871)
);

INVx1_ASAP7_75t_SL g2872 ( 
.A(n_2351),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2799),
.Y(n_2873)
);

OR2x2_ASAP7_75t_L g2874 ( 
.A(n_2648),
.B(n_193),
.Y(n_2874)
);

INVx4_ASAP7_75t_L g2875 ( 
.A(n_2358),
.Y(n_2875)
);

INVx1_ASAP7_75t_SL g2876 ( 
.A(n_2801),
.Y(n_2876)
);

INVx3_ASAP7_75t_SL g2877 ( 
.A(n_2373),
.Y(n_2877)
);

BUFx3_ASAP7_75t_L g2878 ( 
.A(n_2807),
.Y(n_2878)
);

INVx3_ASAP7_75t_L g2879 ( 
.A(n_2623),
.Y(n_2879)
);

NOR2xp33_ASAP7_75t_L g2880 ( 
.A(n_2491),
.B(n_194),
.Y(n_2880)
);

INVx3_ASAP7_75t_L g2881 ( 
.A(n_2623),
.Y(n_2881)
);

AND2x2_ASAP7_75t_L g2882 ( 
.A(n_2380),
.B(n_194),
.Y(n_2882)
);

NAND2x1p5_ASAP7_75t_L g2883 ( 
.A(n_2833),
.B(n_2358),
.Y(n_2883)
);

BUFx3_ASAP7_75t_L g2884 ( 
.A(n_2410),
.Y(n_2884)
);

BUFx6f_ASAP7_75t_L g2885 ( 
.A(n_2345),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2799),
.B(n_195),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2810),
.Y(n_2887)
);

BUFx3_ASAP7_75t_L g2888 ( 
.A(n_2410),
.Y(n_2888)
);

INVx2_ASAP7_75t_SL g2889 ( 
.A(n_2415),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2855),
.Y(n_2890)
);

INVxp67_ASAP7_75t_SL g2891 ( 
.A(n_2810),
.Y(n_2891)
);

INVx3_ASAP7_75t_L g2892 ( 
.A(n_2634),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2814),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2814),
.Y(n_2894)
);

CKINVDCx11_ASAP7_75t_R g2895 ( 
.A(n_2367),
.Y(n_2895)
);

INVxp67_ASAP7_75t_SL g2896 ( 
.A(n_2847),
.Y(n_2896)
);

NAND2xp5_ASAP7_75t_L g2897 ( 
.A(n_2847),
.B(n_195),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2491),
.B(n_196),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2643),
.Y(n_2899)
);

INVx1_ASAP7_75t_SL g2900 ( 
.A(n_2829),
.Y(n_2900)
);

BUFx12f_ASAP7_75t_L g2901 ( 
.A(n_2817),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2725),
.B(n_196),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_2662),
.Y(n_2903)
);

BUFx6f_ASAP7_75t_SL g2904 ( 
.A(n_2817),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2643),
.Y(n_2905)
);

INVx6_ASAP7_75t_L g2906 ( 
.A(n_2386),
.Y(n_2906)
);

INVx3_ASAP7_75t_L g2907 ( 
.A(n_2634),
.Y(n_2907)
);

AOI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2792),
.A2(n_200),
.B1(n_197),
.B2(n_198),
.Y(n_2908)
);

CKINVDCx16_ASAP7_75t_R g2909 ( 
.A(n_2374),
.Y(n_2909)
);

CKINVDCx20_ASAP7_75t_R g2910 ( 
.A(n_2402),
.Y(n_2910)
);

BUFx6f_ASAP7_75t_L g2911 ( 
.A(n_2345),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2645),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2645),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2371),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_2662),
.Y(n_2915)
);

BUFx12f_ASAP7_75t_L g2916 ( 
.A(n_2404),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2371),
.Y(n_2917)
);

BUFx2_ASAP7_75t_R g2918 ( 
.A(n_2620),
.Y(n_2918)
);

INVx4_ASAP7_75t_L g2919 ( 
.A(n_2374),
.Y(n_2919)
);

BUFx3_ASAP7_75t_L g2920 ( 
.A(n_2386),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2403),
.B(n_197),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2821),
.Y(n_2922)
);

INVx1_ASAP7_75t_SL g2923 ( 
.A(n_2830),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2343),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2800),
.Y(n_2925)
);

INVxp67_ASAP7_75t_SL g2926 ( 
.A(n_2450),
.Y(n_2926)
);

BUFx2_ASAP7_75t_L g2927 ( 
.A(n_2569),
.Y(n_2927)
);

INVx3_ASAP7_75t_SL g2928 ( 
.A(n_2504),
.Y(n_2928)
);

NAND2x1p5_ASAP7_75t_L g2929 ( 
.A(n_2796),
.B(n_198),
.Y(n_2929)
);

BUFx2_ASAP7_75t_R g2930 ( 
.A(n_2596),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2802),
.Y(n_2931)
);

BUFx2_ASAP7_75t_SL g2932 ( 
.A(n_2366),
.Y(n_2932)
);

BUFx6f_ASAP7_75t_L g2933 ( 
.A(n_2348),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2379),
.Y(n_2934)
);

BUFx4_ASAP7_75t_SL g2935 ( 
.A(n_2404),
.Y(n_2935)
);

BUFx3_ASAP7_75t_L g2936 ( 
.A(n_2617),
.Y(n_2936)
);

OAI22xp5_ASAP7_75t_L g2937 ( 
.A1(n_2437),
.A2(n_203),
.B1(n_200),
.B2(n_202),
.Y(n_2937)
);

BUFx6f_ASAP7_75t_L g2938 ( 
.A(n_2348),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_L g2939 ( 
.A(n_2348),
.Y(n_2939)
);

BUFx12f_ASAP7_75t_L g2940 ( 
.A(n_2533),
.Y(n_2940)
);

BUFx8_ASAP7_75t_L g2941 ( 
.A(n_2600),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2826),
.Y(n_2942)
);

BUFx3_ASAP7_75t_L g2943 ( 
.A(n_2811),
.Y(n_2943)
);

INVx1_ASAP7_75t_SL g2944 ( 
.A(n_2841),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2379),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2392),
.Y(n_2946)
);

INVx5_ASAP7_75t_L g2947 ( 
.A(n_2471),
.Y(n_2947)
);

BUFx2_ASAP7_75t_SL g2948 ( 
.A(n_2827),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2392),
.Y(n_2949)
);

OR2x6_ASAP7_75t_L g2950 ( 
.A(n_2471),
.B(n_205),
.Y(n_2950)
);

INVx2_ASAP7_75t_SL g2951 ( 
.A(n_2846),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2395),
.Y(n_2952)
);

INVx6_ASAP7_75t_L g2953 ( 
.A(n_2846),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2851),
.Y(n_2954)
);

INVx1_ASAP7_75t_SL g2955 ( 
.A(n_2447),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2389),
.B(n_206),
.Y(n_2956)
);

INVx1_ASAP7_75t_SL g2957 ( 
.A(n_2368),
.Y(n_2957)
);

BUFx3_ASAP7_75t_L g2958 ( 
.A(n_2472),
.Y(n_2958)
);

BUFx6f_ASAP7_75t_L g2959 ( 
.A(n_2365),
.Y(n_2959)
);

CKINVDCx20_ASAP7_75t_R g2960 ( 
.A(n_2503),
.Y(n_2960)
);

NAND2x1p5_ASAP7_75t_L g2961 ( 
.A(n_2437),
.B(n_207),
.Y(n_2961)
);

OR2x2_ASAP7_75t_L g2962 ( 
.A(n_2382),
.B(n_207),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2395),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2396),
.Y(n_2964)
);

INVx6_ASAP7_75t_SL g2965 ( 
.A(n_2434),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2396),
.Y(n_2966)
);

INVx1_ASAP7_75t_SL g2967 ( 
.A(n_2354),
.Y(n_2967)
);

INVx2_ASAP7_75t_L g2968 ( 
.A(n_2804),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2812),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2844),
.Y(n_2970)
);

NAND2xp5_ASAP7_75t_L g2971 ( 
.A(n_2726),
.B(n_208),
.Y(n_2971)
);

INVx3_ASAP7_75t_L g2972 ( 
.A(n_2405),
.Y(n_2972)
);

INVx4_ASAP7_75t_L g2973 ( 
.A(n_2434),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2440),
.Y(n_2974)
);

INVx3_ASAP7_75t_SL g2975 ( 
.A(n_2533),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_2464),
.Y(n_2976)
);

BUFx2_ASAP7_75t_L g2977 ( 
.A(n_2569),
.Y(n_2977)
);

BUFx2_ASAP7_75t_L g2978 ( 
.A(n_2414),
.Y(n_2978)
);

BUFx2_ASAP7_75t_L g2979 ( 
.A(n_2414),
.Y(n_2979)
);

INVx3_ASAP7_75t_L g2980 ( 
.A(n_2405),
.Y(n_2980)
);

NAND2x1p5_ASAP7_75t_L g2981 ( 
.A(n_2719),
.B(n_2468),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2734),
.B(n_209),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2440),
.Y(n_2983)
);

OR2x6_ASAP7_75t_L g2984 ( 
.A(n_2579),
.B(n_211),
.Y(n_2984)
);

INVx3_ASAP7_75t_SL g2985 ( 
.A(n_2579),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2741),
.B(n_212),
.Y(n_2986)
);

INVx1_ASAP7_75t_SL g2987 ( 
.A(n_2364),
.Y(n_2987)
);

BUFx4_ASAP7_75t_SL g2988 ( 
.A(n_2640),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2848),
.Y(n_2989)
);

NAND2x1p5_ASAP7_75t_L g2990 ( 
.A(n_2719),
.B(n_2468),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2850),
.Y(n_2991)
);

BUFx12f_ASAP7_75t_L g2992 ( 
.A(n_2640),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2408),
.Y(n_2993)
);

INVx2_ASAP7_75t_SL g2994 ( 
.A(n_2464),
.Y(n_2994)
);

BUFx6f_ASAP7_75t_L g2995 ( 
.A(n_2365),
.Y(n_2995)
);

NOR2xp33_ASAP7_75t_L g2996 ( 
.A(n_2578),
.B(n_213),
.Y(n_2996)
);

BUFx2_ASAP7_75t_SL g2997 ( 
.A(n_2489),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2456),
.Y(n_2998)
);

BUFx8_ASAP7_75t_L g2999 ( 
.A(n_2364),
.Y(n_2999)
);

BUFx6f_ASAP7_75t_L g3000 ( 
.A(n_2365),
.Y(n_3000)
);

INVx6_ASAP7_75t_SL g3001 ( 
.A(n_2663),
.Y(n_3001)
);

OR2x6_ASAP7_75t_L g3002 ( 
.A(n_2693),
.B(n_214),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2456),
.Y(n_3003)
);

BUFx2_ASAP7_75t_SL g3004 ( 
.A(n_2489),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2429),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2411),
.Y(n_3006)
);

BUFx2_ASAP7_75t_L g3007 ( 
.A(n_2798),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2747),
.B(n_215),
.Y(n_3008)
);

AND2x2_ASAP7_75t_L g3009 ( 
.A(n_2461),
.B(n_215),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2750),
.B(n_216),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2458),
.Y(n_3011)
);

BUFx12f_ASAP7_75t_L g3012 ( 
.A(n_2629),
.Y(n_3012)
);

BUFx3_ASAP7_75t_L g3013 ( 
.A(n_2441),
.Y(n_3013)
);

INVx3_ASAP7_75t_L g3014 ( 
.A(n_2659),
.Y(n_3014)
);

BUFx8_ASAP7_75t_L g3015 ( 
.A(n_2743),
.Y(n_3015)
);

NOR2xp67_ASAP7_75t_SL g3016 ( 
.A(n_2428),
.B(n_216),
.Y(n_3016)
);

INVx4_ASAP7_75t_L g3017 ( 
.A(n_2489),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2595),
.Y(n_3018)
);

BUFx2_ASAP7_75t_SL g3019 ( 
.A(n_2489),
.Y(n_3019)
);

INVx1_ASAP7_75t_SL g3020 ( 
.A(n_2383),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2458),
.Y(n_3021)
);

BUFx2_ASAP7_75t_SL g3022 ( 
.A(n_2427),
.Y(n_3022)
);

BUFx8_ASAP7_75t_L g3023 ( 
.A(n_2481),
.Y(n_3023)
);

BUFx2_ASAP7_75t_SL g3024 ( 
.A(n_2427),
.Y(n_3024)
);

BUFx6f_ASAP7_75t_L g3025 ( 
.A(n_2429),
.Y(n_3025)
);

NAND2x1p5_ASAP7_75t_L g3026 ( 
.A(n_2621),
.B(n_217),
.Y(n_3026)
);

BUFx3_ASAP7_75t_L g3027 ( 
.A(n_2709),
.Y(n_3027)
);

BUFx3_ASAP7_75t_L g3028 ( 
.A(n_2547),
.Y(n_3028)
);

INVx4_ASAP7_75t_L g3029 ( 
.A(n_2621),
.Y(n_3029)
);

BUFx3_ASAP7_75t_L g3030 ( 
.A(n_2547),
.Y(n_3030)
);

INVx6_ASAP7_75t_SL g3031 ( 
.A(n_2663),
.Y(n_3031)
);

NAND2x1p5_ASAP7_75t_L g3032 ( 
.A(n_2714),
.B(n_218),
.Y(n_3032)
);

BUFx6f_ASAP7_75t_L g3033 ( 
.A(n_2429),
.Y(n_3033)
);

BUFx6f_ASAP7_75t_SL g3034 ( 
.A(n_2543),
.Y(n_3034)
);

BUFx2_ASAP7_75t_SL g3035 ( 
.A(n_2729),
.Y(n_3035)
);

BUFx2_ASAP7_75t_L g3036 ( 
.A(n_2840),
.Y(n_3036)
);

INVx4_ASAP7_75t_L g3037 ( 
.A(n_2714),
.Y(n_3037)
);

INVx1_ASAP7_75t_SL g3038 ( 
.A(n_2416),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_2452),
.Y(n_3039)
);

CKINVDCx20_ASAP7_75t_R g3040 ( 
.A(n_2668),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2523),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_3041)
);

NAND2x1p5_ASAP7_75t_L g3042 ( 
.A(n_2714),
.B(n_219),
.Y(n_3042)
);

BUFx6f_ASAP7_75t_L g3043 ( 
.A(n_2438),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2433),
.Y(n_3044)
);

BUFx6f_ASAP7_75t_L g3045 ( 
.A(n_2438),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2438),
.Y(n_3046)
);

INVx1_ASAP7_75t_SL g3047 ( 
.A(n_2416),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2493),
.Y(n_3048)
);

INVx3_ASAP7_75t_SL g3049 ( 
.A(n_2548),
.Y(n_3049)
);

NAND2xp5_ASAP7_75t_SL g3050 ( 
.A(n_2444),
.B(n_220),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2510),
.Y(n_3051)
);

BUFx3_ASAP7_75t_L g3052 ( 
.A(n_2452),
.Y(n_3052)
);

CKINVDCx6p67_ASAP7_75t_R g3053 ( 
.A(n_2693),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2454),
.Y(n_3054)
);

INVx5_ASAP7_75t_L g3055 ( 
.A(n_2516),
.Y(n_3055)
);

INVxp67_ASAP7_75t_SL g3056 ( 
.A(n_2450),
.Y(n_3056)
);

OR2x6_ASAP7_75t_L g3057 ( 
.A(n_2384),
.B(n_222),
.Y(n_3057)
);

BUFx2_ASAP7_75t_L g3058 ( 
.A(n_2852),
.Y(n_3058)
);

BUFx6f_ASAP7_75t_L g3059 ( 
.A(n_2443),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2454),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2442),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2510),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2511),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2767),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2511),
.Y(n_3065)
);

BUFx12f_ASAP7_75t_L g3066 ( 
.A(n_2417),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2603),
.Y(n_3067)
);

INVx5_ASAP7_75t_L g3068 ( 
.A(n_2516),
.Y(n_3068)
);

BUFx3_ASAP7_75t_L g3069 ( 
.A(n_2580),
.Y(n_3069)
);

BUFx6f_ASAP7_75t_L g3070 ( 
.A(n_2443),
.Y(n_3070)
);

NAND2x1p5_ASAP7_75t_L g3071 ( 
.A(n_2412),
.B(n_224),
.Y(n_3071)
);

BUFx12f_ASAP7_75t_L g3072 ( 
.A(n_2401),
.Y(n_3072)
);

INVx2_ASAP7_75t_SL g3073 ( 
.A(n_2716),
.Y(n_3073)
);

INVx3_ASAP7_75t_L g3074 ( 
.A(n_2767),
.Y(n_3074)
);

OR2x6_ASAP7_75t_L g3075 ( 
.A(n_2560),
.B(n_225),
.Y(n_3075)
);

INVxp67_ASAP7_75t_SL g3076 ( 
.A(n_2378),
.Y(n_3076)
);

INVx1_ASAP7_75t_SL g3077 ( 
.A(n_2824),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2677),
.B(n_225),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2446),
.Y(n_3079)
);

NOR2xp33_ASAP7_75t_L g3080 ( 
.A(n_2542),
.B(n_226),
.Y(n_3080)
);

CKINVDCx6p67_ASAP7_75t_R g3081 ( 
.A(n_2601),
.Y(n_3081)
);

BUFx6f_ASAP7_75t_L g3082 ( 
.A(n_2443),
.Y(n_3082)
);

INVx3_ASAP7_75t_SL g3083 ( 
.A(n_2341),
.Y(n_3083)
);

BUFx6f_ASAP7_75t_L g3084 ( 
.A(n_2453),
.Y(n_3084)
);

BUFx12f_ASAP7_75t_L g3085 ( 
.A(n_2421),
.Y(n_3085)
);

INVx1_ASAP7_75t_SL g3086 ( 
.A(n_2412),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2760),
.B(n_227),
.Y(n_3087)
);

INVxp67_ASAP7_75t_SL g3088 ( 
.A(n_2439),
.Y(n_3088)
);

INVx3_ASAP7_75t_L g3089 ( 
.A(n_2520),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_2475),
.B(n_228),
.Y(n_3090)
);

INVx5_ASAP7_75t_L g3091 ( 
.A(n_2516),
.Y(n_3091)
);

BUFx2_ASAP7_75t_L g3092 ( 
.A(n_2435),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2603),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2618),
.Y(n_3094)
);

BUFx6f_ASAP7_75t_L g3095 ( 
.A(n_2453),
.Y(n_3095)
);

AOI22xp33_ASAP7_75t_L g3096 ( 
.A1(n_2556),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2466),
.Y(n_3097)
);

INVx2_ASAP7_75t_SL g3098 ( 
.A(n_2716),
.Y(n_3098)
);

NOR2xp33_ASAP7_75t_L g3099 ( 
.A(n_2496),
.B(n_229),
.Y(n_3099)
);

BUFx2_ASAP7_75t_SL g3100 ( 
.A(n_2466),
.Y(n_3100)
);

INVx2_ASAP7_75t_SL g3101 ( 
.A(n_2716),
.Y(n_3101)
);

BUFx6f_ASAP7_75t_L g3102 ( 
.A(n_2453),
.Y(n_3102)
);

CKINVDCx20_ASAP7_75t_R g3103 ( 
.A(n_2400),
.Y(n_3103)
);

INVx4_ASAP7_75t_L g3104 ( 
.A(n_2519),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2448),
.Y(n_3105)
);

INVx5_ASAP7_75t_L g3106 ( 
.A(n_2519),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2618),
.Y(n_3107)
);

INVx5_ASAP7_75t_L g3108 ( 
.A(n_2519),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2432),
.B(n_230),
.Y(n_3109)
);

CKINVDCx16_ASAP7_75t_R g3110 ( 
.A(n_2390),
.Y(n_3110)
);

BUFx4f_ASAP7_75t_L g3111 ( 
.A(n_2733),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2459),
.Y(n_3112)
);

INVx1_ASAP7_75t_SL g3113 ( 
.A(n_2339),
.Y(n_3113)
);

AND2x6_ASAP7_75t_L g3114 ( 
.A(n_2650),
.B(n_231),
.Y(n_3114)
);

INVx3_ASAP7_75t_L g3115 ( 
.A(n_2520),
.Y(n_3115)
);

BUFx2_ASAP7_75t_L g3116 ( 
.A(n_2486),
.Y(n_3116)
);

BUFx3_ASAP7_75t_L g3117 ( 
.A(n_2580),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2492),
.B(n_232),
.Y(n_3118)
);

INVx1_ASAP7_75t_SL g3119 ( 
.A(n_2353),
.Y(n_3119)
);

INVxp67_ASAP7_75t_SL g3120 ( 
.A(n_2599),
.Y(n_3120)
);

AND2x4_ASAP7_75t_L g3121 ( 
.A(n_2650),
.B(n_232),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2633),
.Y(n_3122)
);

INVx3_ASAP7_75t_L g3123 ( 
.A(n_2532),
.Y(n_3123)
);

BUFx3_ASAP7_75t_L g3124 ( 
.A(n_2597),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2774),
.Y(n_3125)
);

BUFx3_ASAP7_75t_L g3126 ( 
.A(n_2597),
.Y(n_3126)
);

OAI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2625),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_3127)
);

BUFx12f_ASAP7_75t_L g3128 ( 
.A(n_2465),
.Y(n_3128)
);

INVx3_ASAP7_75t_SL g3129 ( 
.A(n_2341),
.Y(n_3129)
);

BUFx4_ASAP7_75t_SL g3130 ( 
.A(n_2420),
.Y(n_3130)
);

INVx3_ASAP7_75t_SL g3131 ( 
.A(n_2350),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2633),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2636),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2575),
.B(n_234),
.Y(n_3134)
);

NAND2x1p5_ASAP7_75t_L g3135 ( 
.A(n_2428),
.B(n_2474),
.Y(n_3135)
);

BUFx4f_ASAP7_75t_SL g3136 ( 
.A(n_2678),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_SL g3137 ( 
.A(n_2678),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_L g3138 ( 
.A1(n_2779),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_3138)
);

BUFx2_ASAP7_75t_SL g3139 ( 
.A(n_2486),
.Y(n_3139)
);

INVx5_ASAP7_75t_L g3140 ( 
.A(n_2550),
.Y(n_3140)
);

HB1xp67_ASAP7_75t_L g3141 ( 
.A(n_2494),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2636),
.Y(n_3142)
);

INVx3_ASAP7_75t_SL g3143 ( 
.A(n_2350),
.Y(n_3143)
);

OAI22xp5_ASAP7_75t_L g3144 ( 
.A1(n_2625),
.A2(n_240),
.B1(n_237),
.B2(n_238),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2644),
.B(n_238),
.Y(n_3145)
);

CKINVDCx11_ASAP7_75t_R g3146 ( 
.A(n_2695),
.Y(n_3146)
);

INVx3_ASAP7_75t_SL g3147 ( 
.A(n_2797),
.Y(n_3147)
);

BUFx2_ASAP7_75t_L g3148 ( 
.A(n_2494),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2577),
.Y(n_3149)
);

BUFx2_ASAP7_75t_SL g3150 ( 
.A(n_2497),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2470),
.Y(n_3151)
);

OAI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_2628),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_3152)
);

INVx5_ASAP7_75t_L g3153 ( 
.A(n_2550),
.Y(n_3153)
);

INVx1_ASAP7_75t_SL g3154 ( 
.A(n_2808),
.Y(n_3154)
);

INVx5_ASAP7_75t_L g3155 ( 
.A(n_2550),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2460),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2582),
.B(n_243),
.Y(n_3157)
);

BUFx2_ASAP7_75t_SL g3158 ( 
.A(n_2497),
.Y(n_3158)
);

INVx1_ASAP7_75t_SL g3159 ( 
.A(n_2836),
.Y(n_3159)
);

BUFx3_ASAP7_75t_L g3160 ( 
.A(n_2577),
.Y(n_3160)
);

INVx5_ASAP7_75t_L g3161 ( 
.A(n_2460),
.Y(n_3161)
);

INVx1_ASAP7_75t_SL g3162 ( 
.A(n_2837),
.Y(n_3162)
);

AOI22xp33_ASAP7_75t_L g3163 ( 
.A1(n_2499),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2484),
.Y(n_3164)
);

BUFx12f_ASAP7_75t_L g3165 ( 
.A(n_2718),
.Y(n_3165)
);

BUFx2_ASAP7_75t_L g3166 ( 
.A(n_2505),
.Y(n_3166)
);

INVx2_ASAP7_75t_SL g3167 ( 
.A(n_2505),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2487),
.Y(n_3168)
);

INVx1_ASAP7_75t_SL g3169 ( 
.A(n_2838),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2381),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2577),
.Y(n_3171)
);

INVx1_ASAP7_75t_SL g3172 ( 
.A(n_2853),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_2626),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_2409),
.Y(n_3174)
);

BUFx3_ASAP7_75t_L g3175 ( 
.A(n_2626),
.Y(n_3175)
);

INVx5_ASAP7_75t_SL g3176 ( 
.A(n_2797),
.Y(n_3176)
);

BUFx8_ASAP7_75t_L g3177 ( 
.A(n_2695),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2611),
.B(n_244),
.Y(n_3178)
);

INVx2_ASAP7_75t_R g3179 ( 
.A(n_2428),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2508),
.B(n_245),
.Y(n_3180)
);

BUFx6f_ASAP7_75t_SL g3181 ( 
.A(n_2730),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2385),
.Y(n_3182)
);

BUFx6f_ASAP7_75t_L g3183 ( 
.A(n_2460),
.Y(n_3183)
);

INVx5_ASAP7_75t_L g3184 ( 
.A(n_2498),
.Y(n_3184)
);

INVx2_ASAP7_75t_SL g3185 ( 
.A(n_2585),
.Y(n_3185)
);

AND2x2_ASAP7_75t_L g3186 ( 
.A(n_2469),
.B(n_246),
.Y(n_3186)
);

BUFx3_ASAP7_75t_L g3187 ( 
.A(n_2626),
.Y(n_3187)
);

BUFx12f_ASAP7_75t_L g3188 ( 
.A(n_2436),
.Y(n_3188)
);

INVx2_ASAP7_75t_SL g3189 ( 
.A(n_2585),
.Y(n_3189)
);

BUFx3_ASAP7_75t_L g3190 ( 
.A(n_2508),
.Y(n_3190)
);

BUFx6f_ASAP7_75t_L g3191 ( 
.A(n_2498),
.Y(n_3191)
);

BUFx3_ASAP7_75t_L g3192 ( 
.A(n_2522),
.Y(n_3192)
);

INVx4_ASAP7_75t_L g3193 ( 
.A(n_2474),
.Y(n_3193)
);

NAND2x1p5_ASAP7_75t_L g3194 ( 
.A(n_2474),
.B(n_246),
.Y(n_3194)
);

BUFx4_ASAP7_75t_SL g3195 ( 
.A(n_2540),
.Y(n_3195)
);

BUFx2_ASAP7_75t_L g3196 ( 
.A(n_2413),
.Y(n_3196)
);

BUFx3_ASAP7_75t_L g3197 ( 
.A(n_2522),
.Y(n_3197)
);

INVx3_ASAP7_75t_L g3198 ( 
.A(n_2532),
.Y(n_3198)
);

BUFx2_ASAP7_75t_L g3199 ( 
.A(n_2413),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2524),
.B(n_247),
.Y(n_3200)
);

AOI22xp33_ASAP7_75t_L g3201 ( 
.A1(n_2704),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_3201)
);

BUFx2_ASAP7_75t_L g3202 ( 
.A(n_2704),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2387),
.Y(n_3203)
);

CKINVDCx8_ASAP7_75t_R g3204 ( 
.A(n_2733),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2418),
.Y(n_3205)
);

NAND2x1p5_ASAP7_75t_L g3206 ( 
.A(n_2557),
.B(n_248),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2526),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2344),
.Y(n_3208)
);

INVx3_ASAP7_75t_L g3209 ( 
.A(n_2498),
.Y(n_3209)
);

INVx2_ASAP7_75t_SL g3210 ( 
.A(n_2809),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2355),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2507),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2513),
.Y(n_3213)
);

BUFx6f_ASAP7_75t_L g3214 ( 
.A(n_2507),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2530),
.Y(n_3215)
);

BUFx4_ASAP7_75t_SL g3216 ( 
.A(n_2606),
.Y(n_3216)
);

CKINVDCx20_ASAP7_75t_R g3217 ( 
.A(n_2612),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2658),
.Y(n_3218)
);

BUFx6f_ASAP7_75t_L g3219 ( 
.A(n_2507),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2349),
.Y(n_3220)
);

CKINVDCx11_ASAP7_75t_R g3221 ( 
.A(n_2436),
.Y(n_3221)
);

INVx2_ASAP7_75t_SL g3222 ( 
.A(n_2809),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2805),
.Y(n_3223)
);

BUFx6f_ASAP7_75t_L g3224 ( 
.A(n_2805),
.Y(n_3224)
);

BUFx5_ASAP7_75t_L g3225 ( 
.A(n_2667),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2681),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_2805),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_2599),
.Y(n_3228)
);

INVxp67_ASAP7_75t_SL g3229 ( 
.A(n_2624),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2684),
.B(n_251),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2683),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2357),
.Y(n_3232)
);

BUFx6f_ASAP7_75t_L g3233 ( 
.A(n_2813),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_2362),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_2624),
.Y(n_3235)
);

INVx3_ASAP7_75t_L g3236 ( 
.A(n_2813),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2370),
.Y(n_3237)
);

INVx5_ASAP7_75t_L g3238 ( 
.A(n_2813),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_L g3239 ( 
.A(n_2710),
.B(n_252),
.Y(n_3239)
);

INVx2_ASAP7_75t_SL g3240 ( 
.A(n_2839),
.Y(n_3240)
);

OR2x6_ASAP7_75t_L g3241 ( 
.A(n_2525),
.B(n_252),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2546),
.Y(n_3242)
);

BUFx3_ASAP7_75t_L g3243 ( 
.A(n_2839),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2554),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_2842),
.Y(n_3245)
);

INVx2_ASAP7_75t_L g3246 ( 
.A(n_2608),
.Y(n_3246)
);

BUFx12f_ASAP7_75t_L g3247 ( 
.A(n_2457),
.Y(n_3247)
);

INVxp67_ASAP7_75t_SL g3248 ( 
.A(n_2638),
.Y(n_3248)
);

CKINVDCx5p33_ASAP7_75t_R g3249 ( 
.A(n_2842),
.Y(n_3249)
);

BUFx3_ASAP7_75t_L g3250 ( 
.A(n_2854),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2588),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_2567),
.Y(n_3252)
);

INVxp67_ASAP7_75t_SL g3253 ( 
.A(n_2638),
.Y(n_3253)
);

BUFx2_ASAP7_75t_SL g3254 ( 
.A(n_2641),
.Y(n_3254)
);

BUFx2_ASAP7_75t_L g3255 ( 
.A(n_2641),
.Y(n_3255)
);

CKINVDCx16_ASAP7_75t_R g3256 ( 
.A(n_2397),
.Y(n_3256)
);

INVx5_ASAP7_75t_L g3257 ( 
.A(n_2815),
.Y(n_3257)
);

INVx3_ASAP7_75t_L g3258 ( 
.A(n_2815),
.Y(n_3258)
);

INVx3_ASAP7_75t_L g3259 ( 
.A(n_2815),
.Y(n_3259)
);

INVx6_ASAP7_75t_SL g3260 ( 
.A(n_2854),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2483),
.Y(n_3261)
);

CKINVDCx11_ASAP7_75t_R g3262 ( 
.A(n_2857),
.Y(n_3262)
);

CKINVDCx5p33_ASAP7_75t_R g3263 ( 
.A(n_2857),
.Y(n_3263)
);

AND2x4_ASAP7_75t_L g3264 ( 
.A(n_2589),
.B(n_253),
.Y(n_3264)
);

INVx5_ASAP7_75t_L g3265 ( 
.A(n_2820),
.Y(n_3265)
);

INVx6_ASAP7_75t_SL g3266 ( 
.A(n_2525),
.Y(n_3266)
);

BUFx12f_ASAP7_75t_L g3267 ( 
.A(n_2730),
.Y(n_3267)
);

BUFx3_ASAP7_75t_L g3268 ( 
.A(n_2538),
.Y(n_3268)
);

BUFx12f_ASAP7_75t_L g3269 ( 
.A(n_2538),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2488),
.Y(n_3270)
);

OR2x2_ASAP7_75t_L g3271 ( 
.A(n_2359),
.B(n_253),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_2593),
.B(n_254),
.Y(n_3272)
);

BUFx24_ASAP7_75t_L g3273 ( 
.A(n_2653),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_2736),
.Y(n_3274)
);

BUFx6f_ASAP7_75t_L g3275 ( 
.A(n_2820),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2769),
.Y(n_3276)
);

INVx5_ASAP7_75t_L g3277 ( 
.A(n_2820),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2642),
.B(n_254),
.Y(n_3278)
);

BUFx4f_ASAP7_75t_SL g3279 ( 
.A(n_2477),
.Y(n_3279)
);

BUFx3_ASAP7_75t_L g3280 ( 
.A(n_2653),
.Y(n_3280)
);

NAND2x1p5_ASAP7_75t_L g3281 ( 
.A(n_2557),
.B(n_255),
.Y(n_3281)
);

BUFx3_ASAP7_75t_L g3282 ( 
.A(n_2657),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2746),
.Y(n_3283)
);

BUFx3_ASAP7_75t_L g3284 ( 
.A(n_2657),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2673),
.Y(n_3285)
);

BUFx6f_ASAP7_75t_L g3286 ( 
.A(n_2823),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2673),
.Y(n_3287)
);

NAND2x1p5_ASAP7_75t_L g3288 ( 
.A(n_2557),
.B(n_255),
.Y(n_3288)
);

BUFx6f_ASAP7_75t_L g3289 ( 
.A(n_2823),
.Y(n_3289)
);

AND2x4_ASAP7_75t_L g3290 ( 
.A(n_2754),
.B(n_256),
.Y(n_3290)
);

BUFx6f_ASAP7_75t_SL g3291 ( 
.A(n_2591),
.Y(n_3291)
);

BUFx6f_ASAP7_75t_L g3292 ( 
.A(n_2823),
.Y(n_3292)
);

INVx3_ASAP7_75t_SL g3293 ( 
.A(n_2666),
.Y(n_3293)
);

INVx2_ASAP7_75t_SL g3294 ( 
.A(n_2549),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_2690),
.Y(n_3295)
);

INVx1_ASAP7_75t_SL g3296 ( 
.A(n_2360),
.Y(n_3296)
);

BUFx6f_ASAP7_75t_L g3297 ( 
.A(n_2690),
.Y(n_3297)
);

BUFx2_ASAP7_75t_L g3298 ( 
.A(n_2666),
.Y(n_3298)
);

BUFx8_ASAP7_75t_L g3299 ( 
.A(n_2591),
.Y(n_3299)
);

BUFx3_ASAP7_75t_L g3300 ( 
.A(n_2671),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_2451),
.A2(n_260),
.B1(n_256),
.B2(n_257),
.Y(n_3301)
);

BUFx2_ASAP7_75t_L g3302 ( 
.A(n_2671),
.Y(n_3302)
);

INVx2_ASAP7_75t_SL g3303 ( 
.A(n_2566),
.Y(n_3303)
);

BUFx12f_ASAP7_75t_L g3304 ( 
.A(n_2615),
.Y(n_3304)
);

INVx1_ASAP7_75t_SL g3305 ( 
.A(n_2676),
.Y(n_3305)
);

INVx1_ASAP7_75t_SL g3306 ( 
.A(n_2676),
.Y(n_3306)
);

INVx3_ASAP7_75t_SL g3307 ( 
.A(n_2518),
.Y(n_3307)
);

INVx1_ASAP7_75t_SL g3308 ( 
.A(n_2375),
.Y(n_3308)
);

BUFx4f_ASAP7_75t_SL g3309 ( 
.A(n_2733),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_2746),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_2356),
.B(n_261),
.Y(n_3311)
);

INVxp67_ASAP7_75t_SL g3312 ( 
.A(n_2518),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_2655),
.B(n_261),
.Y(n_3313)
);

INVx1_ASAP7_75t_L g3314 ( 
.A(n_2899),
.Y(n_3314)
);

CKINVDCx5p33_ASAP7_75t_R g3315 ( 
.A(n_2935),
.Y(n_3315)
);

HB1xp67_ASAP7_75t_L g3316 ( 
.A(n_3007),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2899),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2905),
.Y(n_3318)
);

CKINVDCx6p67_ASAP7_75t_R g3319 ( 
.A(n_2904),
.Y(n_3319)
);

INVx2_ASAP7_75t_L g3320 ( 
.A(n_2860),
.Y(n_3320)
);

NAND2x1p5_ASAP7_75t_L g3321 ( 
.A(n_2861),
.B(n_2637),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3276),
.B(n_2605),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3251),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3251),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_L g3325 ( 
.A(n_2864),
.Y(n_3325)
);

OAI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3241),
.A2(n_2628),
.B1(n_2748),
.B2(n_2553),
.Y(n_3326)
);

BUFx6f_ASAP7_75t_SL g3327 ( 
.A(n_2884),
.Y(n_3327)
);

INVx1_ASAP7_75t_SL g3328 ( 
.A(n_3040),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_SL g3329 ( 
.A1(n_3254),
.A2(n_2731),
.B1(n_2733),
.B2(n_2700),
.Y(n_3329)
);

INVx2_ASAP7_75t_SL g3330 ( 
.A(n_2869),
.Y(n_3330)
);

INVx2_ASAP7_75t_SL g3331 ( 
.A(n_3015),
.Y(n_3331)
);

CKINVDCx20_ASAP7_75t_R g3332 ( 
.A(n_2865),
.Y(n_3332)
);

BUFx3_ASAP7_75t_L g3333 ( 
.A(n_2960),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_3276),
.B(n_2565),
.Y(n_3334)
);

BUFx2_ASAP7_75t_L g3335 ( 
.A(n_2999),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_3034),
.A2(n_3049),
.B1(n_3081),
.B2(n_2915),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_3207),
.Y(n_3337)
);

BUFx12f_ASAP7_75t_L g3338 ( 
.A(n_2895),
.Y(n_3338)
);

AOI22xp33_ASAP7_75t_L g3339 ( 
.A1(n_3034),
.A2(n_2609),
.B1(n_2707),
.B2(n_2748),
.Y(n_3339)
);

AOI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_2903),
.A2(n_2707),
.B1(n_2785),
.B2(n_2391),
.Y(n_3340)
);

BUFx2_ASAP7_75t_L g3341 ( 
.A(n_2999),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3174),
.Y(n_3342)
);

INVx3_ASAP7_75t_L g3343 ( 
.A(n_3017),
.Y(n_3343)
);

CKINVDCx11_ASAP7_75t_R g3344 ( 
.A(n_2877),
.Y(n_3344)
);

BUFx4f_ASAP7_75t_SL g3345 ( 
.A(n_2888),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3048),
.B(n_2376),
.Y(n_3346)
);

INVx6_ASAP7_75t_L g3347 ( 
.A(n_3015),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2863),
.Y(n_3348)
);

CKINVDCx11_ASAP7_75t_R g3349 ( 
.A(n_2858),
.Y(n_3349)
);

OAI22xp5_ASAP7_75t_L g3350 ( 
.A1(n_3241),
.A2(n_2553),
.B1(n_2564),
.B2(n_2558),
.Y(n_3350)
);

BUFx4f_ASAP7_75t_SL g3351 ( 
.A(n_2901),
.Y(n_3351)
);

OAI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3293),
.A2(n_2558),
.B1(n_2564),
.B2(n_2755),
.Y(n_3352)
);

AOI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_3217),
.A2(n_2845),
.B1(n_2602),
.B2(n_2604),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3205),
.Y(n_3354)
);

OAI21xp5_ASAP7_75t_SL g3355 ( 
.A1(n_2961),
.A2(n_2660),
.B(n_2672),
.Y(n_3355)
);

INVx2_ASAP7_75t_SL g3356 ( 
.A(n_2870),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2922),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_2903),
.A2(n_2770),
.B1(n_2531),
.B2(n_2755),
.Y(n_3358)
);

BUFx3_ASAP7_75t_L g3359 ( 
.A(n_2878),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2942),
.Y(n_3360)
);

AOI22xp33_ASAP7_75t_L g3361 ( 
.A1(n_2915),
.A2(n_2770),
.B1(n_2786),
.B2(n_2752),
.Y(n_3361)
);

INVx3_ASAP7_75t_L g3362 ( 
.A(n_3017),
.Y(n_3362)
);

INVx3_ASAP7_75t_SL g3363 ( 
.A(n_2867),
.Y(n_3363)
);

OAI22xp5_ASAP7_75t_L g3364 ( 
.A1(n_3120),
.A2(n_2765),
.B1(n_2561),
.B2(n_2613),
.Y(n_3364)
);

AOI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_3002),
.A2(n_2717),
.B1(n_2685),
.B2(n_2555),
.Y(n_3365)
);

INVx3_ASAP7_75t_L g3366 ( 
.A(n_2981),
.Y(n_3366)
);

AOI22xp33_ASAP7_75t_L g3367 ( 
.A1(n_3002),
.A2(n_2786),
.B1(n_2388),
.B2(n_2772),
.Y(n_3367)
);

INVx6_ASAP7_75t_L g3368 ( 
.A(n_2859),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_2914),
.Y(n_3369)
);

HB1xp67_ASAP7_75t_L g3370 ( 
.A(n_3092),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_2871),
.Y(n_3371)
);

INVx4_ASAP7_75t_L g3372 ( 
.A(n_2875),
.Y(n_3372)
);

INVxp67_ASAP7_75t_SL g3373 ( 
.A(n_2891),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_3053),
.A2(n_2772),
.B1(n_2765),
.B2(n_2485),
.Y(n_3374)
);

OAI22xp5_ASAP7_75t_L g3375 ( 
.A1(n_3229),
.A2(n_2586),
.B1(n_2675),
.B2(n_2646),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_SL g3376 ( 
.A1(n_3181),
.A2(n_2749),
.B1(n_2649),
.B2(n_2545),
.Y(n_3376)
);

INVx1_ASAP7_75t_SL g3377 ( 
.A(n_3262),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3009),
.B(n_2393),
.Y(n_3378)
);

BUFx3_ASAP7_75t_L g3379 ( 
.A(n_2958),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_2984),
.A2(n_2430),
.B1(n_2445),
.B2(n_2424),
.Y(n_3380)
);

CKINVDCx11_ASAP7_75t_R g3381 ( 
.A(n_2928),
.Y(n_3381)
);

INVx4_ASAP7_75t_L g3382 ( 
.A(n_2875),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2914),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_2984),
.A2(n_2698),
.B1(n_2735),
.B2(n_2422),
.Y(n_3384)
);

AOI22xp33_ASAP7_75t_L g3385 ( 
.A1(n_3239),
.A2(n_2698),
.B1(n_2377),
.B2(n_2528),
.Y(n_3385)
);

CKINVDCx11_ASAP7_75t_R g3386 ( 
.A(n_2910),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2993),
.Y(n_3387)
);

BUFx6f_ASAP7_75t_L g3388 ( 
.A(n_2864),
.Y(n_3388)
);

BUFx4f_ASAP7_75t_SL g3389 ( 
.A(n_2859),
.Y(n_3389)
);

OAI21xp5_ASAP7_75t_SL g3390 ( 
.A1(n_3026),
.A2(n_2834),
.B(n_2788),
.Y(n_3390)
);

AOI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3181),
.A2(n_2622),
.B1(n_2639),
.B2(n_2674),
.Y(n_3391)
);

BUFx3_ASAP7_75t_L g3392 ( 
.A(n_3018),
.Y(n_3392)
);

CKINVDCx8_ASAP7_75t_R g3393 ( 
.A(n_2909),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_SL g3394 ( 
.A1(n_3022),
.A2(n_2649),
.B1(n_2574),
.B2(n_2527),
.Y(n_3394)
);

BUFx3_ASAP7_75t_L g3395 ( 
.A(n_2936),
.Y(n_3395)
);

INVx6_ASAP7_75t_L g3396 ( 
.A(n_2941),
.Y(n_3396)
);

OAI22xp5_ASAP7_75t_L g3397 ( 
.A1(n_3248),
.A2(n_2467),
.B1(n_2789),
.B2(n_2776),
.Y(n_3397)
);

CKINVDCx20_ASAP7_75t_R g3398 ( 
.A(n_2941),
.Y(n_3398)
);

BUFx3_ASAP7_75t_L g3399 ( 
.A(n_3013),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2905),
.Y(n_3400)
);

BUFx12f_ASAP7_75t_L g3401 ( 
.A(n_2916),
.Y(n_3401)
);

INVx1_ASAP7_75t_L g3402 ( 
.A(n_2917),
.Y(n_3402)
);

OAI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3136),
.A2(n_2825),
.B1(n_2590),
.B2(n_2361),
.Y(n_3403)
);

AOI22xp33_ASAP7_75t_L g3404 ( 
.A1(n_2904),
.A2(n_2698),
.B1(n_2535),
.B2(n_2495),
.Y(n_3404)
);

INVx2_ASAP7_75t_L g3405 ( 
.A(n_3006),
.Y(n_3405)
);

BUFx3_ASAP7_75t_L g3406 ( 
.A(n_2883),
.Y(n_3406)
);

BUFx2_ASAP7_75t_SL g3407 ( 
.A(n_2947),
.Y(n_3407)
);

CKINVDCx6p67_ASAP7_75t_R g3408 ( 
.A(n_2975),
.Y(n_3408)
);

BUFx8_ASAP7_75t_L g3409 ( 
.A(n_2940),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2917),
.Y(n_3410)
);

AND2x2_ASAP7_75t_L g3411 ( 
.A(n_2956),
.B(n_2462),
.Y(n_3411)
);

INVx6_ASAP7_75t_L g3412 ( 
.A(n_2906),
.Y(n_3412)
);

CKINVDCx11_ASAP7_75t_R g3413 ( 
.A(n_3012),
.Y(n_3413)
);

CKINVDCx20_ASAP7_75t_R g3414 ( 
.A(n_3221),
.Y(n_3414)
);

BUFx2_ASAP7_75t_SL g3415 ( 
.A(n_2947),
.Y(n_3415)
);

INVx2_ASAP7_75t_SL g3416 ( 
.A(n_2862),
.Y(n_3416)
);

INVx8_ASAP7_75t_L g3417 ( 
.A(n_2950),
.Y(n_3417)
);

BUFx2_ASAP7_75t_L g3418 ( 
.A(n_3266),
.Y(n_3418)
);

CKINVDCx8_ASAP7_75t_R g3419 ( 
.A(n_2932),
.Y(n_3419)
);

BUFx2_ASAP7_75t_L g3420 ( 
.A(n_3266),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2934),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3048),
.B(n_2866),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2866),
.B(n_2478),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3137),
.A2(n_2694),
.B1(n_2664),
.B2(n_2665),
.Y(n_3424)
);

INVx6_ASAP7_75t_L g3425 ( 
.A(n_2906),
.Y(n_3425)
);

INVx5_ASAP7_75t_SL g3426 ( 
.A(n_2950),
.Y(n_3426)
);

INVx6_ASAP7_75t_L g3427 ( 
.A(n_3177),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3044),
.Y(n_3428)
);

BUFx12f_ASAP7_75t_L g3429 ( 
.A(n_2992),
.Y(n_3429)
);

BUFx3_ASAP7_75t_L g3430 ( 
.A(n_2920),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_SL g3431 ( 
.A1(n_3024),
.A2(n_3291),
.B1(n_3309),
.B2(n_3139),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2934),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2945),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_2945),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2946),
.Y(n_3435)
);

AOI22xp33_ASAP7_75t_L g3436 ( 
.A1(n_3001),
.A2(n_2698),
.B1(n_2782),
.B2(n_2766),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_SL g3437 ( 
.A1(n_3291),
.A2(n_2771),
.B1(n_2784),
.B2(n_2501),
.Y(n_3437)
);

CKINVDCx20_ASAP7_75t_R g3438 ( 
.A(n_3146),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_3001),
.A2(n_2766),
.B1(n_2762),
.B2(n_2751),
.Y(n_3439)
);

OR2x2_ASAP7_75t_L g3440 ( 
.A(n_2874),
.B(n_2369),
.Y(n_3440)
);

OAI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_3253),
.A2(n_2762),
.B1(n_2778),
.B2(n_2777),
.Y(n_3441)
);

OAI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_2896),
.A2(n_2768),
.B1(n_2795),
.B2(n_2352),
.Y(n_3442)
);

CKINVDCx6p67_ASAP7_75t_R g3443 ( 
.A(n_2985),
.Y(n_3443)
);

AOI22xp33_ASAP7_75t_SL g3444 ( 
.A1(n_3100),
.A2(n_2771),
.B1(n_2559),
.B2(n_2562),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_2946),
.Y(n_3445)
);

CKINVDCx11_ASAP7_75t_R g3446 ( 
.A(n_2890),
.Y(n_3446)
);

BUFx4f_ASAP7_75t_SL g3447 ( 
.A(n_2965),
.Y(n_3447)
);

AOI22xp33_ASAP7_75t_L g3448 ( 
.A1(n_3031),
.A2(n_2563),
.B1(n_2512),
.B2(n_2536),
.Y(n_3448)
);

INVx4_ASAP7_75t_SL g3449 ( 
.A(n_3114),
.Y(n_3449)
);

INVx2_ASAP7_75t_L g3450 ( 
.A(n_3061),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_2949),
.Y(n_3451)
);

BUFx3_ASAP7_75t_L g3452 ( 
.A(n_3023),
.Y(n_3452)
);

NAND2x1p5_ASAP7_75t_L g3453 ( 
.A(n_2947),
.B(n_2637),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3031),
.A2(n_2732),
.B1(n_2727),
.B2(n_2712),
.Y(n_3454)
);

INVx3_ASAP7_75t_L g3455 ( 
.A(n_2990),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_L g3456 ( 
.A1(n_2919),
.A2(n_2559),
.B1(n_2562),
.B2(n_2501),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3176),
.A2(n_2806),
.B1(n_2816),
.B2(n_2803),
.Y(n_3457)
);

AOI22xp33_ASAP7_75t_L g3458 ( 
.A1(n_2919),
.A2(n_2559),
.B1(n_2562),
.B2(n_2501),
.Y(n_3458)
);

OAI22xp5_ASAP7_75t_L g3459 ( 
.A1(n_3176),
.A2(n_2819),
.B1(n_2822),
.B2(n_2818),
.Y(n_3459)
);

INVx2_ASAP7_75t_L g3460 ( 
.A(n_3079),
.Y(n_3460)
);

AOI22xp5_ASAP7_75t_L g3461 ( 
.A1(n_3137),
.A2(n_2775),
.B1(n_2559),
.B2(n_2562),
.Y(n_3461)
);

INVx6_ASAP7_75t_L g3462 ( 
.A(n_3177),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3105),
.Y(n_3463)
);

BUFx4_ASAP7_75t_SL g3464 ( 
.A(n_2868),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2949),
.Y(n_3465)
);

NAND2x1p5_ASAP7_75t_L g3466 ( 
.A(n_3037),
.B(n_2637),
.Y(n_3466)
);

BUFx10_ASAP7_75t_L g3467 ( 
.A(n_3057),
.Y(n_3467)
);

BUFx3_ASAP7_75t_L g3468 ( 
.A(n_3023),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_2973),
.A2(n_2570),
.B1(n_2501),
.B2(n_2581),
.Y(n_3469)
);

AOI22xp33_ASAP7_75t_L g3470 ( 
.A1(n_2973),
.A2(n_2570),
.B1(n_2753),
.B2(n_2476),
.Y(n_3470)
);

OAI21xp5_ASAP7_75t_SL g3471 ( 
.A1(n_3071),
.A2(n_2630),
.B(n_2738),
.Y(n_3471)
);

OR2x2_ASAP7_75t_L g3472 ( 
.A(n_2967),
.B(n_2372),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3112),
.Y(n_3473)
);

BUFx6f_ASAP7_75t_SL g3474 ( 
.A(n_3057),
.Y(n_3474)
);

BUFx2_ASAP7_75t_L g3475 ( 
.A(n_3260),
.Y(n_3475)
);

CKINVDCx20_ASAP7_75t_R g3476 ( 
.A(n_3103),
.Y(n_3476)
);

OAI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3111),
.A2(n_2843),
.B1(n_2849),
.B2(n_2832),
.Y(n_3477)
);

INVx1_ASAP7_75t_SL g3478 ( 
.A(n_3273),
.Y(n_3478)
);

INVx6_ASAP7_75t_L g3479 ( 
.A(n_3299),
.Y(n_3479)
);

BUFx3_ASAP7_75t_L g3480 ( 
.A(n_3274),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_2965),
.A2(n_3299),
.B1(n_3290),
.B2(n_3269),
.Y(n_3481)
);

AOI22xp33_ASAP7_75t_SL g3482 ( 
.A1(n_3150),
.A2(n_3158),
.B1(n_3004),
.B2(n_3019),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_2873),
.B(n_2689),
.Y(n_3483)
);

INVx6_ASAP7_75t_L g3484 ( 
.A(n_3066),
.Y(n_3484)
);

CKINVDCx16_ASAP7_75t_R g3485 ( 
.A(n_3110),
.Y(n_3485)
);

INVx3_ASAP7_75t_L g3486 ( 
.A(n_3037),
.Y(n_3486)
);

INVxp67_ASAP7_75t_SL g3487 ( 
.A(n_3076),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_SL g3488 ( 
.A1(n_2997),
.A2(n_2771),
.B1(n_2570),
.B2(n_2738),
.Y(n_3488)
);

OAI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_3111),
.A2(n_2856),
.B1(n_2756),
.B2(n_2744),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_2952),
.Y(n_3490)
);

OAI22xp5_ASAP7_75t_L g3491 ( 
.A1(n_3307),
.A2(n_2517),
.B1(n_2514),
.B2(n_2759),
.Y(n_3491)
);

BUFx4f_ASAP7_75t_SL g3492 ( 
.A(n_3247),
.Y(n_3492)
);

AOI22xp33_ASAP7_75t_SL g3493 ( 
.A1(n_3267),
.A2(n_2771),
.B1(n_2570),
.B2(n_2363),
.Y(n_3493)
);

INVx2_ASAP7_75t_SL g3494 ( 
.A(n_2988),
.Y(n_3494)
);

AOI22xp33_ASAP7_75t_L g3495 ( 
.A1(n_3290),
.A2(n_2455),
.B1(n_2480),
.B2(n_2654),
.Y(n_3495)
);

OAI22xp33_ASAP7_75t_SL g3496 ( 
.A1(n_3256),
.A2(n_2728),
.B1(n_2509),
.B2(n_2835),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3090),
.B(n_2619),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2952),
.Y(n_3498)
);

BUFx2_ASAP7_75t_SL g3499 ( 
.A(n_2889),
.Y(n_3499)
);

CKINVDCx6p67_ASAP7_75t_R g3500 ( 
.A(n_2948),
.Y(n_3500)
);

CKINVDCx5p33_ASAP7_75t_R g3501 ( 
.A(n_2918),
.Y(n_3501)
);

BUFx3_ASAP7_75t_L g3502 ( 
.A(n_3027),
.Y(n_3502)
);

BUFx8_ASAP7_75t_SL g3503 ( 
.A(n_3125),
.Y(n_3503)
);

AOI22xp33_ASAP7_75t_L g3504 ( 
.A1(n_3072),
.A2(n_2463),
.B1(n_2473),
.B2(n_2584),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_L g3505 ( 
.A1(n_3188),
.A2(n_2594),
.B1(n_2598),
.B2(n_2587),
.Y(n_3505)
);

INVx2_ASAP7_75t_SL g3506 ( 
.A(n_2953),
.Y(n_3506)
);

AOI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3202),
.A2(n_2616),
.B1(n_2652),
.B2(n_2635),
.Y(n_3507)
);

AND2x2_ASAP7_75t_L g3508 ( 
.A(n_3078),
.B(n_2647),
.Y(n_3508)
);

INVx4_ASAP7_75t_L g3509 ( 
.A(n_3064),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2963),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_2882),
.B(n_2661),
.Y(n_3511)
);

AOI22xp33_ASAP7_75t_SL g3512 ( 
.A1(n_3114),
.A2(n_2363),
.B1(n_2506),
.B2(n_2627),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3151),
.Y(n_3513)
);

INVx1_ASAP7_75t_SL g3514 ( 
.A(n_3035),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3164),
.Y(n_3515)
);

BUFx2_ASAP7_75t_L g3516 ( 
.A(n_3260),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3168),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3168),
.Y(n_3518)
);

INVx6_ASAP7_75t_L g3519 ( 
.A(n_3304),
.Y(n_3519)
);

CKINVDCx5p33_ASAP7_75t_R g3520 ( 
.A(n_2930),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_2963),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2873),
.B(n_2431),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_2964),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3085),
.A2(n_2697),
.B1(n_2759),
.B2(n_2592),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3128),
.A2(n_2502),
.B1(n_2500),
.B2(n_2631),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3252),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_2887),
.Y(n_3527)
);

BUFx2_ASAP7_75t_L g3528 ( 
.A(n_2976),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_2964),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_2943),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2966),
.Y(n_3531)
);

INVx5_ASAP7_75t_L g3532 ( 
.A(n_3114),
.Y(n_3532)
);

OAI22xp33_ASAP7_75t_L g3533 ( 
.A1(n_3075),
.A2(n_2342),
.B1(n_2692),
.B2(n_2544),
.Y(n_3533)
);

AOI22xp33_ASAP7_75t_L g3534 ( 
.A1(n_3075),
.A2(n_2670),
.B1(n_2669),
.B2(n_2761),
.Y(n_3534)
);

AOI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3249),
.A2(n_2572),
.B1(n_2573),
.B2(n_2537),
.Y(n_3535)
);

INVx1_ASAP7_75t_SL g3536 ( 
.A(n_2957),
.Y(n_3536)
);

BUFx12f_ASAP7_75t_L g3537 ( 
.A(n_2927),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_2887),
.Y(n_3538)
);

CKINVDCx11_ASAP7_75t_R g3539 ( 
.A(n_3083),
.Y(n_3539)
);

BUFx3_ASAP7_75t_L g3540 ( 
.A(n_2953),
.Y(n_3540)
);

BUFx6f_ASAP7_75t_L g3541 ( 
.A(n_2864),
.Y(n_3541)
);

BUFx2_ASAP7_75t_L g3542 ( 
.A(n_3039),
.Y(n_3542)
);

INVx3_ASAP7_75t_L g3543 ( 
.A(n_3064),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_2966),
.Y(n_3544)
);

AND2x2_ASAP7_75t_L g3545 ( 
.A(n_3192),
.B(n_2568),
.Y(n_3545)
);

AOI22xp33_ASAP7_75t_SL g3546 ( 
.A1(n_3114),
.A2(n_2506),
.B1(n_2419),
.B2(n_2529),
.Y(n_3546)
);

AOI22xp33_ASAP7_75t_SL g3547 ( 
.A1(n_3235),
.A2(n_2506),
.B1(n_2781),
.B2(n_2722),
.Y(n_3547)
);

INVx1_ASAP7_75t_SL g3548 ( 
.A(n_2872),
.Y(n_3548)
);

CKINVDCx16_ASAP7_75t_R g3549 ( 
.A(n_3052),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2974),
.Y(n_3550)
);

BUFx12f_ASAP7_75t_L g3551 ( 
.A(n_2977),
.Y(n_3551)
);

AOI22xp33_ASAP7_75t_L g3552 ( 
.A1(n_2886),
.A2(n_2761),
.B1(n_2687),
.B2(n_2703),
.Y(n_3552)
);

BUFx8_ASAP7_75t_L g3553 ( 
.A(n_3196),
.Y(n_3553)
);

BUFx3_ASAP7_75t_L g3554 ( 
.A(n_3028),
.Y(n_3554)
);

INVx1_ASAP7_75t_L g3555 ( 
.A(n_2974),
.Y(n_3555)
);

AOI22xp33_ASAP7_75t_L g3556 ( 
.A1(n_2886),
.A2(n_2696),
.B1(n_2686),
.B2(n_2680),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_L g3557 ( 
.A1(n_3080),
.A2(n_2425),
.B1(n_2423),
.B2(n_2551),
.Y(n_3557)
);

BUFx8_ASAP7_75t_L g3558 ( 
.A(n_3199),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_2983),
.Y(n_3559)
);

INVx3_ASAP7_75t_SL g3560 ( 
.A(n_3263),
.Y(n_3560)
);

BUFx6f_ASAP7_75t_L g3561 ( 
.A(n_2885),
.Y(n_3561)
);

BUFx3_ASAP7_75t_L g3562 ( 
.A(n_3030),
.Y(n_3562)
);

INVx2_ASAP7_75t_SL g3563 ( 
.A(n_3279),
.Y(n_3563)
);

CKINVDCx6p67_ASAP7_75t_R g3564 ( 
.A(n_3129),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_2983),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_2998),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_2998),
.Y(n_3567)
);

AOI22xp5_ASAP7_75t_L g3568 ( 
.A1(n_3180),
.A2(n_2398),
.B1(n_2407),
.B2(n_2406),
.Y(n_3568)
);

CKINVDCx11_ASAP7_75t_R g3569 ( 
.A(n_3131),
.Y(n_3569)
);

CKINVDCx5p33_ASAP7_75t_R g3570 ( 
.A(n_3195),
.Y(n_3570)
);

BUFx10_ASAP7_75t_L g3571 ( 
.A(n_3121),
.Y(n_3571)
);

CKINVDCx11_ASAP7_75t_R g3572 ( 
.A(n_3143),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3180),
.A2(n_2490),
.B1(n_2724),
.B2(n_2715),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3003),
.Y(n_3574)
);

CKINVDCx11_ASAP7_75t_R g3575 ( 
.A(n_3147),
.Y(n_3575)
);

OAI22xp5_ASAP7_75t_L g3576 ( 
.A1(n_3312),
.A2(n_2722),
.B1(n_2758),
.B2(n_2679),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3003),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3011),
.Y(n_3578)
);

AOI22xp33_ASAP7_75t_L g3579 ( 
.A1(n_2996),
.A2(n_2790),
.B1(n_2758),
.B2(n_2679),
.Y(n_3579)
);

BUFx3_ASAP7_75t_L g3580 ( 
.A(n_3197),
.Y(n_3580)
);

BUFx10_ASAP7_75t_L g3581 ( 
.A(n_3121),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3011),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3021),
.Y(n_3583)
);

CKINVDCx16_ASAP7_75t_R g3584 ( 
.A(n_3054),
.Y(n_3584)
);

OAI22xp33_ASAP7_75t_L g3585 ( 
.A1(n_3255),
.A2(n_2728),
.B1(n_2705),
.B2(n_2713),
.Y(n_3585)
);

BUFx8_ASAP7_75t_L g3586 ( 
.A(n_3036),
.Y(n_3586)
);

AOI22xp33_ASAP7_75t_L g3587 ( 
.A1(n_3165),
.A2(n_2781),
.B1(n_2610),
.B2(n_2583),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_2893),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_2893),
.Y(n_3589)
);

HB1xp67_ASAP7_75t_L g3590 ( 
.A(n_3058),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_2894),
.Y(n_3591)
);

AOI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_3308),
.A2(n_2739),
.B1(n_2740),
.B2(n_2706),
.Y(n_3592)
);

AOI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3298),
.A2(n_2682),
.B1(n_2757),
.B2(n_2745),
.Y(n_3593)
);

INVx4_ASAP7_75t_L g3594 ( 
.A(n_3074),
.Y(n_3594)
);

BUFx2_ASAP7_75t_SL g3595 ( 
.A(n_3204),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3186),
.B(n_264),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_SL g3597 ( 
.A1(n_3302),
.A2(n_2506),
.B1(n_2780),
.B2(n_2773),
.Y(n_3597)
);

BUFx12f_ASAP7_75t_L g3598 ( 
.A(n_3029),
.Y(n_3598)
);

CKINVDCx6p67_ASAP7_75t_R g3599 ( 
.A(n_3060),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_2894),
.Y(n_3600)
);

BUFx12f_ASAP7_75t_L g3601 ( 
.A(n_3029),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3021),
.Y(n_3602)
);

INVx1_ASAP7_75t_SL g3603 ( 
.A(n_2876),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3051),
.Y(n_3604)
);

BUFx12f_ASAP7_75t_L g3605 ( 
.A(n_2929),
.Y(n_3605)
);

BUFx4f_ASAP7_75t_L g3606 ( 
.A(n_3032),
.Y(n_3606)
);

INVx4_ASAP7_75t_SL g3607 ( 
.A(n_3264),
.Y(n_3607)
);

BUFx6f_ASAP7_75t_L g3608 ( 
.A(n_2885),
.Y(n_3608)
);

OAI22xp33_ASAP7_75t_L g3609 ( 
.A1(n_3280),
.A2(n_2764),
.B1(n_2835),
.B2(n_2509),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3051),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3305),
.A2(n_2607),
.B1(n_2780),
.B2(n_2773),
.Y(n_3611)
);

AOI22xp33_ASAP7_75t_SL g3612 ( 
.A1(n_3282),
.A2(n_2780),
.B1(n_2783),
.B2(n_2773),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3062),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3306),
.A2(n_2783),
.B1(n_2614),
.B2(n_2426),
.Y(n_3614)
);

BUFx6f_ASAP7_75t_L g3615 ( 
.A(n_2885),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3268),
.A2(n_2783),
.B1(n_2791),
.B2(n_2763),
.Y(n_3616)
);

CKINVDCx11_ASAP7_75t_R g3617 ( 
.A(n_2955),
.Y(n_3617)
);

INVx8_ASAP7_75t_L g3618 ( 
.A(n_3055),
.Y(n_3618)
);

AOI22xp33_ASAP7_75t_L g3619 ( 
.A1(n_3097),
.A2(n_2791),
.B1(n_2763),
.B2(n_2426),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3062),
.Y(n_3620)
);

AOI22xp33_ASAP7_75t_L g3621 ( 
.A1(n_3116),
.A2(n_2763),
.B1(n_2449),
.B2(n_2482),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3170),
.Y(n_3622)
);

CKINVDCx14_ASAP7_75t_R g3623 ( 
.A(n_2880),
.Y(n_3623)
);

OAI22xp33_ASAP7_75t_L g3624 ( 
.A1(n_3284),
.A2(n_2737),
.B1(n_2794),
.B2(n_2787),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3148),
.A2(n_3166),
.B1(n_3138),
.B2(n_3228),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3063),
.Y(n_3626)
);

OAI22xp33_ASAP7_75t_L g3627 ( 
.A1(n_3300),
.A2(n_2737),
.B1(n_2688),
.B2(n_2449),
.Y(n_3627)
);

AOI22xp33_ASAP7_75t_SL g3628 ( 
.A1(n_3243),
.A2(n_2482),
.B1(n_2340),
.B2(n_2667),
.Y(n_3628)
);

OAI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_3086),
.A2(n_2737),
.B1(n_2688),
.B2(n_2340),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3264),
.A2(n_2667),
.B1(n_2576),
.B2(n_2632),
.Y(n_3630)
);

CKINVDCx5p33_ASAP7_75t_R g3631 ( 
.A(n_3216),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3063),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3065),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3065),
.Y(n_3634)
);

INVxp67_ASAP7_75t_L g3635 ( 
.A(n_2900),
.Y(n_3635)
);

CKINVDCx11_ASAP7_75t_R g3636 ( 
.A(n_2923),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3261),
.B(n_2571),
.Y(n_3637)
);

AOI22xp33_ASAP7_75t_L g3638 ( 
.A1(n_3272),
.A2(n_3099),
.B1(n_3141),
.B2(n_3038),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3067),
.Y(n_3639)
);

OAI22xp33_ASAP7_75t_L g3640 ( 
.A1(n_2908),
.A2(n_2571),
.B1(n_2632),
.B2(n_2576),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3067),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3170),
.Y(n_3642)
);

INVx2_ASAP7_75t_L g3643 ( 
.A(n_3182),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3272),
.A2(n_2667),
.B1(n_2656),
.B2(n_2793),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3093),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3261),
.B(n_2656),
.Y(n_3646)
);

AOI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_3296),
.A2(n_2720),
.B1(n_2723),
.B2(n_2711),
.Y(n_3647)
);

INVx8_ASAP7_75t_L g3648 ( 
.A(n_3055),
.Y(n_3648)
);

AOI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3047),
.A2(n_2720),
.B1(n_2723),
.B2(n_2651),
.Y(n_3649)
);

AOI22xp5_ASAP7_75t_L g3650 ( 
.A1(n_3113),
.A2(n_2742),
.B1(n_2711),
.B2(n_2691),
.Y(n_3650)
);

AOI22xp33_ASAP7_75t_L g3651 ( 
.A1(n_3245),
.A2(n_2651),
.B1(n_2702),
.B2(n_2691),
.Y(n_3651)
);

BUFx2_ASAP7_75t_L g3652 ( 
.A(n_3250),
.Y(n_3652)
);

BUFx3_ASAP7_75t_L g3653 ( 
.A(n_3149),
.Y(n_3653)
);

BUFx2_ASAP7_75t_L g3654 ( 
.A(n_3160),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3171),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_2912),
.Y(n_3656)
);

INVx6_ASAP7_75t_L g3657 ( 
.A(n_3173),
.Y(n_3657)
);

OAI22xp33_ASAP7_75t_L g3658 ( 
.A1(n_2987),
.A2(n_2690),
.B1(n_2699),
.B2(n_2541),
.Y(n_3658)
);

INVx2_ASAP7_75t_L g3659 ( 
.A(n_3182),
.Y(n_3659)
);

INVx3_ASAP7_75t_L g3660 ( 
.A(n_3074),
.Y(n_3660)
);

INVxp67_ASAP7_75t_SL g3661 ( 
.A(n_2926),
.Y(n_3661)
);

INVx4_ASAP7_75t_SL g3662 ( 
.A(n_2994),
.Y(n_3662)
);

BUFx12f_ASAP7_75t_L g3663 ( 
.A(n_3042),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3270),
.B(n_2479),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_2912),
.Y(n_3665)
);

BUFx12f_ASAP7_75t_L g3666 ( 
.A(n_3185),
.Y(n_3666)
);

AOI22xp33_ASAP7_75t_SL g3667 ( 
.A1(n_3189),
.A2(n_2534),
.B1(n_2479),
.B2(n_2651),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_2913),
.Y(n_3668)
);

CKINVDCx11_ASAP7_75t_R g3669 ( 
.A(n_2944),
.Y(n_3669)
);

OAI22xp5_ASAP7_75t_L g3670 ( 
.A1(n_3056),
.A2(n_2699),
.B1(n_2521),
.B2(n_2552),
.Y(n_3670)
);

INVx2_ASAP7_75t_SL g3671 ( 
.A(n_3175),
.Y(n_3671)
);

BUFx6f_ASAP7_75t_L g3672 ( 
.A(n_2911),
.Y(n_3672)
);

INVx2_ASAP7_75t_L g3673 ( 
.A(n_3203),
.Y(n_3673)
);

INVx6_ASAP7_75t_L g3674 ( 
.A(n_3187),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3118),
.B(n_264),
.Y(n_3675)
);

INVx1_ASAP7_75t_L g3676 ( 
.A(n_2913),
.Y(n_3676)
);

INVx4_ASAP7_75t_L g3677 ( 
.A(n_3055),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3270),
.B(n_2534),
.Y(n_3678)
);

BUFx4f_ASAP7_75t_L g3679 ( 
.A(n_3194),
.Y(n_3679)
);

OAI22xp5_ASAP7_75t_L g3680 ( 
.A1(n_3167),
.A2(n_2699),
.B1(n_2521),
.B2(n_2552),
.Y(n_3680)
);

OAI22xp5_ASAP7_75t_L g3681 ( 
.A1(n_3201),
.A2(n_2515),
.B1(n_2742),
.B2(n_2708),
.Y(n_3681)
);

CKINVDCx5p33_ASAP7_75t_R g3682 ( 
.A(n_3130),
.Y(n_3682)
);

BUFx12f_ASAP7_75t_L g3683 ( 
.A(n_2954),
.Y(n_3683)
);

INVx4_ASAP7_75t_L g3684 ( 
.A(n_3068),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3285),
.Y(n_3685)
);

INVx5_ASAP7_75t_L g3686 ( 
.A(n_3068),
.Y(n_3686)
);

BUFx6f_ASAP7_75t_L g3687 ( 
.A(n_2911),
.Y(n_3687)
);

BUFx8_ASAP7_75t_L g3688 ( 
.A(n_2978),
.Y(n_3688)
);

OAI22xp33_ASAP7_75t_L g3689 ( 
.A1(n_3127),
.A2(n_2515),
.B1(n_2721),
.B2(n_2708),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_SL g3690 ( 
.A1(n_3144),
.A2(n_2721),
.B1(n_2702),
.B2(n_267),
.Y(n_3690)
);

BUFx6f_ASAP7_75t_L g3691 ( 
.A(n_2911),
.Y(n_3691)
);

BUFx8_ASAP7_75t_SL g3692 ( 
.A(n_2979),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_SL g3693 ( 
.A1(n_3152),
.A2(n_2721),
.B1(n_267),
.B2(n_265),
.Y(n_3693)
);

BUFx3_ASAP7_75t_L g3694 ( 
.A(n_2951),
.Y(n_3694)
);

BUFx2_ASAP7_75t_L g3695 ( 
.A(n_3088),
.Y(n_3695)
);

BUFx2_ASAP7_75t_L g3696 ( 
.A(n_3190),
.Y(n_3696)
);

OAI22xp5_ASAP7_75t_SL g3697 ( 
.A1(n_2898),
.A2(n_270),
.B1(n_266),
.B2(n_268),
.Y(n_3697)
);

BUFx6f_ASAP7_75t_L g3698 ( 
.A(n_3618),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3474),
.A2(n_2937),
.B1(n_3041),
.B2(n_3096),
.Y(n_3699)
);

BUFx6f_ASAP7_75t_L g3700 ( 
.A(n_3618),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3357),
.Y(n_3701)
);

INVx4_ASAP7_75t_L g3702 ( 
.A(n_3686),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3474),
.A2(n_3210),
.B1(n_3240),
.B2(n_3222),
.Y(n_3703)
);

OAI222xp33_ASAP7_75t_L g3704 ( 
.A1(n_3326),
.A2(n_3288),
.B1(n_3281),
.B2(n_3206),
.C1(n_3313),
.C2(n_3016),
.Y(n_3704)
);

AOI22xp33_ASAP7_75t_SL g3705 ( 
.A1(n_3417),
.A2(n_3350),
.B1(n_3426),
.B2(n_3532),
.Y(n_3705)
);

OAI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_3456),
.A2(n_3458),
.B1(n_3461),
.B2(n_3367),
.Y(n_3706)
);

AOI22xp33_ASAP7_75t_SL g3707 ( 
.A1(n_3417),
.A2(n_2881),
.B1(n_2907),
.B2(n_2892),
.Y(n_3707)
);

AOI22xp33_ASAP7_75t_L g3708 ( 
.A1(n_3439),
.A2(n_3163),
.B1(n_3119),
.B2(n_3159),
.Y(n_3708)
);

AOI222xp33_ASAP7_75t_L g3709 ( 
.A1(n_3697),
.A2(n_3134),
.B1(n_3109),
.B2(n_3020),
.C1(n_3178),
.C2(n_3157),
.Y(n_3709)
);

BUFx12f_ASAP7_75t_L g3710 ( 
.A(n_3386),
.Y(n_3710)
);

AOI222xp33_ASAP7_75t_L g3711 ( 
.A1(n_3426),
.A2(n_3478),
.B1(n_3389),
.B2(n_3606),
.C1(n_3467),
.C2(n_3447),
.Y(n_3711)
);

HB1xp67_ASAP7_75t_L g3712 ( 
.A(n_3695),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3322),
.B(n_3093),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3596),
.B(n_3154),
.Y(n_3714)
);

BUFx12f_ASAP7_75t_L g3715 ( 
.A(n_3349),
.Y(n_3715)
);

AOI22xp33_ASAP7_75t_L g3716 ( 
.A1(n_3329),
.A2(n_3403),
.B1(n_3441),
.B2(n_3679),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3360),
.Y(n_3717)
);

OAI21xp5_ASAP7_75t_SL g3718 ( 
.A1(n_3355),
.A2(n_3301),
.B(n_3050),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_SL g3719 ( 
.A1(n_3532),
.A2(n_3352),
.B1(n_3467),
.B2(n_3571),
.Y(n_3719)
);

AOI222xp33_ASAP7_75t_L g3720 ( 
.A1(n_3606),
.A2(n_3077),
.B1(n_3145),
.B2(n_3278),
.C1(n_3169),
.C2(n_3172),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3337),
.B(n_3094),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3342),
.Y(n_3722)
);

AOI22xp33_ASAP7_75t_SL g3723 ( 
.A1(n_3532),
.A2(n_2881),
.B1(n_2907),
.B2(n_2892),
.Y(n_3723)
);

OAI222xp33_ASAP7_75t_L g3724 ( 
.A1(n_3376),
.A2(n_3287),
.B1(n_3285),
.B2(n_3271),
.C1(n_3162),
.C2(n_2921),
.Y(n_3724)
);

AOI22xp33_ASAP7_75t_L g3725 ( 
.A1(n_3679),
.A2(n_3287),
.B1(n_2980),
.B2(n_2972),
.Y(n_3725)
);

INVx3_ASAP7_75t_L g3726 ( 
.A(n_3509),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_3444),
.A2(n_2972),
.B1(n_2980),
.B2(n_2962),
.Y(n_3727)
);

OAI22xp5_ASAP7_75t_L g3728 ( 
.A1(n_3469),
.A2(n_2897),
.B1(n_2879),
.B2(n_3311),
.Y(n_3728)
);

OAI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_3437),
.A2(n_2879),
.B1(n_2971),
.B2(n_2902),
.Y(n_3729)
);

OR2x2_ASAP7_75t_L g3730 ( 
.A(n_3316),
.B(n_3203),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_L g3731 ( 
.A1(n_3690),
.A2(n_2986),
.B1(n_3008),
.B2(n_2982),
.Y(n_3731)
);

OAI22xp5_ASAP7_75t_L g3732 ( 
.A1(n_3339),
.A2(n_3087),
.B1(n_3010),
.B2(n_3230),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3354),
.B(n_3094),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3323),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3693),
.A2(n_3122),
.B1(n_3132),
.B2(n_3107),
.Y(n_3735)
);

AOI22xp33_ASAP7_75t_L g3736 ( 
.A1(n_3340),
.A2(n_3122),
.B1(n_3132),
.B2(n_3107),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_L g3737 ( 
.A1(n_3378),
.A2(n_3142),
.B1(n_3133),
.B2(n_3200),
.Y(n_3737)
);

AOI22xp33_ASAP7_75t_SL g3738 ( 
.A1(n_3571),
.A2(n_3225),
.B1(n_3014),
.B2(n_3142),
.Y(n_3738)
);

INVx5_ASAP7_75t_SL g3739 ( 
.A(n_3319),
.Y(n_3739)
);

INVxp67_ASAP7_75t_L g3740 ( 
.A(n_3370),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3324),
.Y(n_3741)
);

BUFx2_ASAP7_75t_L g3742 ( 
.A(n_3487),
.Y(n_3742)
);

BUFx3_ASAP7_75t_L g3743 ( 
.A(n_3492),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3604),
.Y(n_3744)
);

OAI21xp33_ASAP7_75t_L g3745 ( 
.A1(n_3394),
.A2(n_3244),
.B(n_3242),
.Y(n_3745)
);

AOI22xp33_ASAP7_75t_L g3746 ( 
.A1(n_3491),
.A2(n_3133),
.B1(n_3303),
.B2(n_3294),
.Y(n_3746)
);

AOI22xp33_ASAP7_75t_L g3747 ( 
.A1(n_3411),
.A2(n_3098),
.B1(n_3101),
.B2(n_3073),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3610),
.Y(n_3748)
);

BUFx3_ASAP7_75t_L g3749 ( 
.A(n_3395),
.Y(n_3749)
);

AND2x2_ASAP7_75t_L g3750 ( 
.A(n_3675),
.B(n_3242),
.Y(n_3750)
);

OAI22xp33_ASAP7_75t_L g3751 ( 
.A1(n_3365),
.A2(n_3014),
.B1(n_3193),
.B2(n_3244),
.Y(n_3751)
);

OAI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3373),
.A2(n_3213),
.B1(n_3215),
.B2(n_3211),
.Y(n_3752)
);

AND2x2_ASAP7_75t_L g3753 ( 
.A(n_3497),
.B(n_2924),
.Y(n_3753)
);

INVx5_ASAP7_75t_SL g3754 ( 
.A(n_3500),
.Y(n_3754)
);

AOI22xp33_ASAP7_75t_L g3755 ( 
.A1(n_3579),
.A2(n_3310),
.B1(n_3283),
.B2(n_3213),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3622),
.Y(n_3756)
);

AOI22xp33_ASAP7_75t_L g3757 ( 
.A1(n_3556),
.A2(n_3511),
.B1(n_3457),
.B2(n_3459),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3334),
.B(n_3211),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3642),
.Y(n_3759)
);

AOI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3375),
.A2(n_3218),
.B1(n_3226),
.B2(n_3215),
.Y(n_3760)
);

OAI21xp5_ASAP7_75t_SL g3761 ( 
.A1(n_3482),
.A2(n_3431),
.B(n_3493),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_SL g3762 ( 
.A1(n_3581),
.A2(n_3225),
.B1(n_3089),
.B2(n_3123),
.Y(n_3762)
);

AOI22xp33_ASAP7_75t_L g3763 ( 
.A1(n_3508),
.A2(n_3226),
.B1(n_3231),
.B2(n_3218),
.Y(n_3763)
);

AND2x2_ASAP7_75t_L g3764 ( 
.A(n_3399),
.B(n_2925),
.Y(n_3764)
);

OAI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_3374),
.A2(n_3231),
.B1(n_3115),
.B2(n_3123),
.Y(n_3765)
);

CKINVDCx20_ASAP7_75t_R g3766 ( 
.A(n_3398),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3509),
.Y(n_3767)
);

BUFx4f_ASAP7_75t_SL g3768 ( 
.A(n_3338),
.Y(n_3768)
);

AOI22xp33_ASAP7_75t_SL g3769 ( 
.A1(n_3581),
.A2(n_3225),
.B1(n_3089),
.B2(n_3198),
.Y(n_3769)
);

OR2x2_ASAP7_75t_L g3770 ( 
.A(n_3590),
.B(n_2931),
.Y(n_3770)
);

OAI21xp33_ASAP7_75t_L g3771 ( 
.A1(n_3353),
.A2(n_2969),
.B(n_2968),
.Y(n_3771)
);

CKINVDCx5p33_ASAP7_75t_R g3772 ( 
.A(n_3503),
.Y(n_3772)
);

AOI22xp33_ASAP7_75t_L g3773 ( 
.A1(n_3552),
.A2(n_2989),
.B1(n_2991),
.B2(n_2970),
.Y(n_3773)
);

CKINVDCx5p33_ASAP7_75t_R g3774 ( 
.A(n_3315),
.Y(n_3774)
);

OAI222xp33_ASAP7_75t_L g3775 ( 
.A1(n_3488),
.A2(n_3193),
.B1(n_3198),
.B2(n_3115),
.C1(n_3135),
.C2(n_3104),
.Y(n_3775)
);

OAI21xp5_ASAP7_75t_SL g3776 ( 
.A1(n_3336),
.A2(n_3220),
.B(n_3208),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3625),
.A2(n_3234),
.B1(n_3237),
.B2(n_3232),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3385),
.A2(n_3246),
.B1(n_3069),
.B2(n_3124),
.Y(n_3778)
);

AOI22xp33_ASAP7_75t_L g3779 ( 
.A1(n_3364),
.A2(n_3117),
.B1(n_3126),
.B2(n_3225),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3534),
.A2(n_3225),
.B1(n_3179),
.B2(n_3104),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3643),
.Y(n_3781)
);

OAI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_3485),
.A2(n_3257),
.B1(n_3155),
.B2(n_3091),
.Y(n_3782)
);

BUFx4f_ASAP7_75t_SL g3783 ( 
.A(n_3332),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3613),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_3526),
.B(n_266),
.Y(n_3785)
);

AOI22xp33_ASAP7_75t_L g3786 ( 
.A1(n_3504),
.A2(n_3212),
.B1(n_3236),
.B2(n_3209),
.Y(n_3786)
);

OAI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3380),
.A2(n_3091),
.B1(n_3106),
.B2(n_3068),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_3422),
.B(n_3091),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3659),
.Y(n_3789)
);

BUFx4f_ASAP7_75t_SL g3790 ( 
.A(n_3401),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3448),
.A2(n_3212),
.B1(n_3236),
.B2(n_3209),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3549),
.B(n_271),
.Y(n_3792)
);

OAI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3358),
.A2(n_3108),
.B1(n_3140),
.B2(n_3106),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3673),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3584),
.B(n_271),
.Y(n_3795)
);

AOI22xp33_ASAP7_75t_L g3796 ( 
.A1(n_3495),
.A2(n_3259),
.B1(n_3258),
.B2(n_3108),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3620),
.B(n_3106),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3626),
.B(n_3632),
.Y(n_3798)
);

AOI22xp33_ASAP7_75t_L g3799 ( 
.A1(n_3623),
.A2(n_3259),
.B1(n_3258),
.B2(n_3140),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3573),
.A2(n_3140),
.B1(n_3153),
.B2(n_3108),
.Y(n_3800)
);

INVx4_ASAP7_75t_L g3801 ( 
.A(n_3686),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3436),
.A2(n_3155),
.B1(n_3161),
.B2(n_3153),
.Y(n_3802)
);

CKINVDCx6p67_ASAP7_75t_R g3803 ( 
.A(n_3363),
.Y(n_3803)
);

AOI22xp33_ASAP7_75t_L g3804 ( 
.A1(n_3533),
.A2(n_3155),
.B1(n_3161),
.B2(n_3153),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_SL g3805 ( 
.A1(n_3407),
.A2(n_3184),
.B1(n_3238),
.B2(n_3161),
.Y(n_3805)
);

NAND2x1p5_ASAP7_75t_L g3806 ( 
.A(n_3686),
.B(n_3184),
.Y(n_3806)
);

INVx2_ASAP7_75t_SL g3807 ( 
.A(n_3484),
.Y(n_3807)
);

OAI21xp5_ASAP7_75t_SL g3808 ( 
.A1(n_3481),
.A2(n_3341),
.B(n_3335),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_3517),
.B(n_272),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3633),
.B(n_3184),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3634),
.B(n_3238),
.Y(n_3811)
);

OAI22xp5_ASAP7_75t_L g3812 ( 
.A1(n_3361),
.A2(n_3257),
.B1(n_3265),
.B2(n_3238),
.Y(n_3812)
);

INVx1_ASAP7_75t_L g3813 ( 
.A(n_3639),
.Y(n_3813)
);

OAI21xp5_ASAP7_75t_SL g3814 ( 
.A1(n_3390),
.A2(n_2938),
.B(n_2933),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3384),
.A2(n_3265),
.B1(n_3277),
.B2(n_3257),
.Y(n_3815)
);

BUFx2_ASAP7_75t_L g3816 ( 
.A(n_3607),
.Y(n_3816)
);

OA222x2_ASAP7_75t_L g3817 ( 
.A1(n_3664),
.A2(n_3277),
.B1(n_3265),
.B2(n_274),
.C1(n_276),
.C2(n_272),
.Y(n_3817)
);

OAI22xp5_ASAP7_75t_SL g3818 ( 
.A1(n_3414),
.A2(n_3277),
.B1(n_2938),
.B2(n_2939),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3641),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3470),
.A2(n_3297),
.B1(n_3295),
.B2(n_3191),
.Y(n_3820)
);

AOI22xp33_ASAP7_75t_L g3821 ( 
.A1(n_3663),
.A2(n_3297),
.B1(n_3295),
.B2(n_2938),
.Y(n_3821)
);

INVxp67_ASAP7_75t_L g3822 ( 
.A(n_3586),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_L g3823 ( 
.A1(n_3678),
.A2(n_3297),
.B1(n_3295),
.B2(n_2939),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3645),
.B(n_2933),
.Y(n_3824)
);

OAI22xp5_ASAP7_75t_L g3825 ( 
.A1(n_3638),
.A2(n_3214),
.B1(n_3219),
.B2(n_3191),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3518),
.Y(n_3826)
);

CKINVDCx11_ASAP7_75t_R g3827 ( 
.A(n_3344),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3423),
.B(n_2933),
.Y(n_3828)
);

AOI22xp33_ASAP7_75t_L g3829 ( 
.A1(n_3477),
.A2(n_2959),
.B1(n_2995),
.B2(n_2939),
.Y(n_3829)
);

NOR2x1_ASAP7_75t_R g3830 ( 
.A(n_3347),
.B(n_2959),
.Y(n_3830)
);

AOI22xp33_ASAP7_75t_L g3831 ( 
.A1(n_3505),
.A2(n_2995),
.B1(n_3000),
.B2(n_2959),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3387),
.Y(n_3832)
);

AOI22xp33_ASAP7_75t_L g3833 ( 
.A1(n_3605),
.A2(n_3000),
.B1(n_3005),
.B2(n_2995),
.Y(n_3833)
);

AOI22xp33_ASAP7_75t_SL g3834 ( 
.A1(n_3415),
.A2(n_3005),
.B1(n_3025),
.B2(n_3000),
.Y(n_3834)
);

BUFx6f_ASAP7_75t_L g3835 ( 
.A(n_3648),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3314),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3314),
.Y(n_3837)
);

AOI22xp33_ASAP7_75t_L g3838 ( 
.A1(n_3507),
.A2(n_3025),
.B1(n_3033),
.B2(n_3005),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_SL g3839 ( 
.A1(n_3594),
.A2(n_3033),
.B1(n_3043),
.B2(n_3025),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3317),
.Y(n_3840)
);

BUFx4f_ASAP7_75t_SL g3841 ( 
.A(n_3429),
.Y(n_3841)
);

OAI22xp5_ASAP7_75t_SL g3842 ( 
.A1(n_3438),
.A2(n_3043),
.B1(n_3045),
.B2(n_3033),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_3369),
.B(n_3043),
.Y(n_3843)
);

HB1xp67_ASAP7_75t_L g3844 ( 
.A(n_3635),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3640),
.A2(n_3046),
.B1(n_3059),
.B2(n_3045),
.Y(n_3845)
);

AOI22xp33_ASAP7_75t_SL g3846 ( 
.A1(n_3594),
.A2(n_3046),
.B1(n_3059),
.B2(n_3045),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3383),
.B(n_3046),
.Y(n_3847)
);

OAI21xp5_ASAP7_75t_SL g3848 ( 
.A1(n_3471),
.A2(n_3070),
.B(n_3059),
.Y(n_3848)
);

AOI22xp33_ASAP7_75t_L g3849 ( 
.A1(n_3442),
.A2(n_3082),
.B1(n_3084),
.B2(n_3070),
.Y(n_3849)
);

AOI22xp33_ASAP7_75t_SL g3850 ( 
.A1(n_3343),
.A2(n_3082),
.B1(n_3084),
.B2(n_3070),
.Y(n_3850)
);

AOI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3557),
.A2(n_3084),
.B1(n_3095),
.B2(n_3082),
.Y(n_3851)
);

AOI211xp5_ASAP7_75t_L g3852 ( 
.A1(n_3514),
.A2(n_3102),
.B(n_3156),
.C(n_3095),
.Y(n_3852)
);

BUFx4f_ASAP7_75t_SL g3853 ( 
.A(n_3409),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3317),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3402),
.B(n_3095),
.Y(n_3855)
);

OAI22xp5_ASAP7_75t_L g3856 ( 
.A1(n_3568),
.A2(n_3214),
.B1(n_3219),
.B2(n_3191),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3318),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3630),
.A2(n_3219),
.B1(n_3223),
.B2(n_3214),
.Y(n_3858)
);

INVx1_ASAP7_75t_L g3859 ( 
.A(n_3318),
.Y(n_3859)
);

OAI21xp5_ASAP7_75t_SL g3860 ( 
.A1(n_3494),
.A2(n_3156),
.B(n_3102),
.Y(n_3860)
);

AOI21xp33_ASAP7_75t_L g3861 ( 
.A1(n_3489),
.A2(n_3156),
.B(n_3102),
.Y(n_3861)
);

BUFx3_ASAP7_75t_L g3862 ( 
.A(n_3484),
.Y(n_3862)
);

AOI222xp33_ASAP7_75t_L g3863 ( 
.A1(n_3351),
.A2(n_275),
.B1(n_277),
.B2(n_273),
.C1(n_274),
.C2(n_276),
.Y(n_3863)
);

AOI22xp33_ASAP7_75t_SL g3864 ( 
.A1(n_3343),
.A2(n_3223),
.B1(n_3224),
.B2(n_3183),
.Y(n_3864)
);

OAI22xp5_ASAP7_75t_L g3865 ( 
.A1(n_3593),
.A2(n_3286),
.B1(n_3289),
.B2(n_3275),
.Y(n_3865)
);

AOI22xp33_ASAP7_75t_L g3866 ( 
.A1(n_3545),
.A2(n_3223),
.B1(n_3224),
.B2(n_3183),
.Y(n_3866)
);

OAI222xp33_ASAP7_75t_L g3867 ( 
.A1(n_3667),
.A2(n_277),
.B1(n_279),
.B2(n_273),
.C1(n_275),
.C2(n_278),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3400),
.Y(n_3868)
);

BUFx5_ASAP7_75t_L g3869 ( 
.A(n_3685),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_L g3870 ( 
.A(n_3328),
.B(n_821),
.Y(n_3870)
);

OAI22xp33_ASAP7_75t_L g3871 ( 
.A1(n_3424),
.A2(n_3479),
.B1(n_3427),
.B2(n_3462),
.Y(n_3871)
);

OAI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3404),
.A2(n_3224),
.B1(n_3227),
.B2(n_3183),
.Y(n_3872)
);

OAI21xp33_ASAP7_75t_L g3873 ( 
.A1(n_3454),
.A2(n_3233),
.B(n_3227),
.Y(n_3873)
);

OAI22xp33_ASAP7_75t_L g3874 ( 
.A1(n_3479),
.A2(n_3233),
.B1(n_3275),
.B2(n_3227),
.Y(n_3874)
);

OAI22xp5_ASAP7_75t_SL g3875 ( 
.A1(n_3393),
.A2(n_3275),
.B1(n_3286),
.B2(n_3233),
.Y(n_3875)
);

AOI22xp33_ASAP7_75t_SL g3876 ( 
.A1(n_3362),
.A2(n_3289),
.B1(n_3292),
.B2(n_3286),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3576),
.A2(n_3292),
.B1(n_3289),
.B2(n_282),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_3449),
.B(n_3292),
.Y(n_3878)
);

NOR2xp33_ASAP7_75t_L g3879 ( 
.A(n_3330),
.B(n_821),
.Y(n_3879)
);

AOI22xp33_ASAP7_75t_L g3880 ( 
.A1(n_3525),
.A2(n_282),
.B1(n_278),
.B2(n_280),
.Y(n_3880)
);

OAI22xp5_ASAP7_75t_L g3881 ( 
.A1(n_3391),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3881)
);

AOI22xp33_ASAP7_75t_SL g3882 ( 
.A1(n_3362),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3882)
);

INVx4_ASAP7_75t_L g3883 ( 
.A(n_3648),
.Y(n_3883)
);

HB1xp67_ASAP7_75t_L g3884 ( 
.A(n_3536),
.Y(n_3884)
);

AOI22xp33_ASAP7_75t_SL g3885 ( 
.A1(n_3586),
.A2(n_290),
.B1(n_287),
.B2(n_289),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3400),
.Y(n_3886)
);

AOI22xp33_ASAP7_75t_L g3887 ( 
.A1(n_3449),
.A2(n_290),
.B1(n_287),
.B2(n_289),
.Y(n_3887)
);

INVx4_ASAP7_75t_L g3888 ( 
.A(n_3607),
.Y(n_3888)
);

AOI22xp33_ASAP7_75t_L g3889 ( 
.A1(n_3636),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_3889)
);

AOI22xp33_ASAP7_75t_L g3890 ( 
.A1(n_3427),
.A2(n_294),
.B1(n_291),
.B2(n_293),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3656),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3656),
.Y(n_3892)
);

OAI22xp5_ASAP7_75t_L g3893 ( 
.A1(n_3592),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_3893)
);

BUFx2_ASAP7_75t_L g3894 ( 
.A(n_3379),
.Y(n_3894)
);

INVx4_ASAP7_75t_L g3895 ( 
.A(n_3372),
.Y(n_3895)
);

INVx2_ASAP7_75t_SL g3896 ( 
.A(n_3347),
.Y(n_3896)
);

INVx4_ASAP7_75t_L g3897 ( 
.A(n_3372),
.Y(n_3897)
);

OAI21xp5_ASAP7_75t_SL g3898 ( 
.A1(n_3377),
.A2(n_295),
.B(n_296),
.Y(n_3898)
);

AOI22xp33_ASAP7_75t_L g3899 ( 
.A1(n_3462),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_SL g3900 ( 
.A1(n_3397),
.A2(n_302),
.B1(n_300),
.B2(n_301),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3665),
.Y(n_3901)
);

HB1xp67_ASAP7_75t_L g3902 ( 
.A(n_3548),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3410),
.B(n_303),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3421),
.B(n_303),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3683),
.A2(n_306),
.B1(n_304),
.B2(n_305),
.Y(n_3905)
);

BUFx2_ASAP7_75t_L g3906 ( 
.A(n_3688),
.Y(n_3906)
);

HB1xp67_ASAP7_75t_L g3907 ( 
.A(n_3603),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3665),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3440),
.A2(n_307),
.B1(n_304),
.B2(n_306),
.Y(n_3909)
);

INVx1_ASAP7_75t_SL g3910 ( 
.A(n_3476),
.Y(n_3910)
);

AOI22xp33_ASAP7_75t_L g3911 ( 
.A1(n_3595),
.A2(n_3669),
.B1(n_3558),
.B2(n_3553),
.Y(n_3911)
);

AOI22xp33_ASAP7_75t_L g3912 ( 
.A1(n_3553),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_3912)
);

AOI22xp33_ASAP7_75t_L g3913 ( 
.A1(n_3558),
.A2(n_3688),
.B1(n_3346),
.B2(n_3472),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3668),
.Y(n_3914)
);

OAI22xp5_ASAP7_75t_L g3915 ( 
.A1(n_3644),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_3915)
);

OAI22xp5_ASAP7_75t_L g3916 ( 
.A1(n_3524),
.A2(n_316),
.B1(n_312),
.B2(n_313),
.Y(n_3916)
);

OAI22xp5_ASAP7_75t_L g3917 ( 
.A1(n_3535),
.A2(n_3546),
.B1(n_3661),
.B2(n_3587),
.Y(n_3917)
);

CKINVDCx20_ASAP7_75t_R g3918 ( 
.A(n_3381),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_3617),
.B(n_317),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3628),
.A2(n_3599),
.B1(n_3564),
.B2(n_3512),
.Y(n_3920)
);

OAI22xp33_ASAP7_75t_L g3921 ( 
.A1(n_3382),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_3921)
);

AOI22xp33_ASAP7_75t_L g3922 ( 
.A1(n_3685),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_3922)
);

INVxp67_ASAP7_75t_L g3923 ( 
.A(n_3359),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3654),
.B(n_320),
.Y(n_3924)
);

INVx5_ASAP7_75t_SL g3925 ( 
.A(n_3408),
.Y(n_3925)
);

AOI22xp33_ASAP7_75t_L g3926 ( 
.A1(n_3666),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3668),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_3486),
.B(n_3496),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3653),
.B(n_835),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3652),
.A2(n_3676),
.B1(n_3542),
.B2(n_3538),
.Y(n_3930)
);

OAI22xp5_ASAP7_75t_L g3931 ( 
.A1(n_3382),
.A2(n_326),
.B1(n_322),
.B2(n_325),
.Y(n_3931)
);

AOI22xp33_ASAP7_75t_L g3932 ( 
.A1(n_3676),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_3932)
);

OAI22xp5_ASAP7_75t_L g3933 ( 
.A1(n_3486),
.A2(n_330),
.B1(n_327),
.B2(n_329),
.Y(n_3933)
);

INVx5_ASAP7_75t_SL g3934 ( 
.A(n_3443),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3432),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_L g3936 ( 
.A1(n_3527),
.A2(n_332),
.B1(n_329),
.B2(n_331),
.Y(n_3936)
);

AOI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3588),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3433),
.Y(n_3938)
);

INVx8_ASAP7_75t_L g3939 ( 
.A(n_3327),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3434),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3435),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3589),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3405),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_SL g3944 ( 
.A1(n_3543),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_3944)
);

AOI222xp33_ASAP7_75t_L g3945 ( 
.A1(n_3409),
.A2(n_340),
.B1(n_342),
.B2(n_337),
.C1(n_338),
.C2(n_341),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3655),
.B(n_341),
.Y(n_3946)
);

BUFx4f_ASAP7_75t_SL g3947 ( 
.A(n_3331),
.Y(n_3947)
);

OAI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3543),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_3948)
);

OR2x2_ASAP7_75t_L g3949 ( 
.A(n_3591),
.B(n_343),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_SL g3950 ( 
.A1(n_3660),
.A2(n_3368),
.B1(n_3396),
.B2(n_3452),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3600),
.A2(n_347),
.B1(n_344),
.B2(n_346),
.Y(n_3951)
);

INVx3_ASAP7_75t_L g3952 ( 
.A(n_3677),
.Y(n_3952)
);

AOI21xp33_ASAP7_75t_L g3953 ( 
.A1(n_3624),
.A2(n_3609),
.B(n_3585),
.Y(n_3953)
);

BUFx4f_ASAP7_75t_SL g3954 ( 
.A(n_3468),
.Y(n_3954)
);

OAI22xp5_ASAP7_75t_L g3955 ( 
.A1(n_3660),
.A2(n_349),
.B1(n_346),
.B2(n_348),
.Y(n_3955)
);

NOR2xp33_ASAP7_75t_L g3956 ( 
.A(n_3333),
.B(n_348),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3428),
.B(n_350),
.Y(n_3957)
);

NAND3xp33_ASAP7_75t_L g3958 ( 
.A(n_3647),
.B(n_351),
.C(n_352),
.Y(n_3958)
);

OAI21xp5_ASAP7_75t_SL g3959 ( 
.A1(n_3453),
.A2(n_353),
.B(n_354),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3696),
.A2(n_358),
.B1(n_355),
.B2(n_357),
.Y(n_3960)
);

AOI22xp5_ASAP7_75t_L g3961 ( 
.A1(n_3522),
.A2(n_359),
.B1(n_355),
.B2(n_358),
.Y(n_3961)
);

AND2x2_ASAP7_75t_L g3962 ( 
.A(n_3450),
.B(n_359),
.Y(n_3962)
);

HB1xp67_ASAP7_75t_L g3963 ( 
.A(n_3320),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3445),
.Y(n_3964)
);

OAI22xp5_ASAP7_75t_L g3965 ( 
.A1(n_3547),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3965)
);

INVx6_ASAP7_75t_L g3966 ( 
.A(n_3368),
.Y(n_3966)
);

OAI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_3619),
.A2(n_3419),
.B1(n_3616),
.B2(n_3612),
.Y(n_3967)
);

HB1xp67_ASAP7_75t_L g3968 ( 
.A(n_3348),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3451),
.Y(n_3969)
);

BUFx12f_ASAP7_75t_L g3970 ( 
.A(n_3396),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3465),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3460),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_L g3973 ( 
.A1(n_3475),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_3973)
);

NAND3xp33_ASAP7_75t_L g3974 ( 
.A(n_3650),
.B(n_364),
.C(n_365),
.Y(n_3974)
);

BUFx2_ASAP7_75t_L g3975 ( 
.A(n_3662),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3463),
.B(n_834),
.Y(n_3976)
);

AOI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3516),
.A2(n_368),
.B1(n_366),
.B2(n_367),
.Y(n_3977)
);

CKINVDCx11_ASAP7_75t_R g3978 ( 
.A(n_3413),
.Y(n_3978)
);

HB1xp67_ASAP7_75t_L g3979 ( 
.A(n_3371),
.Y(n_3979)
);

AOI222xp33_ASAP7_75t_L g3980 ( 
.A1(n_3327),
.A2(n_368),
.B1(n_370),
.B2(n_366),
.C1(n_367),
.C2(n_369),
.Y(n_3980)
);

HB1xp67_ASAP7_75t_L g3981 ( 
.A(n_3473),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3662),
.B(n_370),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3513),
.Y(n_3983)
);

INVx3_ASAP7_75t_L g3984 ( 
.A(n_3677),
.Y(n_3984)
);

OAI21xp33_ASAP7_75t_L g3985 ( 
.A1(n_3490),
.A2(n_371),
.B(n_372),
.Y(n_3985)
);

AOI22xp33_ASAP7_75t_L g3986 ( 
.A1(n_3692),
.A2(n_377),
.B1(n_374),
.B2(n_376),
.Y(n_3986)
);

HB1xp67_ASAP7_75t_L g3987 ( 
.A(n_3515),
.Y(n_3987)
);

INVx4_ASAP7_75t_L g3988 ( 
.A(n_3366),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3528),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_3989)
);

OAI21xp5_ASAP7_75t_SL g3990 ( 
.A1(n_3321),
.A2(n_378),
.B(n_380),
.Y(n_3990)
);

AOI22xp33_ASAP7_75t_L g3991 ( 
.A1(n_3537),
.A2(n_382),
.B1(n_380),
.B2(n_381),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3498),
.Y(n_3992)
);

OAI21xp33_ASAP7_75t_L g3993 ( 
.A1(n_3510),
.A2(n_382),
.B(n_383),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_L g3994 ( 
.A1(n_3551),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3580),
.A2(n_387),
.B1(n_384),
.B2(n_385),
.Y(n_3995)
);

OAI22xp5_ASAP7_75t_L g3996 ( 
.A1(n_3621),
.A2(n_389),
.B1(n_387),
.B2(n_388),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3684),
.Y(n_3997)
);

HB1xp67_ASAP7_75t_L g3998 ( 
.A(n_3521),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3523),
.Y(n_3999)
);

BUFx6f_ASAP7_75t_L g4000 ( 
.A(n_3325),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3529),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3539),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_4002)
);

OAI22xp5_ASAP7_75t_L g4003 ( 
.A1(n_3530),
.A2(n_392),
.B1(n_390),
.B2(n_391),
.Y(n_4003)
);

AOI22xp33_ASAP7_75t_L g4004 ( 
.A1(n_3569),
.A2(n_396),
.B1(n_394),
.B2(n_395),
.Y(n_4004)
);

BUFx2_ASAP7_75t_L g4005 ( 
.A(n_3684),
.Y(n_4005)
);

BUFx4f_ASAP7_75t_SL g4006 ( 
.A(n_3598),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3531),
.Y(n_4007)
);

AOI22xp33_ASAP7_75t_SL g4008 ( 
.A1(n_3499),
.A2(n_397),
.B1(n_394),
.B2(n_396),
.Y(n_4008)
);

AOI22xp33_ASAP7_75t_L g4009 ( 
.A1(n_3572),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_4009)
);

BUFx6f_ASAP7_75t_L g4010 ( 
.A(n_3325),
.Y(n_4010)
);

AOI22xp5_ASAP7_75t_L g4011 ( 
.A1(n_3959),
.A2(n_3990),
.B1(n_3706),
.B2(n_3699),
.Y(n_4011)
);

INVx2_ASAP7_75t_L g4012 ( 
.A(n_3981),
.Y(n_4012)
);

AOI22xp33_ASAP7_75t_L g4013 ( 
.A1(n_3757),
.A2(n_3689),
.B1(n_3418),
.B2(n_3420),
.Y(n_4013)
);

AOI22xp33_ASAP7_75t_L g4014 ( 
.A1(n_3709),
.A2(n_3694),
.B1(n_3562),
.B2(n_3554),
.Y(n_4014)
);

OAI22xp5_ASAP7_75t_L g4015 ( 
.A1(n_3716),
.A2(n_3570),
.B1(n_3682),
.B2(n_3651),
.Y(n_4015)
);

AOI22xp33_ASAP7_75t_L g4016 ( 
.A1(n_3727),
.A2(n_3550),
.B1(n_3555),
.B2(n_3544),
.Y(n_4016)
);

AOI22xp33_ASAP7_75t_L g4017 ( 
.A1(n_3863),
.A2(n_3565),
.B1(n_3566),
.B2(n_3559),
.Y(n_4017)
);

OAI222xp33_ASAP7_75t_L g4018 ( 
.A1(n_3742),
.A2(n_3577),
.B1(n_3574),
.B2(n_3582),
.C1(n_3578),
.C2(n_3567),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3945),
.A2(n_3917),
.B1(n_3900),
.B2(n_3980),
.Y(n_4019)
);

OAI22xp33_ASAP7_75t_L g4020 ( 
.A1(n_3898),
.A2(n_3501),
.B1(n_3345),
.B2(n_3631),
.Y(n_4020)
);

OAI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3705),
.A2(n_3649),
.B1(n_3597),
.B2(n_3560),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3712),
.B(n_3583),
.Y(n_4022)
);

NAND3xp33_ASAP7_75t_L g4023 ( 
.A(n_3720),
.B(n_3602),
.C(n_3671),
.Y(n_4023)
);

OAI22xp5_ASAP7_75t_L g4024 ( 
.A1(n_3895),
.A2(n_3356),
.B1(n_3627),
.B2(n_3455),
.Y(n_4024)
);

OAI21xp5_ASAP7_75t_L g4025 ( 
.A1(n_3867),
.A2(n_3611),
.B(n_3483),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3701),
.Y(n_4026)
);

OAI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3895),
.A2(n_3520),
.B1(n_3519),
.B2(n_3366),
.Y(n_4027)
);

AOI22xp33_ASAP7_75t_SL g4028 ( 
.A1(n_3920),
.A2(n_3519),
.B1(n_3455),
.B2(n_3601),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3717),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3987),
.Y(n_4030)
);

OAI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3897),
.A2(n_3637),
.B1(n_3646),
.B2(n_3466),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3963),
.B(n_3968),
.Y(n_4032)
);

OAI22xp5_ASAP7_75t_L g4033 ( 
.A1(n_3897),
.A2(n_3629),
.B1(n_3674),
.B2(n_3657),
.Y(n_4033)
);

AOI22xp33_ASAP7_75t_SL g4034 ( 
.A1(n_3726),
.A2(n_3406),
.B1(n_3480),
.B2(n_3392),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_L g4035 ( 
.A1(n_3729),
.A2(n_3681),
.B1(n_3657),
.B2(n_3674),
.Y(n_4035)
);

OAI22xp5_ASAP7_75t_L g4036 ( 
.A1(n_3760),
.A2(n_3502),
.B1(n_3563),
.B2(n_3658),
.Y(n_4036)
);

AOI22xp33_ASAP7_75t_L g4037 ( 
.A1(n_3871),
.A2(n_3575),
.B1(n_3614),
.B2(n_3446),
.Y(n_4037)
);

AOI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_3718),
.A2(n_3416),
.B1(n_3506),
.B2(n_3670),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3722),
.Y(n_4039)
);

OAI221xp5_ASAP7_75t_L g4040 ( 
.A1(n_3885),
.A2(n_3540),
.B1(n_3430),
.B2(n_3412),
.C(n_3425),
.Y(n_4040)
);

AOI22xp33_ASAP7_75t_L g4041 ( 
.A1(n_3728),
.A2(n_3680),
.B1(n_3388),
.B2(n_3541),
.Y(n_4041)
);

AOI22xp33_ASAP7_75t_L g4042 ( 
.A1(n_3881),
.A2(n_3691),
.B1(n_3388),
.B2(n_3541),
.Y(n_4042)
);

OAI211xp5_ASAP7_75t_SL g4043 ( 
.A1(n_3808),
.A2(n_3464),
.B(n_3425),
.C(n_3412),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3998),
.Y(n_4044)
);

AOI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_3731),
.A2(n_3388),
.B1(n_3541),
.B2(n_3325),
.Y(n_4045)
);

AOI22xp33_ASAP7_75t_SL g4046 ( 
.A1(n_3726),
.A2(n_3608),
.B1(n_3615),
.B2(n_3561),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3745),
.A2(n_3691),
.B1(n_3608),
.B2(n_3615),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3734),
.Y(n_4048)
);

NAND3xp33_ASAP7_75t_L g4049 ( 
.A(n_3974),
.B(n_3691),
.C(n_3608),
.Y(n_4049)
);

OAI22xp5_ASAP7_75t_L g4050 ( 
.A1(n_3760),
.A2(n_3615),
.B1(n_3672),
.B2(n_3561),
.Y(n_4050)
);

NOR3xp33_ASAP7_75t_L g4051 ( 
.A(n_3724),
.B(n_3982),
.C(n_3732),
.Y(n_4051)
);

AOI22xp33_ASAP7_75t_L g4052 ( 
.A1(n_3745),
.A2(n_3672),
.B1(n_3687),
.B2(n_3561),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_L g4053 ( 
.A1(n_3714),
.A2(n_3687),
.B1(n_3672),
.B2(n_402),
.Y(n_4053)
);

AOI22xp33_ASAP7_75t_L g4054 ( 
.A1(n_3735),
.A2(n_3687),
.B1(n_402),
.B2(n_399),
.Y(n_4054)
);

AOI22xp33_ASAP7_75t_L g4055 ( 
.A1(n_3746),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_3753),
.B(n_403),
.Y(n_4056)
);

AOI22xp5_ASAP7_75t_L g4057 ( 
.A1(n_3761),
.A2(n_408),
.B1(n_404),
.B2(n_407),
.Y(n_4057)
);

AOI221xp5_ASAP7_75t_L g4058 ( 
.A1(n_3737),
.A2(n_410),
.B1(n_407),
.B2(n_409),
.C(n_411),
.Y(n_4058)
);

AOI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3882),
.A2(n_3931),
.B1(n_3921),
.B2(n_3965),
.Y(n_4059)
);

AOI22xp33_ASAP7_75t_L g4060 ( 
.A1(n_4008),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4060)
);

AOI22xp33_ASAP7_75t_L g4061 ( 
.A1(n_3953),
.A2(n_415),
.B1(n_412),
.B2(n_414),
.Y(n_4061)
);

AOI22xp33_ASAP7_75t_L g4062 ( 
.A1(n_3916),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_4062)
);

AOI22xp33_ASAP7_75t_L g4063 ( 
.A1(n_3944),
.A2(n_419),
.B1(n_416),
.B2(n_418),
.Y(n_4063)
);

AOI22xp33_ASAP7_75t_SL g4064 ( 
.A1(n_3767),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3979),
.Y(n_4065)
);

AOI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_3912),
.A2(n_426),
.B1(n_422),
.B2(n_423),
.Y(n_4066)
);

AOI22xp33_ASAP7_75t_L g4067 ( 
.A1(n_3708),
.A2(n_426),
.B1(n_422),
.B2(n_423),
.Y(n_4067)
);

NAND3xp33_ASAP7_75t_L g4068 ( 
.A(n_3958),
.B(n_428),
.C(n_429),
.Y(n_4068)
);

INVx2_ASAP7_75t_L g4069 ( 
.A(n_3756),
.Y(n_4069)
);

AOI22xp33_ASAP7_75t_L g4070 ( 
.A1(n_3985),
.A2(n_430),
.B1(n_428),
.B2(n_429),
.Y(n_4070)
);

AOI22xp33_ASAP7_75t_L g4071 ( 
.A1(n_3985),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3741),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3764),
.B(n_3750),
.Y(n_4073)
);

AOI22xp33_ASAP7_75t_L g4074 ( 
.A1(n_3993),
.A2(n_436),
.B1(n_433),
.B2(n_434),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3999),
.B(n_433),
.Y(n_4075)
);

AOI22xp33_ASAP7_75t_L g4076 ( 
.A1(n_3993),
.A2(n_438),
.B1(n_434),
.B2(n_437),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_4003),
.A2(n_439),
.B1(n_437),
.B2(n_438),
.Y(n_4077)
);

AOI22xp33_ASAP7_75t_L g4078 ( 
.A1(n_3915),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_4078)
);

AOI22xp33_ASAP7_75t_L g4079 ( 
.A1(n_3893),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_4079)
);

OAI221xp5_ASAP7_75t_SL g4080 ( 
.A1(n_3961),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.C(n_446),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_SL g4081 ( 
.A1(n_3767),
.A2(n_446),
.B1(n_443),
.B2(n_445),
.Y(n_4081)
);

AOI22xp33_ASAP7_75t_L g4082 ( 
.A1(n_3719),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_4082)
);

AOI22xp33_ASAP7_75t_SL g4083 ( 
.A1(n_3816),
.A2(n_450),
.B1(n_448),
.B2(n_449),
.Y(n_4083)
);

AOI22xp33_ASAP7_75t_L g4084 ( 
.A1(n_3736),
.A2(n_3844),
.B1(n_3899),
.B2(n_3890),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_L g4085 ( 
.A1(n_3986),
.A2(n_452),
.B1(n_450),
.B2(n_451),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3842),
.B(n_451),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_3961),
.A2(n_454),
.B1(n_452),
.B2(n_453),
.Y(n_4087)
);

AOI22xp33_ASAP7_75t_L g4088 ( 
.A1(n_3879),
.A2(n_458),
.B1(n_454),
.B2(n_456),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_4001),
.B(n_456),
.Y(n_4089)
);

NOR3xp33_ASAP7_75t_L g4090 ( 
.A(n_3704),
.B(n_458),
.C(n_459),
.Y(n_4090)
);

AOI22xp33_ASAP7_75t_L g4091 ( 
.A1(n_3884),
.A2(n_463),
.B1(n_460),
.B2(n_461),
.Y(n_4091)
);

AOI22xp5_ASAP7_75t_L g4092 ( 
.A1(n_4002),
.A2(n_467),
.B1(n_465),
.B2(n_466),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3759),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3730),
.B(n_834),
.Y(n_4094)
);

AOI22xp33_ASAP7_75t_L g4095 ( 
.A1(n_3902),
.A2(n_468),
.B1(n_466),
.B2(n_467),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3781),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3744),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_4007),
.B(n_468),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3748),
.Y(n_4099)
);

OAI22xp5_ASAP7_75t_L g4100 ( 
.A1(n_3707),
.A2(n_472),
.B1(n_469),
.B2(n_470),
.Y(n_4100)
);

AOI22xp33_ASAP7_75t_L g4101 ( 
.A1(n_3907),
.A2(n_473),
.B1(n_470),
.B2(n_472),
.Y(n_4101)
);

HB1xp67_ASAP7_75t_L g4102 ( 
.A(n_3770),
.Y(n_4102)
);

OAI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_3887),
.A2(n_478),
.B1(n_474),
.B2(n_476),
.Y(n_4103)
);

INVx2_ASAP7_75t_L g4104 ( 
.A(n_3789),
.Y(n_4104)
);

AOI22xp33_ASAP7_75t_L g4105 ( 
.A1(n_3771),
.A2(n_479),
.B1(n_474),
.B2(n_476),
.Y(n_4105)
);

AOI22xp33_ASAP7_75t_L g4106 ( 
.A1(n_4004),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_SL g4107 ( 
.A(n_3952),
.B(n_481),
.Y(n_4107)
);

OAI22xp5_ASAP7_75t_L g4108 ( 
.A1(n_3888),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_4108)
);

OAI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3933),
.A2(n_485),
.B(n_487),
.Y(n_4109)
);

AOI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_4009),
.A2(n_489),
.B1(n_487),
.B2(n_488),
.Y(n_4110)
);

OAI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3888),
.A2(n_492),
.B1(n_488),
.B2(n_490),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_3784),
.B(n_490),
.Y(n_4112)
);

AOI222xp33_ASAP7_75t_L g4113 ( 
.A1(n_3919),
.A2(n_495),
.B1(n_497),
.B2(n_493),
.C1(n_494),
.C2(n_496),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3889),
.A2(n_497),
.B1(n_493),
.B2(n_494),
.Y(n_4114)
);

OAI22xp5_ASAP7_75t_L g4115 ( 
.A1(n_3725),
.A2(n_501),
.B1(n_499),
.B2(n_500),
.Y(n_4115)
);

AOI22xp33_ASAP7_75t_L g4116 ( 
.A1(n_3996),
.A2(n_502),
.B1(n_499),
.B2(n_500),
.Y(n_4116)
);

OAI22xp5_ASAP7_75t_L g4117 ( 
.A1(n_3950),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3813),
.Y(n_4118)
);

OAI221xp5_ASAP7_75t_L g4119 ( 
.A1(n_3991),
.A2(n_507),
.B1(n_505),
.B2(n_506),
.C(n_508),
.Y(n_4119)
);

OAI21xp5_ASAP7_75t_SL g4120 ( 
.A1(n_3711),
.A2(n_505),
.B(n_507),
.Y(n_4120)
);

AOI22xp33_ASAP7_75t_L g4121 ( 
.A1(n_3994),
.A2(n_3905),
.B1(n_3926),
.B2(n_3913),
.Y(n_4121)
);

AOI22xp33_ASAP7_75t_L g4122 ( 
.A1(n_3948),
.A2(n_510),
.B1(n_508),
.B2(n_509),
.Y(n_4122)
);

AOI22xp33_ASAP7_75t_L g4123 ( 
.A1(n_3955),
.A2(n_512),
.B1(n_509),
.B2(n_511),
.Y(n_4123)
);

INVx2_ASAP7_75t_SL g4124 ( 
.A(n_3749),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3794),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3819),
.B(n_513),
.Y(n_4126)
);

OAI22xp33_ASAP7_75t_L g4127 ( 
.A1(n_3883),
.A2(n_518),
.B1(n_514),
.B2(n_515),
.Y(n_4127)
);

OAI22xp5_ASAP7_75t_L g4128 ( 
.A1(n_3930),
.A2(n_519),
.B1(n_515),
.B2(n_518),
.Y(n_4128)
);

AOI22xp33_ASAP7_75t_SL g4129 ( 
.A1(n_3752),
.A2(n_523),
.B1(n_520),
.B2(n_522),
.Y(n_4129)
);

AOI22xp33_ASAP7_75t_L g4130 ( 
.A1(n_3924),
.A2(n_524),
.B1(n_522),
.B2(n_523),
.Y(n_4130)
);

OAI22x1_ASAP7_75t_L g4131 ( 
.A1(n_3906),
.A2(n_528),
.B1(n_526),
.B2(n_527),
.Y(n_4131)
);

OAI22xp5_ASAP7_75t_L g4132 ( 
.A1(n_3804),
.A2(n_530),
.B1(n_526),
.B2(n_529),
.Y(n_4132)
);

INVxp67_ASAP7_75t_L g4133 ( 
.A(n_3894),
.Y(n_4133)
);

AOI22xp33_ASAP7_75t_L g4134 ( 
.A1(n_3956),
.A2(n_531),
.B1(n_529),
.B2(n_530),
.Y(n_4134)
);

AOI22xp33_ASAP7_75t_L g4135 ( 
.A1(n_3880),
.A2(n_533),
.B1(n_531),
.B2(n_532),
.Y(n_4135)
);

AOI22xp33_ASAP7_75t_L g4136 ( 
.A1(n_3989),
.A2(n_536),
.B1(n_534),
.B2(n_535),
.Y(n_4136)
);

NOR2xp67_ASAP7_75t_L g4137 ( 
.A(n_3883),
.B(n_3702),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_3740),
.B(n_833),
.Y(n_4138)
);

AOI22xp33_ASAP7_75t_L g4139 ( 
.A1(n_3751),
.A2(n_537),
.B1(n_534),
.B2(n_536),
.Y(n_4139)
);

AOI22xp33_ASAP7_75t_L g4140 ( 
.A1(n_3960),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.Y(n_4140)
);

AOI22xp33_ASAP7_75t_L g4141 ( 
.A1(n_3896),
.A2(n_542),
.B1(n_539),
.B2(n_541),
.Y(n_4141)
);

OAI221xp5_ASAP7_75t_L g4142 ( 
.A1(n_3747),
.A2(n_543),
.B1(n_541),
.B2(n_542),
.C(n_544),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3826),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3935),
.B(n_545),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3938),
.B(n_546),
.Y(n_4145)
);

OAI222xp33_ASAP7_75t_L g4146 ( 
.A1(n_3928),
.A2(n_546),
.B1(n_547),
.B2(n_548),
.C1(n_550),
.C2(n_551),
.Y(n_4146)
);

AOI22xp33_ASAP7_75t_L g4147 ( 
.A1(n_3792),
.A2(n_550),
.B1(n_547),
.B2(n_548),
.Y(n_4147)
);

NAND3xp33_ASAP7_75t_L g4148 ( 
.A(n_3776),
.B(n_552),
.C(n_553),
.Y(n_4148)
);

AOI22xp33_ASAP7_75t_L g4149 ( 
.A1(n_3795),
.A2(n_555),
.B1(n_552),
.B2(n_554),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_3832),
.B(n_832),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_3995),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_4151)
);

AOI22xp33_ASAP7_75t_L g4152 ( 
.A1(n_3973),
.A2(n_558),
.B1(n_556),
.B2(n_557),
.Y(n_4152)
);

AOI22xp33_ASAP7_75t_L g4153 ( 
.A1(n_3977),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.Y(n_4153)
);

AOI22xp33_ASAP7_75t_SL g4154 ( 
.A1(n_3975),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.Y(n_4154)
);

OAI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_3909),
.A2(n_561),
.B(n_562),
.Y(n_4155)
);

AOI22xp33_ASAP7_75t_L g4156 ( 
.A1(n_3877),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_4156)
);

AOI22xp33_ASAP7_75t_SL g4157 ( 
.A1(n_3939),
.A2(n_567),
.B1(n_565),
.B2(n_566),
.Y(n_4157)
);

OR2x2_ASAP7_75t_L g4158 ( 
.A(n_3940),
.B(n_565),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3941),
.Y(n_4159)
);

OAI22xp5_ASAP7_75t_L g4160 ( 
.A1(n_3763),
.A2(n_569),
.B1(n_566),
.B2(n_568),
.Y(n_4160)
);

AOI22xp33_ASAP7_75t_L g4161 ( 
.A1(n_3755),
.A2(n_3765),
.B1(n_3788),
.B2(n_3791),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3943),
.B(n_3972),
.Y(n_4162)
);

AOI222xp33_ASAP7_75t_L g4163 ( 
.A1(n_3853),
.A2(n_568),
.B1(n_569),
.B2(n_570),
.C1(n_571),
.C2(n_572),
.Y(n_4163)
);

BUFx12f_ASAP7_75t_L g4164 ( 
.A(n_3978),
.Y(n_4164)
);

AOI22xp33_ASAP7_75t_L g4165 ( 
.A1(n_3777),
.A2(n_573),
.B1(n_571),
.B2(n_572),
.Y(n_4165)
);

AOI22xp33_ASAP7_75t_L g4166 ( 
.A1(n_3870),
.A2(n_576),
.B1(n_573),
.B2(n_575),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3964),
.B(n_575),
.Y(n_4167)
);

AOI22xp33_ASAP7_75t_SL g4168 ( 
.A1(n_3939),
.A2(n_580),
.B1(n_577),
.B2(n_579),
.Y(n_4168)
);

NOR3xp33_ASAP7_75t_L g4169 ( 
.A(n_3929),
.B(n_579),
.C(n_580),
.Y(n_4169)
);

AOI22xp33_ASAP7_75t_SL g4170 ( 
.A1(n_3939),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_4170)
);

OAI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_3849),
.A2(n_584),
.B1(n_581),
.B2(n_583),
.Y(n_4171)
);

AO222x2_ASAP7_75t_SL g4172 ( 
.A1(n_3768),
.A2(n_585),
.B1(n_586),
.B2(n_588),
.C1(n_590),
.C2(n_591),
.Y(n_4172)
);

OAI221xp5_ASAP7_75t_L g4173 ( 
.A1(n_3786),
.A2(n_592),
.B1(n_585),
.B2(n_591),
.C(n_593),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_SL g4174 ( 
.A1(n_4005),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_3946),
.A2(n_596),
.B1(n_594),
.B2(n_595),
.Y(n_4175)
);

AND2x4_ASAP7_75t_L g4176 ( 
.A(n_3836),
.B(n_596),
.Y(n_4176)
);

AOI22xp33_ASAP7_75t_L g4177 ( 
.A1(n_3967),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_4177)
);

AOI22xp5_ASAP7_75t_L g4178 ( 
.A1(n_3796),
.A2(n_601),
.B1(n_597),
.B2(n_600),
.Y(n_4178)
);

AOI22xp33_ASAP7_75t_L g4179 ( 
.A1(n_3873),
.A2(n_602),
.B1(n_600),
.B2(n_601),
.Y(n_4179)
);

OA21x2_ASAP7_75t_L g4180 ( 
.A1(n_3829),
.A2(n_602),
.B(n_603),
.Y(n_4180)
);

AOI22xp33_ASAP7_75t_L g4181 ( 
.A1(n_3869),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3969),
.B(n_606),
.Y(n_4182)
);

AOI22xp33_ASAP7_75t_SL g4183 ( 
.A1(n_3869),
.A2(n_610),
.B1(n_606),
.B2(n_607),
.Y(n_4183)
);

AOI22xp33_ASAP7_75t_L g4184 ( 
.A1(n_3869),
.A2(n_611),
.B1(n_607),
.B2(n_610),
.Y(n_4184)
);

NOR2xp33_ASAP7_75t_L g4185 ( 
.A(n_3910),
.B(n_611),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_SL g4186 ( 
.A1(n_3830),
.A2(n_612),
.B(n_613),
.Y(n_4186)
);

AOI221xp5_ASAP7_75t_L g4187 ( 
.A1(n_3758),
.A2(n_613),
.B1(n_614),
.B2(n_615),
.C(n_616),
.Y(n_4187)
);

OAI221xp5_ASAP7_75t_SL g4188 ( 
.A1(n_3911),
.A2(n_615),
.B1(n_617),
.B2(n_619),
.C(n_620),
.Y(n_4188)
);

AOI22xp33_ASAP7_75t_L g4189 ( 
.A1(n_3869),
.A2(n_622),
.B1(n_617),
.B2(n_621),
.Y(n_4189)
);

AOI222xp33_ASAP7_75t_L g4190 ( 
.A1(n_3822),
.A2(n_621),
.B1(n_623),
.B2(n_624),
.C1(n_625),
.C2(n_627),
.Y(n_4190)
);

AOI22xp33_ASAP7_75t_SL g4191 ( 
.A1(n_3869),
.A2(n_628),
.B1(n_624),
.B2(n_627),
.Y(n_4191)
);

AOI22xp33_ASAP7_75t_L g4192 ( 
.A1(n_3966),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_4192)
);

AOI22xp33_ASAP7_75t_L g4193 ( 
.A1(n_3966),
.A2(n_3779),
.B1(n_3932),
.B2(n_3922),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_3988),
.A2(n_631),
.B1(n_629),
.B2(n_630),
.Y(n_4194)
);

AND2x2_ASAP7_75t_L g4195 ( 
.A(n_3983),
.B(n_631),
.Y(n_4195)
);

OAI22xp5_ASAP7_75t_L g4196 ( 
.A1(n_3988),
.A2(n_634),
.B1(n_632),
.B2(n_633),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_3971),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3992),
.Y(n_4198)
);

AOI22xp33_ASAP7_75t_SL g4199 ( 
.A1(n_3818),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_4199)
);

AOI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3773),
.A2(n_638),
.B1(n_635),
.B2(n_637),
.Y(n_4200)
);

INVx2_ASAP7_75t_SL g4201 ( 
.A(n_3698),
.Y(n_4201)
);

AOI22xp33_ASAP7_75t_L g4202 ( 
.A1(n_3785),
.A2(n_3937),
.B1(n_3942),
.B2(n_3936),
.Y(n_4202)
);

NAND3xp33_ASAP7_75t_L g4203 ( 
.A(n_3951),
.B(n_638),
.C(n_639),
.Y(n_4203)
);

AOI22xp33_ASAP7_75t_L g4204 ( 
.A1(n_3797),
.A2(n_644),
.B1(n_641),
.B2(n_642),
.Y(n_4204)
);

AOI22xp33_ASAP7_75t_SL g4205 ( 
.A1(n_3952),
.A2(n_644),
.B1(n_641),
.B2(n_642),
.Y(n_4205)
);

OA21x2_ASAP7_75t_L g4206 ( 
.A1(n_3848),
.A2(n_645),
.B(n_646),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3837),
.Y(n_4207)
);

AOI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_3787),
.A2(n_647),
.B1(n_645),
.B2(n_646),
.Y(n_4208)
);

OAI21xp5_ASAP7_75t_SL g4209 ( 
.A1(n_3775),
.A2(n_647),
.B(n_649),
.Y(n_4209)
);

AOI22xp33_ASAP7_75t_SL g4210 ( 
.A1(n_3856),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_3713),
.B(n_650),
.Y(n_4211)
);

OAI222xp33_ASAP7_75t_L g4212 ( 
.A1(n_3825),
.A2(n_651),
.B1(n_652),
.B2(n_654),
.C1(n_655),
.C2(n_656),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3840),
.Y(n_4213)
);

OAI221xp5_ASAP7_75t_L g4214 ( 
.A1(n_3703),
.A2(n_654),
.B1(n_655),
.B2(n_657),
.C(n_659),
.Y(n_4214)
);

AND2x2_ASAP7_75t_L g4215 ( 
.A(n_4073),
.B(n_3854),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4102),
.B(n_3857),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4012),
.B(n_3859),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4030),
.B(n_3868),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_4065),
.B(n_3886),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4044),
.B(n_3891),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_R g4221 ( 
.A(n_4164),
.B(n_3772),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4032),
.B(n_3892),
.Y(n_4222)
);

AND2x2_ASAP7_75t_L g4223 ( 
.A(n_4133),
.B(n_3901),
.Y(n_4223)
);

OAI221xp5_ASAP7_75t_L g4224 ( 
.A1(n_4120),
.A2(n_3814),
.B1(n_3778),
.B2(n_3831),
.C(n_3923),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4162),
.B(n_3908),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_4026),
.B(n_4029),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4039),
.B(n_3914),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4048),
.B(n_3927),
.Y(n_4228)
);

OAI22xp5_ASAP7_75t_L g4229 ( 
.A1(n_4017),
.A2(n_3780),
.B1(n_3845),
.B2(n_3838),
.Y(n_4229)
);

AND2x2_ASAP7_75t_L g4230 ( 
.A(n_4072),
.B(n_3817),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4097),
.B(n_3798),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4099),
.B(n_3721),
.Y(n_4232)
);

AND2x2_ASAP7_75t_L g4233 ( 
.A(n_4118),
.B(n_4159),
.Y(n_4233)
);

NAND3xp33_ASAP7_75t_L g4234 ( 
.A(n_4051),
.B(n_3851),
.C(n_3903),
.Y(n_4234)
);

NAND2xp5_ASAP7_75t_L g4235 ( 
.A(n_4197),
.B(n_3733),
.Y(n_4235)
);

OAI21xp5_ASAP7_75t_SL g4236 ( 
.A1(n_4209),
.A2(n_3860),
.B(n_3700),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_4198),
.B(n_3817),
.Y(n_4237)
);

OAI21xp33_ASAP7_75t_L g4238 ( 
.A1(n_4019),
.A2(n_3811),
.B(n_3810),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4022),
.B(n_4069),
.Y(n_4239)
);

NAND2xp5_ASAP7_75t_L g4240 ( 
.A(n_4207),
.B(n_3828),
.Y(n_4240)
);

AND2x2_ASAP7_75t_L g4241 ( 
.A(n_4093),
.B(n_3984),
.Y(n_4241)
);

OAI21xp33_ASAP7_75t_L g4242 ( 
.A1(n_4011),
.A2(n_3904),
.B(n_3807),
.Y(n_4242)
);

OAI21xp33_ASAP7_75t_SL g4243 ( 
.A1(n_4137),
.A2(n_3801),
.B(n_3702),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_4213),
.B(n_3809),
.Y(n_4244)
);

NAND3xp33_ASAP7_75t_L g4245 ( 
.A(n_4028),
.B(n_3823),
.C(n_3801),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_4096),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_4104),
.B(n_3824),
.Y(n_4247)
);

NOR3xp33_ASAP7_75t_L g4248 ( 
.A(n_4146),
.B(n_4188),
.C(n_4148),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_4125),
.B(n_3984),
.Y(n_4249)
);

NAND3xp33_ASAP7_75t_L g4250 ( 
.A(n_4023),
.B(n_3852),
.C(n_3949),
.Y(n_4250)
);

OAI221xp5_ASAP7_75t_SL g4251 ( 
.A1(n_4172),
.A2(n_3799),
.B1(n_3833),
.B2(n_3800),
.C(n_3821),
.Y(n_4251)
);

BUFx3_ASAP7_75t_L g4252 ( 
.A(n_4124),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4143),
.B(n_3843),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_4094),
.B(n_3847),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_4176),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4056),
.B(n_3997),
.Y(n_4256)
);

OAI221xp5_ASAP7_75t_SL g4257 ( 
.A1(n_4020),
.A2(n_3866),
.B1(n_3803),
.B2(n_3815),
.C(n_3802),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_4016),
.B(n_3855),
.Y(n_4258)
);

OAI21xp33_ASAP7_75t_L g4259 ( 
.A1(n_4057),
.A2(n_4185),
.B(n_4168),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4161),
.B(n_3957),
.Y(n_4260)
);

AND2x2_ASAP7_75t_L g4261 ( 
.A(n_4138),
.B(n_3997),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_SL g4262 ( 
.A(n_4034),
.B(n_3698),
.Y(n_4262)
);

AOI221xp5_ASAP7_75t_L g4263 ( 
.A1(n_4188),
.A2(n_3976),
.B1(n_3962),
.B2(n_3782),
.C(n_3820),
.Y(n_4263)
);

OAI22xp5_ASAP7_75t_L g4264 ( 
.A1(n_4129),
.A2(n_3738),
.B1(n_3769),
.B2(n_3762),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4034),
.B(n_3698),
.Y(n_4265)
);

OAI21xp5_ASAP7_75t_SL g4266 ( 
.A1(n_4043),
.A2(n_3835),
.B(n_3700),
.Y(n_4266)
);

NAND3xp33_ASAP7_75t_L g4267 ( 
.A(n_4090),
.B(n_4014),
.C(n_4163),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4176),
.B(n_3700),
.Y(n_4268)
);

OAI21xp5_ASAP7_75t_SL g4269 ( 
.A1(n_4043),
.A2(n_3835),
.B(n_3805),
.Y(n_4269)
);

NAND4xp25_ASAP7_75t_SL g4270 ( 
.A(n_4037),
.B(n_4190),
.C(n_3918),
.D(n_4169),
.Y(n_4270)
);

NOR2xp33_ASAP7_75t_L g4271 ( 
.A(n_4040),
.B(n_3710),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4211),
.B(n_3865),
.Y(n_4272)
);

OAI22xp5_ASAP7_75t_L g4273 ( 
.A1(n_4129),
.A2(n_4191),
.B1(n_4183),
.B2(n_4080),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_4150),
.B(n_3872),
.Y(n_4274)
);

OAI21xp5_ASAP7_75t_SL g4275 ( 
.A1(n_4027),
.A2(n_3835),
.B(n_3806),
.Y(n_4275)
);

OAI22xp5_ASAP7_75t_L g4276 ( 
.A1(n_4183),
.A2(n_3846),
.B1(n_3839),
.B2(n_3850),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_L g4277 ( 
.A(n_4195),
.B(n_3858),
.Y(n_4277)
);

AOI221xp5_ASAP7_75t_L g4278 ( 
.A1(n_4131),
.A2(n_3862),
.B1(n_3793),
.B2(n_3874),
.C(n_3812),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4201),
.B(n_4010),
.Y(n_4279)
);

NOR3xp33_ASAP7_75t_L g4280 ( 
.A(n_4146),
.B(n_3827),
.C(n_3861),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4031),
.B(n_3864),
.Y(n_4281)
);

OAI221xp5_ASAP7_75t_L g4282 ( 
.A1(n_4121),
.A2(n_3743),
.B1(n_3723),
.B2(n_3876),
.C(n_3834),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_SL g4283 ( 
.A(n_4024),
.B(n_4046),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4038),
.B(n_4000),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4112),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4045),
.B(n_4000),
.Y(n_4286)
);

OAI21xp5_ASAP7_75t_SL g4287 ( 
.A1(n_4157),
.A2(n_3878),
.B(n_3754),
.Y(n_4287)
);

INVx2_ASAP7_75t_L g4288 ( 
.A(n_4158),
.Y(n_4288)
);

NAND3xp33_ASAP7_75t_L g4289 ( 
.A(n_4191),
.B(n_4010),
.C(n_4000),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4013),
.B(n_4010),
.Y(n_4290)
);

AND2x2_ASAP7_75t_L g4291 ( 
.A(n_4041),
.B(n_3754),
.Y(n_4291)
);

NAND3xp33_ASAP7_75t_L g4292 ( 
.A(n_4157),
.B(n_3774),
.C(n_3766),
.Y(n_4292)
);

NAND3xp33_ASAP7_75t_L g4293 ( 
.A(n_4168),
.B(n_3947),
.C(n_3875),
.Y(n_4293)
);

OAI221xp5_ASAP7_75t_SL g4294 ( 
.A1(n_4059),
.A2(n_3934),
.B1(n_3925),
.B2(n_3739),
.C(n_3970),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_L g4295 ( 
.A(n_4015),
.B(n_3715),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_4126),
.B(n_3925),
.Y(n_4296)
);

OA21x2_ASAP7_75t_L g4297 ( 
.A1(n_4018),
.A2(n_3739),
.B(n_3954),
.Y(n_4297)
);

NOR3xp33_ASAP7_75t_L g4298 ( 
.A(n_4080),
.B(n_4086),
.C(n_4212),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4144),
.B(n_3934),
.Y(n_4299)
);

AND2x2_ASAP7_75t_L g4300 ( 
.A(n_4035),
.B(n_657),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4145),
.B(n_661),
.Y(n_4301)
);

AND2x2_ASAP7_75t_L g4302 ( 
.A(n_4036),
.B(n_661),
.Y(n_4302)
);

NAND3xp33_ASAP7_75t_L g4303 ( 
.A(n_4154),
.B(n_3783),
.C(n_662),
.Y(n_4303)
);

NAND3xp33_ASAP7_75t_L g4304 ( 
.A(n_4154),
.B(n_4210),
.C(n_4049),
.Y(n_4304)
);

AND2x2_ASAP7_75t_L g4305 ( 
.A(n_4206),
.B(n_662),
.Y(n_4305)
);

OAI221xp5_ASAP7_75t_L g4306 ( 
.A1(n_4170),
.A2(n_3841),
.B1(n_3790),
.B2(n_4006),
.C(n_666),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_SL g4307 ( 
.A(n_4033),
.B(n_663),
.Y(n_4307)
);

AND2x2_ASAP7_75t_L g4308 ( 
.A(n_4206),
.B(n_664),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4167),
.B(n_824),
.Y(n_4309)
);

NAND4xp25_ASAP7_75t_SL g4310 ( 
.A(n_4113),
.B(n_667),
.C(n_664),
.D(n_665),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_4182),
.B(n_665),
.Y(n_4311)
);

NAND3xp33_ASAP7_75t_L g4312 ( 
.A(n_4242),
.B(n_4210),
.C(n_4177),
.Y(n_4312)
);

AND2x2_ASAP7_75t_SL g4313 ( 
.A(n_4297),
.B(n_4180),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4230),
.B(n_4075),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4233),
.Y(n_4315)
);

NAND3xp33_ASAP7_75t_L g4316 ( 
.A(n_4267),
.B(n_4179),
.C(n_4199),
.Y(n_4316)
);

INVx2_ASAP7_75t_L g4317 ( 
.A(n_4241),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4237),
.B(n_4089),
.Y(n_4318)
);

NOR3xp33_ASAP7_75t_L g4319 ( 
.A(n_4294),
.B(n_4306),
.C(n_4270),
.Y(n_4319)
);

INVx4_ASAP7_75t_SL g4320 ( 
.A(n_4265),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4215),
.B(n_4098),
.Y(n_4321)
);

NOR2xp33_ASAP7_75t_L g4322 ( 
.A(n_4295),
.B(n_4021),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4239),
.B(n_4047),
.Y(n_4323)
);

NOR3xp33_ASAP7_75t_L g4324 ( 
.A(n_4257),
.B(n_4212),
.C(n_4068),
.Y(n_4324)
);

OR2x2_ASAP7_75t_L g4325 ( 
.A(n_4216),
.B(n_4050),
.Y(n_4325)
);

OAI21xp5_ASAP7_75t_L g4326 ( 
.A1(n_4236),
.A2(n_4275),
.B(n_4287),
.Y(n_4326)
);

AOI22xp33_ASAP7_75t_L g4327 ( 
.A1(n_4298),
.A2(n_4193),
.B1(n_4087),
.B2(n_4025),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4226),
.Y(n_4328)
);

OR2x2_ASAP7_75t_L g4329 ( 
.A(n_4222),
.B(n_4052),
.Y(n_4329)
);

OAI21xp5_ASAP7_75t_L g4330 ( 
.A1(n_4236),
.A2(n_4186),
.B(n_4083),
.Y(n_4330)
);

INVxp67_ASAP7_75t_L g4331 ( 
.A(n_4252),
.Y(n_4331)
);

AO21x2_ASAP7_75t_L g4332 ( 
.A1(n_4283),
.A2(n_4018),
.B(n_4107),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_4225),
.B(n_4180),
.Y(n_4333)
);

AOI211xp5_ASAP7_75t_L g4334 ( 
.A1(n_4275),
.A2(n_4127),
.B(n_4117),
.C(n_4111),
.Y(n_4334)
);

NAND3xp33_ASAP7_75t_L g4335 ( 
.A(n_4248),
.B(n_4084),
.C(n_4105),
.Y(n_4335)
);

AOI22xp5_ASAP7_75t_L g4336 ( 
.A1(n_4280),
.A2(n_4100),
.B1(n_4108),
.B2(n_4194),
.Y(n_4336)
);

NOR3xp33_ASAP7_75t_SL g4337 ( 
.A(n_4269),
.B(n_4214),
.C(n_4142),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4218),
.B(n_4070),
.Y(n_4338)
);

NAND3xp33_ASAP7_75t_L g4339 ( 
.A(n_4304),
.B(n_4074),
.C(n_4071),
.Y(n_4339)
);

NOR3xp33_ASAP7_75t_L g4340 ( 
.A(n_4303),
.B(n_4259),
.C(n_4234),
.Y(n_4340)
);

OR2x2_ASAP7_75t_L g4341 ( 
.A(n_4217),
.B(n_4053),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4288),
.B(n_4076),
.Y(n_4342)
);

AOI22xp33_ASAP7_75t_L g4343 ( 
.A1(n_4273),
.A2(n_4173),
.B1(n_4203),
.B2(n_4109),
.Y(n_4343)
);

AOI22xp5_ASAP7_75t_L g4344 ( 
.A1(n_4287),
.A2(n_4196),
.B1(n_4174),
.B2(n_4082),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4223),
.B(n_4042),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4246),
.Y(n_4346)
);

NOR3xp33_ASAP7_75t_L g4347 ( 
.A(n_4292),
.B(n_4119),
.C(n_4128),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4249),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_4256),
.B(n_4208),
.Y(n_4349)
);

OAI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4293),
.A2(n_4081),
.B1(n_4064),
.B2(n_4205),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4255),
.Y(n_4351)
);

AND2x2_ASAP7_75t_L g4352 ( 
.A(n_4261),
.B(n_4139),
.Y(n_4352)
);

AND2x2_ASAP7_75t_L g4353 ( 
.A(n_4284),
.B(n_4178),
.Y(n_4353)
);

AOI221xp5_ASAP7_75t_L g4354 ( 
.A1(n_4273),
.A2(n_4160),
.B1(n_4166),
.B2(n_4149),
.C(n_4147),
.Y(n_4354)
);

OA21x2_ASAP7_75t_L g4355 ( 
.A1(n_4269),
.A2(n_4281),
.B(n_4272),
.Y(n_4355)
);

NAND3xp33_ASAP7_75t_L g4356 ( 
.A(n_4264),
.B(n_4058),
.C(n_4181),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4285),
.B(n_4200),
.Y(n_4357)
);

INVx1_ASAP7_75t_SL g4358 ( 
.A(n_4221),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4290),
.B(n_4054),
.Y(n_4359)
);

AO21x2_ASAP7_75t_L g4360 ( 
.A1(n_4305),
.A2(n_4155),
.B(n_4171),
.Y(n_4360)
);

NAND3xp33_ASAP7_75t_L g4361 ( 
.A(n_4264),
.B(n_4189),
.C(n_4184),
.Y(n_4361)
);

NOR3xp33_ASAP7_75t_L g4362 ( 
.A(n_4276),
.B(n_4132),
.C(n_4115),
.Y(n_4362)
);

NAND4xp75_ASAP7_75t_L g4363 ( 
.A(n_4297),
.B(n_4092),
.C(n_4187),
.D(n_4202),
.Y(n_4363)
);

NAND4xp75_ASAP7_75t_L g4364 ( 
.A(n_4262),
.B(n_4130),
.C(n_4175),
.D(n_4134),
.Y(n_4364)
);

OR2x2_ASAP7_75t_L g4365 ( 
.A(n_4219),
.B(n_668),
.Y(n_4365)
);

AND2x2_ASAP7_75t_L g4366 ( 
.A(n_4268),
.B(n_4204),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4286),
.B(n_4091),
.Y(n_4367)
);

NAND3xp33_ASAP7_75t_L g4368 ( 
.A(n_4276),
.B(n_4061),
.C(n_4095),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_4244),
.B(n_4067),
.Y(n_4369)
);

AO21x2_ASAP7_75t_L g4370 ( 
.A1(n_4308),
.A2(n_4103),
.B(n_4101),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4247),
.Y(n_4371)
);

OR2x2_ASAP7_75t_L g4372 ( 
.A(n_4220),
.B(n_670),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_4253),
.Y(n_4373)
);

NOR2x1_ASAP7_75t_L g4374 ( 
.A(n_4266),
.B(n_4060),
.Y(n_4374)
);

NAND3xp33_ASAP7_75t_L g4375 ( 
.A(n_4250),
.B(n_4238),
.C(n_4289),
.Y(n_4375)
);

NAND4xp25_ASAP7_75t_SL g4376 ( 
.A(n_4243),
.B(n_4088),
.C(n_4085),
.D(n_4063),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4279),
.B(n_4192),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4227),
.Y(n_4378)
);

OR2x2_ASAP7_75t_L g4379 ( 
.A(n_4240),
.B(n_671),
.Y(n_4379)
);

BUFx2_ASAP7_75t_L g4380 ( 
.A(n_4291),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_4228),
.Y(n_4381)
);

AOI22xp33_ASAP7_75t_L g4382 ( 
.A1(n_4310),
.A2(n_4079),
.B1(n_4077),
.B2(n_4066),
.Y(n_4382)
);

OR2x2_ASAP7_75t_L g4383 ( 
.A(n_4231),
.B(n_671),
.Y(n_4383)
);

AND2x2_ASAP7_75t_L g4384 ( 
.A(n_4254),
.B(n_4232),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_L g4385 ( 
.A(n_4271),
.B(n_4114),
.Y(n_4385)
);

AOI21xp5_ASAP7_75t_L g4386 ( 
.A1(n_4307),
.A2(n_4165),
.B(n_4055),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_4380),
.B(n_4296),
.Y(n_4387)
);

INVx1_ASAP7_75t_L g4388 ( 
.A(n_4346),
.Y(n_4388)
);

INVx2_ASAP7_75t_L g4389 ( 
.A(n_4351),
.Y(n_4389)
);

NAND4xp75_ASAP7_75t_L g4390 ( 
.A(n_4326),
.B(n_4278),
.C(n_4302),
.D(n_4300),
.Y(n_4390)
);

INVx1_ASAP7_75t_L g4391 ( 
.A(n_4346),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4328),
.B(n_4235),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4328),
.B(n_4258),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4381),
.Y(n_4394)
);

XOR2x2_ASAP7_75t_L g4395 ( 
.A(n_4358),
.B(n_4282),
.Y(n_4395)
);

NAND3xp33_ASAP7_75t_SL g4396 ( 
.A(n_4319),
.B(n_4266),
.C(n_4224),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4381),
.Y(n_4397)
);

XOR2x2_ASAP7_75t_L g4398 ( 
.A(n_4322),
.B(n_4299),
.Y(n_4398)
);

NOR4xp25_ASAP7_75t_L g4399 ( 
.A(n_4335),
.B(n_4251),
.C(n_4309),
.D(n_4301),
.Y(n_4399)
);

INVx1_ASAP7_75t_SL g4400 ( 
.A(n_4329),
.Y(n_4400)
);

INVx1_ASAP7_75t_L g4401 ( 
.A(n_4371),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4373),
.Y(n_4402)
);

INVx4_ASAP7_75t_L g4403 ( 
.A(n_4332),
.Y(n_4403)
);

INVx2_ASAP7_75t_SL g4404 ( 
.A(n_4317),
.Y(n_4404)
);

AND2x2_ASAP7_75t_SL g4405 ( 
.A(n_4355),
.B(n_4263),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4315),
.Y(n_4406)
);

AND2x2_ASAP7_75t_L g4407 ( 
.A(n_4348),
.B(n_4323),
.Y(n_4407)
);

OR2x2_ASAP7_75t_L g4408 ( 
.A(n_4315),
.B(n_4274),
.Y(n_4408)
);

NOR3xp33_ASAP7_75t_L g4409 ( 
.A(n_4375),
.B(n_4245),
.C(n_4311),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4378),
.Y(n_4410)
);

NAND4xp75_ASAP7_75t_L g4411 ( 
.A(n_4374),
.B(n_4355),
.C(n_4313),
.D(n_4330),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4325),
.Y(n_4412)
);

NAND4xp75_ASAP7_75t_L g4413 ( 
.A(n_4344),
.B(n_4337),
.C(n_4336),
.D(n_4385),
.Y(n_4413)
);

INVx2_ASAP7_75t_L g4414 ( 
.A(n_4333),
.Y(n_4414)
);

CKINVDCx20_ASAP7_75t_R g4415 ( 
.A(n_4331),
.Y(n_4415)
);

NAND4xp75_ASAP7_75t_SL g4416 ( 
.A(n_4363),
.B(n_4229),
.C(n_4110),
.D(n_4106),
.Y(n_4416)
);

NAND4xp75_ASAP7_75t_L g4417 ( 
.A(n_4367),
.B(n_4260),
.C(n_4277),
.D(n_4229),
.Y(n_4417)
);

XOR2x2_ASAP7_75t_L g4418 ( 
.A(n_4340),
.B(n_4141),
.Y(n_4418)
);

AND2x4_ASAP7_75t_L g4419 ( 
.A(n_4320),
.B(n_4156),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4384),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4345),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4314),
.Y(n_4422)
);

XOR2x2_ASAP7_75t_L g4423 ( 
.A(n_4316),
.B(n_4152),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_4318),
.B(n_4122),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4332),
.B(n_4123),
.Y(n_4425)
);

INVx2_ASAP7_75t_L g4426 ( 
.A(n_4341),
.Y(n_4426)
);

NOR2x1_ASAP7_75t_L g4427 ( 
.A(n_4372),
.B(n_672),
.Y(n_4427)
);

NAND4xp75_ASAP7_75t_SL g4428 ( 
.A(n_4359),
.B(n_677),
.C(n_674),
.D(n_675),
.Y(n_4428)
);

NAND3xp33_ASAP7_75t_L g4429 ( 
.A(n_4324),
.B(n_4062),
.C(n_4078),
.Y(n_4429)
);

INVx2_ASAP7_75t_L g4430 ( 
.A(n_4338),
.Y(n_4430)
);

AND2x4_ASAP7_75t_L g4431 ( 
.A(n_4320),
.B(n_4116),
.Y(n_4431)
);

CKINVDCx20_ASAP7_75t_R g4432 ( 
.A(n_4321),
.Y(n_4432)
);

NOR3xp33_ASAP7_75t_L g4433 ( 
.A(n_4339),
.B(n_678),
.C(n_680),
.Y(n_4433)
);

NAND4xp75_ASAP7_75t_L g4434 ( 
.A(n_4353),
.B(n_4140),
.C(n_4136),
.D(n_4151),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_4342),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4327),
.B(n_4349),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4365),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4383),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4357),
.B(n_4153),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4352),
.Y(n_4440)
);

BUFx2_ASAP7_75t_L g4441 ( 
.A(n_4379),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4377),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4369),
.B(n_4135),
.Y(n_4443)
);

XNOR2xp5_ASAP7_75t_L g4444 ( 
.A(n_4350),
.B(n_678),
.Y(n_4444)
);

NOR3xp33_ASAP7_75t_L g4445 ( 
.A(n_4368),
.B(n_681),
.C(n_682),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4366),
.B(n_4370),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4370),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4360),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4343),
.B(n_681),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4360),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4362),
.B(n_683),
.Y(n_4451)
);

XOR2x2_ASAP7_75t_L g4452 ( 
.A(n_4413),
.B(n_4361),
.Y(n_4452)
);

INVx1_ASAP7_75t_L g4453 ( 
.A(n_4388),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4446),
.B(n_4356),
.Y(n_4454)
);

OR2x2_ASAP7_75t_L g4455 ( 
.A(n_4400),
.B(n_4312),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4404),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_4400),
.B(n_4347),
.Y(n_4457)
);

XNOR2xp5_ASAP7_75t_L g4458 ( 
.A(n_4395),
.B(n_4334),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4426),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_4391),
.Y(n_4460)
);

INVx1_ASAP7_75t_L g4461 ( 
.A(n_4394),
.Y(n_4461)
);

INVxp67_ASAP7_75t_L g4462 ( 
.A(n_4396),
.Y(n_4462)
);

CKINVDCx16_ASAP7_75t_R g4463 ( 
.A(n_4415),
.Y(n_4463)
);

XNOR2xp5_ASAP7_75t_L g4464 ( 
.A(n_4398),
.B(n_4364),
.Y(n_4464)
);

INVx2_ASAP7_75t_L g4465 ( 
.A(n_4406),
.Y(n_4465)
);

INVx1_ASAP7_75t_SL g4466 ( 
.A(n_4432),
.Y(n_4466)
);

HB1xp67_ASAP7_75t_L g4467 ( 
.A(n_4412),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4389),
.Y(n_4468)
);

HB1xp67_ASAP7_75t_L g4469 ( 
.A(n_4397),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4401),
.Y(n_4470)
);

BUFx2_ASAP7_75t_L g4471 ( 
.A(n_4402),
.Y(n_4471)
);

XNOR2xp5_ASAP7_75t_L g4472 ( 
.A(n_4444),
.B(n_4354),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4410),
.Y(n_4473)
);

XOR2x2_ASAP7_75t_L g4474 ( 
.A(n_4416),
.B(n_4386),
.Y(n_4474)
);

OA22x2_ASAP7_75t_L g4475 ( 
.A1(n_4403),
.A2(n_4376),
.B1(n_4382),
.B2(n_685),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4393),
.Y(n_4476)
);

INVx1_ASAP7_75t_SL g4477 ( 
.A(n_4387),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4414),
.Y(n_4478)
);

XOR2x2_ASAP7_75t_L g4479 ( 
.A(n_4411),
.B(n_683),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4408),
.Y(n_4480)
);

INVx1_ASAP7_75t_SL g4481 ( 
.A(n_4441),
.Y(n_4481)
);

XNOR2xp5_ASAP7_75t_L g4482 ( 
.A(n_4390),
.B(n_684),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4393),
.Y(n_4483)
);

XOR2x2_ASAP7_75t_L g4484 ( 
.A(n_4417),
.B(n_684),
.Y(n_4484)
);

XOR2x2_ASAP7_75t_L g4485 ( 
.A(n_4436),
.B(n_686),
.Y(n_4485)
);

INVx1_ASAP7_75t_L g4486 ( 
.A(n_4392),
.Y(n_4486)
);

INVxp67_ASAP7_75t_L g4487 ( 
.A(n_4451),
.Y(n_4487)
);

XOR2x2_ASAP7_75t_L g4488 ( 
.A(n_4418),
.B(n_687),
.Y(n_4488)
);

INVx3_ASAP7_75t_L g4489 ( 
.A(n_4403),
.Y(n_4489)
);

OR2x6_ASAP7_75t_L g4490 ( 
.A(n_4427),
.B(n_4419),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4430),
.B(n_4435),
.Y(n_4491)
);

AND2x2_ASAP7_75t_L g4492 ( 
.A(n_4442),
.B(n_687),
.Y(n_4492)
);

AOI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_4475),
.A2(n_4405),
.B1(n_4409),
.B2(n_4399),
.Y(n_4493)
);

INVx1_ASAP7_75t_L g4494 ( 
.A(n_4467),
.Y(n_4494)
);

OA22x2_ASAP7_75t_L g4495 ( 
.A1(n_4462),
.A2(n_4448),
.B1(n_4447),
.B2(n_4450),
.Y(n_4495)
);

INVx1_ASAP7_75t_SL g4496 ( 
.A(n_4463),
.Y(n_4496)
);

AOI22xp5_ASAP7_75t_L g4497 ( 
.A1(n_4452),
.A2(n_4399),
.B1(n_4423),
.B2(n_4425),
.Y(n_4497)
);

AOI22xp5_ASAP7_75t_L g4498 ( 
.A1(n_4458),
.A2(n_4425),
.B1(n_4431),
.B2(n_4419),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4469),
.Y(n_4499)
);

INVx3_ASAP7_75t_L g4500 ( 
.A(n_4471),
.Y(n_4500)
);

OA22x2_ASAP7_75t_L g4501 ( 
.A1(n_4490),
.A2(n_4431),
.B1(n_4422),
.B2(n_4438),
.Y(n_4501)
);

OAI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4490),
.A2(n_4421),
.B1(n_4440),
.B2(n_4420),
.Y(n_4502)
);

AO22x2_ASAP7_75t_L g4503 ( 
.A1(n_4455),
.A2(n_4454),
.B1(n_4481),
.B2(n_4489),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4480),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4473),
.Y(n_4505)
);

XOR2x2_ASAP7_75t_L g4506 ( 
.A(n_4464),
.B(n_4474),
.Y(n_4506)
);

NOR2x1_ASAP7_75t_L g4507 ( 
.A(n_4489),
.B(n_4427),
.Y(n_4507)
);

XOR2x2_ASAP7_75t_L g4508 ( 
.A(n_4488),
.B(n_4434),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_4473),
.Y(n_4509)
);

OAI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_4457),
.A2(n_4437),
.B1(n_4424),
.B2(n_4392),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4468),
.Y(n_4511)
);

AOI22xp5_ASAP7_75t_L g4512 ( 
.A1(n_4479),
.A2(n_4429),
.B1(n_4443),
.B2(n_4445),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_SL g4513 ( 
.A(n_4466),
.B(n_4484),
.Y(n_4513)
);

OA22x2_ASAP7_75t_L g4514 ( 
.A1(n_4472),
.A2(n_4449),
.B1(n_4424),
.B2(n_4439),
.Y(n_4514)
);

INVx1_ASAP7_75t_L g4515 ( 
.A(n_4461),
.Y(n_4515)
);

INVx2_ASAP7_75t_L g4516 ( 
.A(n_4478),
.Y(n_4516)
);

INVx2_ASAP7_75t_SL g4517 ( 
.A(n_4456),
.Y(n_4517)
);

INVx1_ASAP7_75t_L g4518 ( 
.A(n_4460),
.Y(n_4518)
);

INVxp67_ASAP7_75t_SL g4519 ( 
.A(n_4482),
.Y(n_4519)
);

AO22x1_ASAP7_75t_L g4520 ( 
.A1(n_4487),
.A2(n_4433),
.B1(n_4407),
.B2(n_4428),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4486),
.Y(n_4521)
);

OA22x2_ASAP7_75t_L g4522 ( 
.A1(n_4477),
.A2(n_4429),
.B1(n_689),
.B2(n_690),
.Y(n_4522)
);

AOI22xp5_ASAP7_75t_L g4523 ( 
.A1(n_4485),
.A2(n_688),
.B1(n_689),
.B2(n_690),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_SL g4524 ( 
.A(n_4492),
.B(n_688),
.Y(n_4524)
);

OA22x2_ASAP7_75t_L g4525 ( 
.A1(n_4476),
.A2(n_4483),
.B1(n_4486),
.B2(n_4459),
.Y(n_4525)
);

BUFx2_ASAP7_75t_L g4526 ( 
.A(n_4476),
.Y(n_4526)
);

INVx2_ASAP7_75t_L g4527 ( 
.A(n_4491),
.Y(n_4527)
);

XNOR2xp5_ASAP7_75t_L g4528 ( 
.A(n_4483),
.B(n_691),
.Y(n_4528)
);

INVx3_ASAP7_75t_L g4529 ( 
.A(n_4465),
.Y(n_4529)
);

OAI22x1_ASAP7_75t_L g4530 ( 
.A1(n_4470),
.A2(n_691),
.B1(n_692),
.B2(n_695),
.Y(n_4530)
);

OA22x2_ASAP7_75t_L g4531 ( 
.A1(n_4470),
.A2(n_696),
.B1(n_697),
.B2(n_698),
.Y(n_4531)
);

AOI22x1_ASAP7_75t_L g4532 ( 
.A1(n_4453),
.A2(n_696),
.B1(n_697),
.B2(n_698),
.Y(n_4532)
);

XOR2x2_ASAP7_75t_L g4533 ( 
.A(n_4453),
.B(n_699),
.Y(n_4533)
);

HB1xp67_ASAP7_75t_L g4534 ( 
.A(n_4471),
.Y(n_4534)
);

AOI22x1_ASAP7_75t_L g4535 ( 
.A1(n_4458),
.A2(n_700),
.B1(n_701),
.B2(n_702),
.Y(n_4535)
);

OAI22x1_ASAP7_75t_L g4536 ( 
.A1(n_4458),
.A2(n_701),
.B1(n_705),
.B2(n_706),
.Y(n_4536)
);

XOR2x2_ASAP7_75t_L g4537 ( 
.A(n_4452),
.B(n_705),
.Y(n_4537)
);

AOI322xp5_ASAP7_75t_L g4538 ( 
.A1(n_4497),
.A2(n_823),
.A3(n_707),
.B1(n_708),
.B2(n_709),
.C1(n_711),
.C2(n_712),
.Y(n_4538)
);

INVx2_ASAP7_75t_L g4539 ( 
.A(n_4500),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4494),
.Y(n_4540)
);

HB1xp67_ASAP7_75t_L g4541 ( 
.A(n_4526),
.Y(n_4541)
);

INVx2_ASAP7_75t_SL g4542 ( 
.A(n_4496),
.Y(n_4542)
);

HB1xp67_ASAP7_75t_L g4543 ( 
.A(n_4526),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_4534),
.Y(n_4544)
);

INVx2_ASAP7_75t_L g4545 ( 
.A(n_4527),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4499),
.Y(n_4546)
);

OA22x2_ASAP7_75t_L g4547 ( 
.A1(n_4493),
.A2(n_706),
.B1(n_707),
.B2(n_708),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4504),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4515),
.Y(n_4549)
);

INVx2_ASAP7_75t_L g4550 ( 
.A(n_4529),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4518),
.Y(n_4551)
);

INVx2_ASAP7_75t_L g4552 ( 
.A(n_4511),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_4505),
.Y(n_4553)
);

HB1xp67_ASAP7_75t_L g4554 ( 
.A(n_4503),
.Y(n_4554)
);

INVx2_ASAP7_75t_L g4555 ( 
.A(n_4516),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4509),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4521),
.Y(n_4557)
);

HB1xp67_ASAP7_75t_L g4558 ( 
.A(n_4503),
.Y(n_4558)
);

NAND2x1_ASAP7_75t_SL g4559 ( 
.A(n_4507),
.B(n_820),
.Y(n_4559)
);

INVx5_ASAP7_75t_L g4560 ( 
.A(n_4508),
.Y(n_4560)
);

INVxp67_ASAP7_75t_SL g4561 ( 
.A(n_4522),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4517),
.Y(n_4562)
);

INVx1_ASAP7_75t_L g4563 ( 
.A(n_4525),
.Y(n_4563)
);

INVx2_ASAP7_75t_L g4564 ( 
.A(n_4531),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4510),
.Y(n_4565)
);

HB1xp67_ASAP7_75t_L g4566 ( 
.A(n_4513),
.Y(n_4566)
);

INVx2_ASAP7_75t_L g4567 ( 
.A(n_4530),
.Y(n_4567)
);

INVx1_ASAP7_75t_L g4568 ( 
.A(n_4541),
.Y(n_4568)
);

AND4x1_ASAP7_75t_L g4569 ( 
.A(n_4562),
.B(n_4512),
.C(n_4498),
.D(n_4523),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4541),
.Y(n_4570)
);

AOI22xp5_ASAP7_75t_L g4571 ( 
.A1(n_4542),
.A2(n_4514),
.B1(n_4519),
.B2(n_4506),
.Y(n_4571)
);

INVx2_ASAP7_75t_L g4572 ( 
.A(n_4539),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4543),
.Y(n_4573)
);

AO22x1_ASAP7_75t_L g4574 ( 
.A1(n_4561),
.A2(n_4501),
.B1(n_4502),
.B2(n_4528),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4543),
.Y(n_4575)
);

INVx5_ASAP7_75t_L g4576 ( 
.A(n_4560),
.Y(n_4576)
);

AOI22xp5_ASAP7_75t_L g4577 ( 
.A1(n_4561),
.A2(n_4566),
.B1(n_4564),
.B2(n_4565),
.Y(n_4577)
);

INVx1_ASAP7_75t_SL g4578 ( 
.A(n_4559),
.Y(n_4578)
);

AOI221xp5_ASAP7_75t_L g4579 ( 
.A1(n_4566),
.A2(n_4536),
.B1(n_4528),
.B2(n_4520),
.C(n_4524),
.Y(n_4579)
);

INVx1_ASAP7_75t_L g4580 ( 
.A(n_4554),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4554),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4558),
.Y(n_4582)
);

INVx2_ASAP7_75t_L g4583 ( 
.A(n_4544),
.Y(n_4583)
);

OA22x2_ASAP7_75t_L g4584 ( 
.A1(n_4558),
.A2(n_4537),
.B1(n_4533),
.B2(n_4495),
.Y(n_4584)
);

OAI322xp33_ASAP7_75t_L g4585 ( 
.A1(n_4563),
.A2(n_4564),
.A3(n_4547),
.B1(n_4567),
.B2(n_4546),
.C1(n_4540),
.C2(n_4548),
.Y(n_4585)
);

OAI222xp33_ASAP7_75t_L g4586 ( 
.A1(n_4560),
.A2(n_4535),
.B1(n_4532),
.B2(n_712),
.C1(n_713),
.C2(n_715),
.Y(n_4586)
);

OA22x2_ASAP7_75t_L g4587 ( 
.A1(n_4550),
.A2(n_709),
.B1(n_711),
.B2(n_715),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4549),
.Y(n_4588)
);

INVx1_ASAP7_75t_SL g4589 ( 
.A(n_4560),
.Y(n_4589)
);

AOI221xp5_ASAP7_75t_L g4590 ( 
.A1(n_4560),
.A2(n_716),
.B1(n_717),
.B2(n_718),
.C(n_719),
.Y(n_4590)
);

INVxp33_ASAP7_75t_SL g4591 ( 
.A(n_4589),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4568),
.Y(n_4592)
);

AOI22xp33_ASAP7_75t_SL g4593 ( 
.A1(n_4584),
.A2(n_4547),
.B1(n_4545),
.B2(n_4551),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4570),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4573),
.Y(n_4595)
);

OAI22x1_ASAP7_75t_L g4596 ( 
.A1(n_4571),
.A2(n_4557),
.B1(n_4556),
.B2(n_4553),
.Y(n_4596)
);

AOI22x1_ASAP7_75t_L g4597 ( 
.A1(n_4578),
.A2(n_4555),
.B1(n_4552),
.B2(n_4538),
.Y(n_4597)
);

HB1xp67_ASAP7_75t_L g4598 ( 
.A(n_4575),
.Y(n_4598)
);

AOI22x1_ASAP7_75t_L g4599 ( 
.A1(n_4580),
.A2(n_816),
.B1(n_717),
.B2(n_718),
.Y(n_4599)
);

AOI311xp33_ASAP7_75t_L g4600 ( 
.A1(n_4581),
.A2(n_716),
.A3(n_719),
.B(n_720),
.C(n_721),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4583),
.Y(n_4601)
);

AOI22xp5_ASAP7_75t_L g4602 ( 
.A1(n_4579),
.A2(n_722),
.B1(n_723),
.B2(n_724),
.Y(n_4602)
);

AOI22xp5_ASAP7_75t_L g4603 ( 
.A1(n_4574),
.A2(n_722),
.B1(n_723),
.B2(n_725),
.Y(n_4603)
);

AND4x1_ASAP7_75t_L g4604 ( 
.A(n_4577),
.B(n_725),
.C(n_726),
.D(n_727),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4572),
.Y(n_4605)
);

O2A1O1Ixp5_ASAP7_75t_SL g4606 ( 
.A1(n_4582),
.A2(n_4576),
.B(n_4588),
.C(n_4585),
.Y(n_4606)
);

INVx1_ASAP7_75t_L g4607 ( 
.A(n_4587),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4576),
.Y(n_4608)
);

OA22x2_ASAP7_75t_L g4609 ( 
.A1(n_4569),
.A2(n_726),
.B1(n_727),
.B2(n_728),
.Y(n_4609)
);

HB1xp67_ASAP7_75t_L g4610 ( 
.A(n_4576),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4590),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4598),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4605),
.Y(n_4613)
);

AOI31xp33_ASAP7_75t_L g4614 ( 
.A1(n_4593),
.A2(n_4586),
.A3(n_730),
.B(n_731),
.Y(n_4614)
);

AO22x1_ASAP7_75t_L g4615 ( 
.A1(n_4607),
.A2(n_728),
.B1(n_730),
.B2(n_731),
.Y(n_4615)
);

NOR2x1_ASAP7_75t_L g4616 ( 
.A(n_4608),
.B(n_733),
.Y(n_4616)
);

NOR4xp25_ASAP7_75t_L g4617 ( 
.A(n_4592),
.B(n_733),
.C(n_734),
.D(n_735),
.Y(n_4617)
);

AOI22xp5_ASAP7_75t_L g4618 ( 
.A1(n_4603),
.A2(n_4591),
.B1(n_4609),
.B2(n_4602),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4610),
.Y(n_4619)
);

NOR2xp33_ASAP7_75t_L g4620 ( 
.A(n_4604),
.B(n_734),
.Y(n_4620)
);

A2O1A1Ixp33_ASAP7_75t_SL g4621 ( 
.A1(n_4594),
.A2(n_735),
.B(n_736),
.C(n_737),
.Y(n_4621)
);

NOR4xp25_ASAP7_75t_L g4622 ( 
.A(n_4595),
.B(n_736),
.C(n_737),
.D(n_738),
.Y(n_4622)
);

NOR3xp33_ASAP7_75t_L g4623 ( 
.A(n_4611),
.B(n_816),
.C(n_738),
.Y(n_4623)
);

INVx1_ASAP7_75t_L g4624 ( 
.A(n_4601),
.Y(n_4624)
);

OA22x2_ASAP7_75t_L g4625 ( 
.A1(n_4596),
.A2(n_813),
.B1(n_741),
.B2(n_742),
.Y(n_4625)
);

INVxp67_ASAP7_75t_SL g4626 ( 
.A(n_4619),
.Y(n_4626)
);

NOR2x1_ASAP7_75t_L g4627 ( 
.A(n_4616),
.B(n_4606),
.Y(n_4627)
);

NAND2xp5_ASAP7_75t_SL g4628 ( 
.A(n_4614),
.B(n_4597),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4615),
.B(n_4599),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4613),
.Y(n_4630)
);

AOI22xp5_ASAP7_75t_L g4631 ( 
.A1(n_4618),
.A2(n_4600),
.B1(n_743),
.B2(n_744),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4624),
.Y(n_4632)
);

NOR2x1_ASAP7_75t_L g4633 ( 
.A(n_4612),
.B(n_4600),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4625),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4620),
.Y(n_4635)
);

OA22x2_ASAP7_75t_L g4636 ( 
.A1(n_4623),
.A2(n_740),
.B1(n_744),
.B2(n_745),
.Y(n_4636)
);

INVx1_ASAP7_75t_L g4637 ( 
.A(n_4626),
.Y(n_4637)
);

OR2x2_ASAP7_75t_L g4638 ( 
.A(n_4634),
.B(n_4617),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4630),
.Y(n_4639)
);

AO22x1_ASAP7_75t_L g4640 ( 
.A1(n_4627),
.A2(n_4622),
.B1(n_4621),
.B2(n_748),
.Y(n_4640)
);

INVxp67_ASAP7_75t_L g4641 ( 
.A(n_4633),
.Y(n_4641)
);

NAND2x1_ASAP7_75t_L g4642 ( 
.A(n_4632),
.B(n_740),
.Y(n_4642)
);

AOI22xp5_ASAP7_75t_L g4643 ( 
.A1(n_4628),
.A2(n_745),
.B1(n_748),
.B2(n_749),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4639),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4637),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4643),
.Y(n_4646)
);

INVxp67_ASAP7_75t_SL g4647 ( 
.A(n_4641),
.Y(n_4647)
);

INVx1_ASAP7_75t_L g4648 ( 
.A(n_4642),
.Y(n_4648)
);

AOI22xp5_ASAP7_75t_L g4649 ( 
.A1(n_4647),
.A2(n_4631),
.B1(n_4629),
.B2(n_4635),
.Y(n_4649)
);

OAI22x1_ASAP7_75t_L g4650 ( 
.A1(n_4648),
.A2(n_4638),
.B1(n_4640),
.B2(n_4636),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4650),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4649),
.Y(n_4652)
);

AOI22xp33_ASAP7_75t_SL g4653 ( 
.A1(n_4652),
.A2(n_4646),
.B1(n_4645),
.B2(n_4644),
.Y(n_4653)
);

BUFx3_ASAP7_75t_L g4654 ( 
.A(n_4653),
.Y(n_4654)
);

AOI22xp5_ASAP7_75t_SL g4655 ( 
.A1(n_4654),
.A2(n_4651),
.B1(n_751),
.B2(n_752),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4655),
.Y(n_4656)
);

AOI221xp5_ASAP7_75t_L g4657 ( 
.A1(n_4656),
.A2(n_750),
.B1(n_752),
.B2(n_753),
.C(n_754),
.Y(n_4657)
);

AOI211xp5_ASAP7_75t_L g4658 ( 
.A1(n_4657),
.A2(n_753),
.B(n_754),
.C(n_755),
.Y(n_4658)
);


endmodule