module fake_jpeg_9485_n_120 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_120);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_120;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_41),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_4),
.B1(n_7),
.B2(n_45),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_61),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_71),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_1),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_3),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_94),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_50),
.B1(n_55),
.B2(n_53),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_67),
.A2(n_51),
.B1(n_58),
.B2(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_87),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_48),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_48),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_24),
.C(n_28),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_30),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_13),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_23),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_104),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_101),
.B1(n_77),
.B2(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_96),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_101),
.B1(n_76),
.B2(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_102),
.C(n_94),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_31),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_105),
.B1(n_99),
.B2(n_89),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_103),
.A3(n_34),
.B1(n_35),
.B2(n_37),
.C1(n_38),
.C2(n_40),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_100),
.C(n_42),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_32),
.C(n_43),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_44),
.B1(n_74),
.B2(n_82),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_78),
.Y(n_120)
);


endmodule