module real_jpeg_29311_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_335, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_335;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_0),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_0),
.A2(n_148),
.B(n_161),
.Y(n_160)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_1),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_31),
.B1(n_33),
.B2(n_133),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_133),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_1),
.A2(n_63),
.B1(n_65),
.B2(n_133),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_3),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_33),
.Y(n_173)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_33),
.B(n_173),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_131),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_3),
.A2(n_11),
.B(n_63),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_3),
.B(n_89),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_3),
.A2(n_110),
.B1(n_116),
.B2(n_225),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_5),
.A2(n_31),
.B1(n_33),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_5),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_126),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_126),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_5),
.A2(n_63),
.B1(n_65),
.B2(n_126),
.Y(n_217)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_37),
.B1(n_63),
.B2(n_65),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_7),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_8),
.A2(n_52),
.B1(n_63),
.B2(n_65),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_55),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_55),
.B1(n_63),
.B2(n_65),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_10),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_13),
.A2(n_31),
.B1(n_33),
.B2(n_50),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_14),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_128),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_14),
.A2(n_63),
.B1(n_65),
.B2(n_128),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_128),
.Y(n_265)
);

INVx11_ASAP7_75t_SL g64 ( 
.A(n_15),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_75),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_70),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_23),
.A2(n_38),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_23),
.A2(n_38),
.B1(n_139),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_23),
.A2(n_265),
.B(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_24),
.A2(n_30),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_24),
.A2(n_86),
.B(n_285),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_25),
.B(n_33),
.Y(n_145)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g130 ( 
.A(n_27),
.B(n_131),
.CON(n_130),
.SN(n_130)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_29),
.A2(n_31),
.B1(n_130),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_30),
.B(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_31),
.A2(n_45),
.A3(n_48),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_34),
.A2(n_38),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_38),
.B(n_131),
.Y(n_158)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_58),
.B2(n_69),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_58),
.C(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_43),
.A2(n_77),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_51),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_44),
.A2(n_56),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_44),
.A2(n_56),
.B1(n_125),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_44),
.A2(n_56),
.B1(n_157),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_44),
.A2(n_56),
.B1(n_79),
.B2(n_304),
.Y(n_303)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g174 ( 
.A(n_46),
.B(n_49),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_46),
.A2(n_61),
.B(n_131),
.C(n_201),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_51),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_53),
.A2(n_89),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_58),
.A2(n_69),
.B1(n_76),
.B2(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_67),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_59),
.A2(n_67),
.B(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_59),
.A2(n_62),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_59),
.A2(n_181),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_59),
.A2(n_62),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_59),
.A2(n_62),
.B1(n_180),
.B2(n_199),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_59),
.A2(n_62),
.B1(n_105),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_59),
.A2(n_121),
.B(n_258),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_62),
.B(n_131),
.Y(n_223)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_65),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_68),
.B(n_122),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.C(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_71),
.A2(n_318),
.B1(n_320),
.B2(n_321),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_71),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_75),
.B(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_76),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_77),
.A2(n_80),
.B(n_90),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_314),
.A3(n_326),
.B1(n_332),
.B2(n_333),
.C(n_335),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_296),
.B(n_313),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_271),
.B(n_295),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_162),
.B(n_248),
.C(n_270),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_149),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_101),
.B(n_149),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_134),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_118),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_103),
.B(n_118),
.C(n_134),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_104),
.B(n_109),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_106),
.B(n_191),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B(n_114),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_113),
.B1(n_116),
.B2(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_117),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_110),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_110),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_110),
.A2(n_212),
.B1(n_217),
.B2(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_110),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_111),
.B(n_131),
.Y(n_229)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_115),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_129),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_143),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_136),
.B(n_141),
.C(n_143),
.Y(n_268)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_150),
.A2(n_151),
.B1(n_243),
.B2(n_245),
.Y(n_242)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_156),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_186),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_158),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_161),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_247),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_240),
.B(n_246),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_192),
.B(n_239),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_182),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_182),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.C(n_178),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_167),
.A2(n_168),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_170),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_211),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_179),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_183),
.B(n_189),
.C(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_233),
.B(n_238),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_213),
.B(n_232),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_202),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_195),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_207),
.C(n_208),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_210),
.B(n_256),
.Y(n_255)
);

INVx5_ASAP7_75t_SL g290 ( 
.A(n_211),
.Y(n_290)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_221),
.B(n_231),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_215),
.B(n_219),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_226),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_250),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_268),
.B2(n_269),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_259),
.B2(n_260),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_260),
.C(n_269),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_263),
.C(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_273),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_294),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_286),
.B2(n_287),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_287),
.C(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_280),
.C(n_282),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_283),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_281),
.Y(n_304)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_288),
.A2(n_289),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_292),
.Y(n_307)
);

AOI21xp33_ASAP7_75t_L g323 ( 
.A1(n_289),
.A2(n_307),
.B(n_310),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_300),
.B1(n_311),
.B2(n_312),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_306),
.C(n_312),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B(n_305),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_316),
.C(n_322),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_305),
.A2(n_316),
.B1(n_317),
.B2(n_331),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_324),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_324),
.Y(n_333)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_318),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_323),
.B1(n_329),
.B2(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule