module fake_jpeg_18486_n_32 (n_3, n_2, n_1, n_0, n_4, n_5, n_32);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_32;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_2),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_8),
.B1(n_7),
.B2(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_7),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_19),
.B(n_8),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_22),
.C(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_17),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_15),
.C(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_19),
.C(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_15),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.C(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_11),
.Y(n_28)
);

OAI311xp33_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_10),
.A3(n_1),
.B1(n_3),
.C1(n_5),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_9),
.A3(n_12),
.B1(n_5),
.B2(n_3),
.C1(n_10),
.C2(n_0),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_9),
.B1(n_12),
.B2(n_0),
.Y(n_32)
);


endmodule