module fake_jpeg_4802_n_160 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_160);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_15),
.B1(n_14),
.B2(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_23),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_15),
.B1(n_21),
.B2(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_52),
.B1(n_36),
.B2(n_26),
.Y(n_73)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_18),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_17),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_58),
.B(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_15),
.B1(n_21),
.B2(n_27),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_14),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_29),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_57),
.Y(n_76)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_29),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_36),
.B1(n_38),
.B2(n_44),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_41),
.Y(n_80)
);

OAI22x1_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_38),
.B1(n_27),
.B2(n_36),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_51),
.B1(n_50),
.B2(n_57),
.Y(n_96)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_70),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_58),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_78),
.B1(n_51),
.B2(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_24),
.B1(n_22),
.B2(n_31),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_87),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_49),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_92),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_60),
.A2(n_40),
.B1(n_52),
.B2(n_48),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_96),
.B1(n_74),
.B2(n_63),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_40),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_46),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_65),
.C(n_42),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_43),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_51),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_31),
.B1(n_22),
.B2(n_42),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_104),
.C(n_98),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_72),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_111),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_61),
.C(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_108),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_112),
.B1(n_114),
.B2(n_99),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_33),
.CI(n_14),
.CON(n_107),
.SN(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_33),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_83),
.A2(n_66),
.B(n_33),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_90),
.B(n_95),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_33),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_31),
.B1(n_62),
.B2(n_22),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_81),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_25),
.B1(n_14),
.B2(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_119),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_89),
.B(n_93),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_96),
.C(n_85),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_120),
.B(n_125),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_111),
.B1(n_101),
.B2(n_112),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_121),
.A2(n_103),
.B1(n_114),
.B2(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_97),
.B(n_84),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_25),
.C(n_1),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_4),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_107),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_126),
.B(n_25),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_119),
.Y(n_140)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_117),
.B(n_116),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_141),
.B(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_121),
.C(n_124),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_143),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_118),
.B(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_144),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_148),
.B(n_149),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_128),
.Y(n_148)
);

NOR2x1_ASAP7_75t_R g149 ( 
.A(n_143),
.B(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_132),
.C(n_135),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_150),
.B1(n_147),
.B2(n_146),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_151),
.B(n_4),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_10),
.B(n_11),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_155),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_157),
.C(n_11),
.Y(n_160)
);


endmodule