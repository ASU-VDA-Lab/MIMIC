module real_aes_16921_n_14 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_14);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_14;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_46;
wire n_25;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_0), .B(n_5), .C(n_20), .Y(n_19) );
NOR5xp2_ASAP7_75t_SL g17 ( .A(n_1), .B(n_10), .C(n_18), .D(n_22), .E(n_23), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_1), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_2), .B(n_25), .Y(n_24) );
NAND2xp33_ASAP7_75t_R g29 ( .A(n_2), .B(n_4), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_2), .Y(n_42) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_3), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_4), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_4), .B(n_42), .Y(n_41) );
AOI221xp5_ASAP7_75t_SL g14 ( .A1(n_6), .A2(n_8), .B1(n_15), .B2(n_26), .C(n_30), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_7), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g46 ( .A(n_9), .Y(n_46) );
CKINVDCx5p33_ASAP7_75t_R g38 ( .A(n_10), .Y(n_38) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_11), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_12), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_13), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_16), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g16 ( .A(n_17), .B(n_24), .Y(n_16) );
NAND2xp33_ASAP7_75t_R g27 ( .A(n_17), .B(n_28), .Y(n_27) );
CKINVDCx5p33_ASAP7_75t_R g45 ( .A(n_17), .Y(n_45) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_18), .Y(n_37) );
NAND2xp33_ASAP7_75t_R g18 ( .A(n_19), .B(n_21), .Y(n_18) );
NAND2xp33_ASAP7_75t_R g34 ( .A(n_22), .B(n_35), .Y(n_34) );
NAND2xp33_ASAP7_75t_R g36 ( .A(n_23), .B(n_37), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_27), .Y(n_26) );
CKINVDCx16_ASAP7_75t_R g28 ( .A(n_29), .Y(n_28) );
OAI32xp33_ASAP7_75t_L g30 ( .A1(n_31), .A2(n_39), .A3(n_40), .B1(n_43), .B2(n_46), .Y(n_30) );
NAND2xp33_ASAP7_75t_R g31 ( .A(n_32), .B(n_38), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_33), .B(n_34), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
NOR2xp33_ASAP7_75t_R g44 ( .A(n_40), .B(n_45), .Y(n_44) );
CKINVDCx5p33_ASAP7_75t_R g40 ( .A(n_41), .Y(n_40) );
INVxp33_ASAP7_75t_L g43 ( .A(n_44), .Y(n_43) );
endmodule