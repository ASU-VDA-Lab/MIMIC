module fake_netlist_1_1259_n_46 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_30;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g15 ( .A(n_0), .B(n_8), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_7), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_6), .Y(n_19) );
INVx3_ASAP7_75t_L g20 ( .A(n_6), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_4), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_12), .A2(n_13), .B1(n_10), .B2(n_4), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_16), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_17), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_17), .B(n_0), .Y(n_25) );
INVx2_ASAP7_75t_L g26 ( .A(n_16), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_23), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_25), .Y(n_31) );
A2O1A1Ixp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_29), .B(n_27), .C(n_26), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_31), .B(n_27), .Y(n_33) );
AOI22xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_31), .B1(n_30), .B2(n_17), .Y(n_34) );
OAI22xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_31), .B1(n_22), .B2(n_15), .Y(n_35) );
OAI21xp33_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_22), .B(n_19), .Y(n_36) );
OAI322xp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_19), .A3(n_21), .B1(n_18), .B2(n_20), .C1(n_24), .C2(n_26), .Y(n_37) );
OAI22xp5_ASAP7_75t_L g38 ( .A1(n_34), .A2(n_20), .B1(n_21), .B2(n_18), .Y(n_38) );
XNOR2x1_ASAP7_75t_L g39 ( .A(n_36), .B(n_20), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_38), .Y(n_40) );
AOI222xp33_ASAP7_75t_L g41 ( .A1(n_39), .A2(n_16), .B1(n_2), .B2(n_3), .C1(n_5), .C2(n_7), .Y(n_41) );
BUFx2_ASAP7_75t_L g42 ( .A(n_37), .Y(n_42) );
AND2x2_ASAP7_75t_L g43 ( .A(n_41), .B(n_1), .Y(n_43) );
AOI22xp33_ASAP7_75t_L g44 ( .A1(n_42), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_44) );
A2O1A1Ixp33_ASAP7_75t_L g45 ( .A1(n_43), .A2(n_42), .B(n_40), .C(n_8), .Y(n_45) );
OA22x2_ASAP7_75t_L g46 ( .A1(n_45), .A2(n_44), .B1(n_11), .B2(n_14), .Y(n_46) );
endmodule