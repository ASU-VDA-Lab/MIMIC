module fake_jpeg_1889_n_245 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_245);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_245;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_41),
.B(n_62),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_23),
.B(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_65),
.Y(n_113)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_23),
.B(n_14),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_69),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_16),
.B(n_0),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_20),
.A2(n_13),
.B(n_12),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_19),
.C(n_17),
.Y(n_83)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_73),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_34),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_76),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_1),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_38),
.B1(n_37),
.B2(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_102),
.B1(n_61),
.B2(n_74),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_82),
.A2(n_94),
.B1(n_116),
.B2(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_49),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_100),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g90 ( 
.A1(n_46),
.A2(n_38),
.B1(n_37),
.B2(n_39),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_113),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_52),
.B(n_28),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_55),
.A2(n_26),
.B1(n_18),
.B2(n_4),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_102),
.B1(n_111),
.B2(n_85),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_51),
.B(n_4),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_9),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_57),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_76),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_138),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_68),
.B1(n_73),
.B2(n_60),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_121),
.A2(n_139),
.B1(n_146),
.B2(n_137),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_125),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_132),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_105),
.B1(n_81),
.B2(n_78),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_110),
.Y(n_136)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_136),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_110),
.C(n_113),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_141),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_115),
.B1(n_88),
.B2(n_80),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_114),
.B(n_139),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_89),
.C(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_143),
.Y(n_173)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_92),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_144),
.B(n_145),
.Y(n_164)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_84),
.B(n_96),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_96),
.B(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_134),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_78),
.A3(n_114),
.B1(n_105),
.B2(n_81),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_122),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_159),
.B(n_160),
.C(n_169),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_114),
.B1(n_139),
.B2(n_119),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_161),
.B(n_117),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_169),
.B1(n_161),
.B2(n_158),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_121),
.B1(n_126),
.B2(n_122),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_123),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_174),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_179),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_176),
.A2(n_165),
.B(n_166),
.Y(n_202)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_144),
.C(n_132),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_182),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_131),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_188),
.Y(n_201)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_118),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_125),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_190),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_145),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_186),
.B(n_187),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_143),
.C(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_192),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_160),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_159),
.B1(n_170),
.B2(n_167),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_164),
.A3(n_155),
.B1(n_157),
.B2(n_165),
.C1(n_166),
.C2(n_153),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g207 ( 
.A1(n_195),
.A2(n_176),
.A3(n_175),
.B1(n_168),
.B2(n_157),
.C1(n_189),
.C2(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_205),
.Y(n_212)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_202),
.A2(n_189),
.B(n_178),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_211),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_186),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_187),
.B1(n_189),
.B2(n_192),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_213),
.A2(n_204),
.B1(n_201),
.B2(n_196),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_197),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_215),
.B(n_216),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_168),
.C(n_153),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_205),
.C(n_202),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_219),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_198),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_209),
.B(n_224),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_225),
.C(n_218),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_193),
.C(n_204),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_225),
.A2(n_212),
.B(n_215),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_227),
.A2(n_230),
.B(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_221),
.A2(n_216),
.B1(n_193),
.B2(n_214),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_227),
.A2(n_220),
.B1(n_199),
.B2(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_235),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_206),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_223),
.B(n_210),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_234),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_219),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_237),
.B(n_233),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_240),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_241),
.B(n_203),
.C(n_227),
.Y(n_243)
);

FAx1_ASAP7_75t_SL g244 ( 
.A(n_243),
.B(n_203),
.CI(n_242),
.CON(n_244),
.SN(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_244),
.B(n_243),
.Y(n_245)
);


endmodule