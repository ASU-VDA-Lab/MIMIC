module fake_jpeg_21803_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_18),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_45),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_0),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g62 ( 
.A(n_43),
.B(n_26),
.Y(n_62)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_21),
.B(n_0),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_51),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_21),
.B1(n_28),
.B2(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_57),
.B1(n_60),
.B2(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_58),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_45),
.B1(n_40),
.B2(n_49),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_62),
.A2(n_70),
.B(n_43),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_66),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_43),
.Y(n_99)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_72),
.Y(n_86)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_82),
.Y(n_135)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_80),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_43),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_101),
.Y(n_109)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_44),
.B1(n_50),
.B2(n_66),
.Y(n_123)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_45),
.B1(n_43),
.B2(n_40),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_89),
.B(n_63),
.C(n_60),
.Y(n_108)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_65),
.A2(n_30),
.B1(n_23),
.B2(n_31),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_102),
.B1(n_105),
.B2(n_34),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_98),
.B(n_100),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_48),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_26),
.B1(n_24),
.B2(n_35),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_104),
.Y(n_136)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_65),
.A2(n_27),
.B1(n_33),
.B2(n_34),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_75),
.B1(n_74),
.B2(n_80),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_108),
.A2(n_24),
.B(n_76),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_61),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_111),
.B(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_122),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_54),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_76),
.B(n_100),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_57),
.B(n_53),
.C(n_56),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_119),
.A2(n_121),
.B1(n_124),
.B2(n_53),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_48),
.B1(n_50),
.B2(n_44),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_51),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_125),
.B1(n_108),
.B2(n_122),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_44),
.B1(n_71),
.B2(n_72),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_126),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_51),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_103),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_37),
.B1(n_25),
.B2(n_20),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_137),
.B(n_140),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_159),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_154),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_92),
.B1(n_93),
.B2(n_104),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_151),
.B1(n_155),
.B2(n_166),
.Y(n_168)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_150),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_86),
.C(n_85),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_109),
.C(n_115),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_158),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_147),
.A2(n_157),
.B(n_160),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_112),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_149),
.A2(n_163),
.B1(n_165),
.B2(n_130),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_96),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_87),
.B1(n_83),
.B2(n_82),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_139),
.B(n_110),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_106),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_90),
.Y(n_156)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_103),
.B(n_90),
.C(n_51),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_47),
.Y(n_158)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_161),
.B(n_162),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_112),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_114),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_112),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_172),
.B(n_186),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_164),
.A2(n_132),
.B1(n_113),
.B2(n_116),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_179),
.B(n_193),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_151),
.B(n_20),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_183),
.C(n_185),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_155),
.A2(n_116),
.B1(n_113),
.B2(n_128),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_181),
.A2(n_198),
.B1(n_173),
.B2(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_90),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_184),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_103),
.C(n_47),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_133),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_47),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_192),
.C(n_199),
.Y(n_217)
);

AOI22x1_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_118),
.B1(n_117),
.B2(n_131),
.Y(n_188)
);

AOI22x1_ASAP7_75t_L g230 ( 
.A1(n_188),
.A2(n_36),
.B1(n_32),
.B2(n_29),
.Y(n_230)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_189),
.B(n_194),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_117),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_196),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_114),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_133),
.Y(n_192)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_146),
.B(n_1),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_144),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_149),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_166),
.A2(n_118),
.B1(n_131),
.B2(n_120),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_143),
.B(n_107),
.C(n_17),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_201),
.A2(n_205),
.B1(n_218),
.B2(n_230),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_157),
.Y(n_203)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_204),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_142),
.B(n_148),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_181),
.CI(n_178),
.CON(n_233),
.SN(n_233)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_141),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_165),
.B(n_163),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_149),
.C(n_36),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_187),
.C(n_177),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_221),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_199),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_20),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_168),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_36),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_192),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_228),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_178),
.B(n_2),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_188),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_180),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_241),
.Y(n_266)
);

AO22x1_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_230),
.B1(n_205),
.B2(n_208),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_244),
.C(n_247),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_226),
.B(n_175),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_237),
.B(n_228),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_216),
.A2(n_168),
.B1(n_185),
.B2(n_174),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_196),
.C(n_193),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_20),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_249),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_32),
.C(n_37),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_32),
.C(n_37),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_250),
.C(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_201),
.B(n_25),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_25),
.C(n_3),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_202),
.C(n_203),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_8),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_255),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_8),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_256),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_218),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_264),
.C(n_249),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_R g264 ( 
.A(n_256),
.B(n_230),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_252),
.A2(n_204),
.B1(n_206),
.B2(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_202),
.C(n_206),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_270),
.C(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_271),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_215),
.C(n_212),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_246),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_257),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_219),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_232),
.B(n_231),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_266),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_224),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_277),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_228),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_279),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_274),
.C(n_245),
.Y(n_305)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_296),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_289),
.C(n_294),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_8),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_266),
.C(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_292),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_2),
.B(n_3),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_241),
.C(n_248),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_SL g295 ( 
.A(n_264),
.B(n_233),
.C(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_272),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_276),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_285),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_298),
.A2(n_306),
.B(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_263),
.C(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_263),
.C(n_268),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_274),
.C(n_259),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_284),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_308)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_308),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_9),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_295),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_4),
.C(n_5),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_290),
.C(n_310),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_296),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_318),
.C(n_320),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_283),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_280),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_291),
.C(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_322),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_302),
.B(n_286),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_305),
.B(n_292),
.CI(n_282),
.CON(n_324),
.SN(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_325),
.B(n_327),
.Y(n_336)
);

NOR3x1_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_281),
.C(n_300),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_326),
.A2(n_328),
.B(n_320),
.C(n_313),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_303),
.Y(n_327)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_317),
.B(n_281),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_10),
.B1(n_13),
.B2(n_7),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_317),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_11),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_331),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_334),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_337),
.B(n_338),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_332),
.B(n_315),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_339),
.A2(n_340),
.B1(n_333),
.B2(n_335),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_328),
.A2(n_315),
.B(n_12),
.Y(n_340)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_342),
.A2(n_336),
.B(n_12),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_344),
.A2(n_345),
.B1(n_9),
.B2(n_10),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_343),
.A2(n_341),
.B(n_9),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_10),
.C(n_13),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_5),
.A3(n_6),
.B1(n_15),
.B2(n_337),
.C1(n_341),
.C2(n_326),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_15),
.Y(n_349)
);


endmodule