module fake_jpeg_29799_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVxp67_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_15),
.Y(n_57)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_20),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_12),
.B(n_5),
.Y(n_41)
);

AND2x6_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_15),
.Y(n_65)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_29),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_59),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_65),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g83 ( 
.A(n_60),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_32),
.A2(n_37),
.B1(n_43),
.B2(n_40),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_56),
.B1(n_38),
.B2(n_63),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_14),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_81),
.B1(n_53),
.B2(n_45),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_31),
.B(n_38),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_31),
.C(n_12),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_75),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_25),
.C(n_17),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_26),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_22),
.B1(n_26),
.B2(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_49),
.B(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_46),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_95),
.B(n_83),
.Y(n_106)
);

HAxp5_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_51),
.CON(n_95),
.SN(n_95)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_70),
.B1(n_81),
.B2(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_73),
.C(n_75),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.C(n_104),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_67),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_77),
.C(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_112),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_108),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_70),
.C(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_96),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

AOI221xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_95),
.B1(n_94),
.B2(n_88),
.C(n_81),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_105),
.Y(n_116)
);

AO221x1_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_90),
.B1(n_99),
.B2(n_109),
.C(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_87),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_88),
.B(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

AOI321xp33_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_101),
.A3(n_108),
.B1(n_111),
.B2(n_83),
.C(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_126),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_121),
.C(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_125),
.C(n_48),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_121),
.B(n_115),
.C(n_114),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_129),
.B1(n_131),
.B2(n_123),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_134),
.B(n_8),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_48),
.C(n_56),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_8),
.C(n_10),
.Y(n_134)
);

AOI31xp67_ASAP7_75t_SL g137 ( 
.A1(n_135),
.A2(n_136),
.A3(n_11),
.B(n_51),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_137),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_72),
.B(n_78),
.C(n_22),
.Y(n_139)
);

AOI221xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_72),
.B1(n_78),
.B2(n_26),
.C(n_22),
.Y(n_140)
);


endmodule