module fake_jpeg_1294_n_418 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_418);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_418;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_9),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_59),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_36),
.B(n_15),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_42),
.B(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_54),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_24),
.B(n_1),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_60),
.A2(n_23),
.B(n_17),
.C(n_19),
.Y(n_101)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_24),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_16),
.B1(n_24),
.B2(n_38),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_81),
.A2(n_91),
.B1(n_108),
.B2(n_114),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_85),
.B(n_101),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_16),
.B1(n_58),
.B2(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_39),
.B(n_48),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_59),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_16),
.B1(n_35),
.B2(n_34),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_41),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_38),
.B(n_35),
.C(n_20),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_101),
.B(n_111),
.C(n_105),
.Y(n_122)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_67),
.A2(n_38),
.B1(n_35),
.B2(n_31),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_50),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_117),
.B(n_95),
.C(n_90),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_87),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_146),
.C(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_60),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_139),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g173 ( 
.A(n_122),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_125),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_130),
.B(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_77),
.A2(n_40),
.B1(n_46),
.B2(n_43),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_76),
.B1(n_102),
.B2(n_110),
.Y(n_159)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_82),
.B(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_135),
.B(n_136),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_66),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_70),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_137),
.B(n_138),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_65),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_73),
.B(n_47),
.C(n_63),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g181 ( 
.A1(n_140),
.A2(n_30),
.B1(n_18),
.B2(n_3),
.Y(n_181)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_86),
.A2(n_56),
.B1(n_55),
.B2(n_28),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_150),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_63),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_116),
.B(n_14),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_51),
.B1(n_43),
.B2(n_74),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_153),
.B1(n_157),
.B2(n_92),
.Y(n_180)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_88),
.B(n_80),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_96),
.A2(n_51),
.B1(n_71),
.B2(n_72),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_93),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_63),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_103),
.A2(n_74),
.B1(n_72),
.B2(n_57),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_159),
.A2(n_172),
.B1(n_196),
.B2(n_157),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_104),
.B1(n_90),
.B2(n_75),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_162),
.B(n_164),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_110),
.B1(n_102),
.B2(n_100),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_165),
.A2(n_170),
.B1(n_171),
.B2(n_175),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_124),
.A2(n_100),
.B1(n_76),
.B2(n_95),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_92),
.B1(n_47),
.B2(n_64),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_154),
.A2(n_143),
.B1(n_121),
.B2(n_122),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_92),
.B1(n_47),
.B2(n_20),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_186),
.Y(n_234)
);

AOI32xp33_ASAP7_75t_L g187 ( 
.A1(n_118),
.A2(n_123),
.A3(n_140),
.B1(n_120),
.B2(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_140),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_139),
.A2(n_30),
.B1(n_18),
.B2(n_4),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_188),
.A2(n_152),
.B1(n_147),
.B2(n_149),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_189),
.B(n_190),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_117),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_18),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_191),
.B(n_192),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_117),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_15),
.B1(n_30),
.B2(n_4),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_117),
.B1(n_140),
.B2(n_156),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_204),
.B(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_131),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_203),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_221),
.B1(n_184),
.B2(n_174),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_205),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_194),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_211),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_151),
.B(n_119),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_134),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_213),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_158),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_158),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_215),
.B(n_222),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_177),
.B(n_192),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_217),
.A2(n_228),
.B(n_197),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_218),
.B(n_224),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_148),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_173),
.A2(n_125),
.B1(n_127),
.B2(n_133),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_155),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_141),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_142),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_229),
.Y(n_247)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_232),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_159),
.B1(n_162),
.B2(n_165),
.Y(n_245)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_190),
.A2(n_153),
.B(n_30),
.C(n_5),
.D(n_6),
.Y(n_228)
);

AO22x1_ASAP7_75t_SL g229 ( 
.A1(n_177),
.A2(n_30),
.B1(n_2),
.B2(n_6),
.Y(n_229)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_178),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_211),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_169),
.B1(n_184),
.B2(n_174),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_243),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_191),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_246),
.C(n_255),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_250),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_201),
.B(n_175),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_163),
.B1(n_183),
.B2(n_181),
.Y(n_249)
);

OAI22x1_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_265),
.B1(n_230),
.B2(n_229),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_171),
.B1(n_188),
.B2(n_170),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_224),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_252),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_231),
.A2(n_197),
.B1(n_183),
.B2(n_163),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_254),
.A2(n_259),
.B1(n_269),
.B2(n_208),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_185),
.C(n_178),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_1),
.C(n_2),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_267),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_1),
.B1(n_2),
.B2(n_6),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_215),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_209),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_227),
.A2(n_2),
.B1(n_7),
.B2(n_8),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

AOI22x1_ASAP7_75t_SL g265 ( 
.A1(n_203),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_266),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_219),
.B(n_8),
.C(n_10),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_217),
.Y(n_271)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_272),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_266),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_277),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_276),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_268),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_278),
.B(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_218),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_222),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_262),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_260),
.B(n_223),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_287),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g287 ( 
.A1(n_236),
.A2(n_234),
.A3(n_230),
.B1(n_210),
.B2(n_229),
.C1(n_199),
.C2(n_205),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_257),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_291),
.B1(n_293),
.B2(n_292),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_265),
.Y(n_290)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_290),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_207),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_239),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_248),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_232),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_241),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_294),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_241),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_295),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_236),
.A2(n_198),
.B1(n_234),
.B2(n_230),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_299),
.B1(n_247),
.B2(n_260),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_304),
.A2(n_311),
.B1(n_316),
.B2(n_285),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_291),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_240),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_309),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_242),
.C(n_255),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_320),
.C(n_321),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_237),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_247),
.B1(n_250),
.B2(n_242),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_237),
.B(n_243),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_312),
.A2(n_314),
.B(n_323),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_280),
.B(n_246),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_313),
.B(n_276),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_288),
.A2(n_249),
.B(n_228),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_298),
.A2(n_221),
.B1(n_254),
.B2(n_233),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_258),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_271),
.B(n_256),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_278),
.B(n_256),
.C(n_251),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_324),
.B(n_279),
.C(n_281),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_301),
.B(n_284),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_327),
.B(n_334),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_273),
.B1(n_288),
.B2(n_295),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_275),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_333),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_274),
.Y(n_332)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_277),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_297),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_345),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_337),
.B(n_340),
.Y(n_352)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_306),
.Y(n_338)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_339),
.A2(n_343),
.B1(n_346),
.B2(n_347),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_283),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_341),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_294),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_342),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_313),
.C(n_320),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_336),
.C(n_330),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_286),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_316),
.B1(n_322),
.B2(n_317),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_326),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_303),
.A2(n_290),
.B1(n_300),
.B2(n_293),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_299),
.Y(n_364)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_340),
.Y(n_351)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_351),
.Y(n_367)
);

AOI322xp5_ASAP7_75t_L g354 ( 
.A1(n_329),
.A2(n_303),
.A3(n_315),
.B1(n_314),
.B2(n_323),
.C1(n_332),
.C2(n_326),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_354),
.B(n_328),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_365),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_323),
.C(n_312),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_348),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_329),
.A2(n_321),
.B(n_325),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_363),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_364),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_286),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_370),
.Y(n_387)
);

OA22x2_ASAP7_75t_L g368 ( 
.A1(n_362),
.A2(n_359),
.B1(n_349),
.B2(n_355),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_377),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_335),
.C(n_344),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_345),
.C(n_331),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_372),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_333),
.C(n_310),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_379),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_226),
.Y(n_375)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_375),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_325),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_358),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_270),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_384),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_361),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_390),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_351),
.C(n_360),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_368),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_391),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_373),
.A2(n_362),
.B1(n_299),
.B2(n_364),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_386),
.B(n_382),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_365),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_369),
.A2(n_363),
.B1(n_251),
.B2(n_248),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_381),
.B(n_369),
.Y(n_393)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_393),
.Y(n_404)
);

NAND3xp33_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_373),
.C(n_356),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_395),
.C(n_399),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_378),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_272),
.B1(n_270),
.B2(n_202),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_397),
.A2(n_235),
.B1(n_206),
.B2(n_12),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_388),
.B(n_356),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_400),
.A2(n_383),
.B(n_390),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_267),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_401),
.A2(n_396),
.B(n_398),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_402),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_403),
.B(n_407),
.Y(n_412)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_394),
.A2(n_269),
.B(n_259),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_405),
.A2(n_12),
.B(n_13),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_408),
.B(n_10),
.C(n_11),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_406),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_410),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_413),
.B(n_411),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_415),
.A2(n_412),
.B(n_404),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_12),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_417),
.B(n_13),
.Y(n_418)
);


endmodule