module fake_jpeg_12803_n_39 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_39);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_8),
.B(n_10),
.Y(n_17)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_11),
.B(n_9),
.C(n_7),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_6),
.C(n_2),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_15),
.B1(n_17),
.B2(n_14),
.Y(n_23)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_16),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_18),
.B(n_20),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_24),
.C(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_15),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_21),
.B(n_22),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_34),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_1),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_26),
.C2(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_3),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_37),
.B(n_5),
.Y(n_39)
);


endmodule