module fake_jpeg_22323_n_191 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_191);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_191;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_38),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_36),
.Y(n_48)
);

OR2x4_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_35),
.A2(n_39),
.B(n_24),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.C(n_3),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_4),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_14),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_16),
.B1(n_20),
.B2(n_29),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_66),
.B1(n_71),
.B2(n_73),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_22),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_68),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_20),
.B1(n_29),
.B2(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_33),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_20),
.B1(n_29),
.B2(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_15),
.B1(n_24),
.B2(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_64),
.Y(n_83)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_33),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_63),
.A2(n_52),
.B(n_47),
.C(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_19),
.B1(n_17),
.B2(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_67),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_23),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_18),
.B1(n_31),
.B2(n_7),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_75),
.B(n_76),
.Y(n_111)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_80),
.Y(n_117)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_95),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_9),
.B(n_10),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_91),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_50),
.A2(n_33),
.B1(n_42),
.B2(n_43),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_78),
.B1(n_88),
.B2(n_80),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_31),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_98),
.C(n_9),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_4),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_73),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_99),
.B(n_67),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_71),
.A2(n_43),
.B1(n_31),
.B2(n_8),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_49),
.B1(n_60),
.B2(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_6),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_12),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_6),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_70),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_70),
.B1(n_51),
.B2(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_104),
.B1(n_118),
.B2(n_119),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_113),
.B(n_119),
.C(n_112),
.Y(n_136)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_9),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_112),
.C(n_116),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_109),
.B(n_93),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_95),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_10),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_115),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_47),
.Y(n_112)
);

XNOR2x2_ASAP7_75t_SL g113 ( 
.A(n_75),
.B(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_12),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_114),
.B(n_98),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_76),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_52),
.C(n_74),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_89),
.B1(n_92),
.B2(n_99),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_52),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_83),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_13),
.B1(n_74),
.B2(n_100),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_133),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_137),
.B(n_114),
.Y(n_144)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_147)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_149),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_137),
.B(n_127),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_102),
.B1(n_116),
.B2(n_101),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_145),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_112),
.B(n_103),
.C(n_109),
.D(n_122),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_149),
.C(n_131),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_112),
.C(n_106),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_122),
.B1(n_106),
.B2(n_105),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_122),
.B1(n_121),
.B2(n_107),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_155),
.B1(n_153),
.B2(n_151),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_139),
.B1(n_130),
.B2(n_141),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_134),
.A3(n_128),
.B1(n_124),
.B2(n_138),
.C1(n_77),
.C2(n_96),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_158),
.C(n_161),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_160),
.B(n_150),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_133),
.B(n_135),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_125),
.C(n_97),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_124),
.C(n_123),
.Y(n_164)
);

OAI321xp33_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_122),
.A3(n_120),
.B1(n_135),
.B2(n_110),
.C(n_77),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_148),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_172),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_147),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_166),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_154),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_174),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_154),
.B1(n_146),
.B2(n_142),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_162),
.C(n_142),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_96),
.C(n_84),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_175),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_185),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_169),
.C(n_170),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_132),
.C(n_13),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_171),
.B(n_79),
.Y(n_185)
);

AOI321xp33_ASAP7_75t_SL g186 ( 
.A1(n_182),
.A2(n_179),
.A3(n_176),
.B1(n_84),
.B2(n_132),
.C(n_115),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_74),
.B(n_187),
.Y(n_190)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_189),
.Y(n_191)
);


endmodule