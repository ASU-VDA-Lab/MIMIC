module fake_netlist_1_12335_n_722 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_722);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_722;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_8), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_35), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_88), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_70), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_34), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_103), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_101), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_17), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_20), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_4), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_62), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_24), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_4), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_86), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_11), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_57), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_21), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_26), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_98), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_30), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_8), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_33), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_58), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_1), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_60), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_76), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_79), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_42), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_65), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_67), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_46), .Y(n_143) );
NOR2xp67_ASAP7_75t_L g144 ( .A(n_77), .B(n_16), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_2), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_16), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_3), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_52), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_25), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_116), .B(n_19), .Y(n_153) );
OA21x2_ASAP7_75t_L g154 ( .A1(n_118), .A2(n_53), .B(n_105), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_107), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_114), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_108), .B(n_0), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_123), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_111), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_113), .B(n_3), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_111), .B(n_5), .Y(n_163) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_127), .A2(n_55), .B(n_104), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_114), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_134), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_107), .Y(n_169) );
AOI22xp5_ASAP7_75t_SL g170 ( .A1(n_136), .A2(n_6), .B1(n_7), .B2(n_9), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
CKINVDCx6p67_ASAP7_75t_R g174 ( .A(n_169), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_169), .B(n_110), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_165), .B(n_110), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_155), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_165), .B(n_137), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_154), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_153), .Y(n_181) );
INVx3_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_167), .B(n_138), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_167), .B(n_112), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_159), .B(n_112), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_156), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_168), .B(n_139), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_153), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_175), .B(n_168), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_196), .B(n_139), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_179), .B(n_158), .Y(n_199) );
INVx8_ASAP7_75t_L g200 ( .A(n_196), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_174), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_182), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_194), .A2(n_166), .B1(n_163), .B2(n_136), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_179), .B(n_160), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_196), .B(n_140), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_182), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_182), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_192), .B(n_160), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_194), .B(n_163), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_192), .B(n_160), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_194), .B(n_140), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_185), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_196), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_192), .B(n_151), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_174), .A2(n_166), .B1(n_170), .B2(n_162), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_178), .A2(n_153), .B1(n_162), .B2(n_145), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_176), .B(n_151), .Y(n_217) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_174), .A2(n_120), .B1(n_117), .B2(n_124), .Y(n_218) );
NAND2xp33_ASAP7_75t_L g219 ( .A(n_196), .B(n_153), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_178), .B(n_161), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_191), .B(n_153), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_190), .B(n_153), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_190), .B(n_153), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_196), .B(n_115), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_181), .B(n_161), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_189), .B(n_119), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_181), .B(n_121), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_189), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_201), .B(n_196), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_208), .A2(n_193), .B(n_188), .C(n_187), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_210), .A2(n_193), .B(n_188), .C(n_187), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_215), .A2(n_188), .B(n_187), .C(n_148), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_188), .B(n_187), .C(n_186), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_209), .B(n_181), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_212), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_218), .B(n_195), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_211), .B(n_195), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_223), .A2(n_195), .B(n_186), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_214), .B(n_204), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_201), .B(n_170), .Y(n_242) );
AOI22x1_ASAP7_75t_L g243 ( .A1(n_212), .A2(n_186), .B1(n_184), .B2(n_183), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_213), .B(n_125), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_224), .A2(n_184), .B(n_183), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g246 ( .A(n_203), .B(n_9), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_213), .B(n_128), .Y(n_247) );
AOI221x1_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_180), .B1(n_183), .B2(n_184), .C(n_150), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_199), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_217), .B(n_157), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_202), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_221), .B(n_132), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_227), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_202), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_227), .A2(n_147), .B(n_141), .C(n_142), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_221), .B(n_180), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_230), .Y(n_257) );
AOI21x1_ASAP7_75t_L g258 ( .A1(n_230), .A2(n_154), .B(n_164), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
AO22x1_ASAP7_75t_L g260 ( .A1(n_202), .A2(n_180), .B1(n_143), .B2(n_146), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_216), .B(n_180), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_237), .B(n_213), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_245), .A2(n_219), .B(n_226), .Y(n_263) );
AOI211x1_ASAP7_75t_L g264 ( .A1(n_241), .A2(n_149), .B(n_228), .C(n_198), .Y(n_264) );
BUFx10_ASAP7_75t_L g265 ( .A(n_231), .Y(n_265) );
AO21x1_ASAP7_75t_L g266 ( .A1(n_261), .A2(n_219), .B(n_220), .Y(n_266) );
BUFx2_ASAP7_75t_L g267 ( .A(n_257), .Y(n_267) );
AO31x2_ASAP7_75t_L g268 ( .A1(n_248), .A2(n_220), .A3(n_207), .B(n_206), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_250), .B(n_207), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_257), .A2(n_180), .B1(n_157), .B2(n_229), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_231), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_253), .B(n_180), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_231), .Y(n_273) );
OAI21x1_ASAP7_75t_SL g274 ( .A1(n_237), .A2(n_164), .B(n_180), .Y(n_274) );
OAI21x1_ASAP7_75t_SL g275 ( .A1(n_234), .A2(n_164), .B(n_200), .Y(n_275) );
BUFx3_ASAP7_75t_L g276 ( .A(n_251), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_243), .A2(n_164), .B(n_225), .Y(n_277) );
AO31x2_ASAP7_75t_L g278 ( .A1(n_248), .A2(n_235), .A3(n_233), .B(n_232), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_251), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_243), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_246), .B(n_205), .Y(n_281) );
AOI221x1_ASAP7_75t_L g282 ( .A1(n_261), .A2(n_126), .B1(n_135), .B2(n_173), .C(n_172), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_164), .B(n_144), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_258), .A2(n_240), .B(n_256), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_236), .A2(n_172), .B(n_171), .Y(n_285) );
NOR2x1_ASAP7_75t_L g286 ( .A(n_238), .B(n_171), .Y(n_286) );
AO21x2_ASAP7_75t_L g287 ( .A1(n_275), .A2(n_255), .B(n_259), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_272), .Y(n_288) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_275), .A2(n_239), .B(n_259), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_282), .A2(n_247), .B(n_244), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_280), .A2(n_260), .B(n_254), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_267), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_270), .A2(n_242), .B1(n_249), .B2(n_126), .Y(n_293) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_282), .A2(n_252), .B(n_260), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_280), .A2(n_173), .B(n_177), .Y(n_295) );
NAND2x1p5_ASAP7_75t_L g296 ( .A(n_279), .B(n_251), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_267), .B(n_242), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_284), .A2(n_254), .B(n_177), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_272), .Y(n_299) );
AO21x2_ASAP7_75t_L g300 ( .A1(n_266), .A2(n_177), .B(n_135), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_279), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_284), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_277), .A2(n_254), .B(n_200), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_266), .A2(n_126), .B(n_135), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_277), .A2(n_200), .B(n_63), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
AO21x2_ASAP7_75t_L g307 ( .A1(n_274), .A2(n_135), .B(n_11), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_269), .B(n_200), .Y(n_308) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_292), .Y(n_309) );
NAND2x1_ASAP7_75t_L g310 ( .A(n_302), .B(n_279), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_302), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_288), .B(n_278), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_288), .B(n_279), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_302), .Y(n_315) );
OA21x2_ASAP7_75t_L g316 ( .A1(n_303), .A2(n_283), .B(n_274), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_299), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_292), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_292), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_303), .A2(n_283), .B(n_263), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
OAI21x1_ASAP7_75t_L g323 ( .A1(n_305), .A2(n_286), .B(n_262), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_296), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_302), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_298), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_297), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_299), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_301), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_301), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_301), .B(n_276), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_306), .Y(n_335) );
INVx2_ASAP7_75t_SL g336 ( .A(n_310), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_313), .B(n_304), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_312), .B(n_300), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_313), .B(n_287), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_324), .B(n_298), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_317), .B(n_287), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_327), .B(n_297), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_311), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_317), .B(n_319), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_329), .B(n_287), .Y(n_348) );
OAI221xp5_ASAP7_75t_L g349 ( .A1(n_318), .A2(n_293), .B1(n_281), .B2(n_291), .C(n_308), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_329), .B(n_287), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_324), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_311), .Y(n_352) );
NOR4xp25_ASAP7_75t_SL g353 ( .A(n_318), .B(n_306), .C(n_307), .D(n_304), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_312), .B(n_287), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_331), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_314), .B(n_298), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_335), .B(n_287), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_330), .B(n_304), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_315), .B(n_325), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_314), .B(n_298), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_332), .A2(n_293), .B1(n_308), .B2(n_289), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_322), .A2(n_291), .B1(n_264), .B2(n_294), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_309), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_323), .A2(n_304), .B(n_307), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_331), .B(n_304), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_325), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_320), .B(n_271), .Y(n_369) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_322), .A2(n_303), .B(n_305), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_333), .B(n_300), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_300), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_335), .B(n_300), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_314), .B(n_300), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_320), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_325), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_328), .B(n_314), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_347), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_346), .B(n_334), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_342), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_338), .B(n_307), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_338), .B(n_307), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_351), .B(n_334), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_365), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_307), .Y(n_387) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_343), .B(n_316), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_346), .B(n_334), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_337), .B(n_326), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_365), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_344), .A2(n_289), .B1(n_334), .B2(n_271), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_337), .B(n_326), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_347), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_376), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_376), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_367), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_367), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_377), .B(n_289), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_371), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_371), .B(n_326), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_369), .B(n_306), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_379), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_372), .B(n_326), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_342), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_358), .B(n_264), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_357), .B(n_326), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_375), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_373), .B(n_316), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_374), .B(n_316), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_374), .B(n_316), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_378), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_359), .B(n_321), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_375), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
OR2x2_ASAP7_75t_L g421 ( .A(n_377), .B(n_321), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_359), .B(n_321), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_361), .B(n_321), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_361), .B(n_295), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g426 ( .A(n_336), .B(n_10), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_358), .B(n_278), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_351), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_345), .Y(n_429) );
AND2x2_ASAP7_75t_SL g430 ( .A(n_370), .B(n_294), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_339), .B(n_295), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_339), .B(n_295), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_341), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_341), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_348), .B(n_278), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_345), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_348), .B(n_295), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_350), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_350), .B(n_278), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_354), .B(n_278), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_345), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_351), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_354), .B(n_295), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_352), .Y(n_444) );
INVx3_ASAP7_75t_SL g445 ( .A(n_340), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_352), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_386), .B(n_352), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_445), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_380), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_403), .B(n_363), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_403), .B(n_363), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_415), .B(n_357), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_380), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_382), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_395), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_397), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_407), .B(n_355), .Y(n_458) );
AND2x2_ASAP7_75t_SL g459 ( .A(n_442), .B(n_370), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_407), .B(n_355), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_417), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_420), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_391), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_398), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_413), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_382), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_415), .B(n_357), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_416), .B(n_357), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_399), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_416), .B(n_362), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_381), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_389), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_412), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_393), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_362), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_411), .B(n_362), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_445), .B(n_412), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_411), .B(n_362), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_393), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_400), .B(n_355), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_400), .B(n_340), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_401), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_401), .B(n_340), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_385), .B(n_336), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_402), .B(n_360), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_402), .B(n_360), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_404), .B(n_340), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_433), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_409), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_433), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_434), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_434), .B(n_360), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_438), .B(n_368), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_438), .Y(n_495) );
NOR2xp67_ASAP7_75t_L g496 ( .A(n_428), .B(n_336), .Y(n_496) );
INVxp33_ASAP7_75t_L g497 ( .A(n_385), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_426), .B(n_343), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_368), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_446), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_404), .B(n_379), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_408), .B(n_379), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_409), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_392), .A2(n_349), .B1(n_353), .B2(n_368), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_388), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_408), .B(n_379), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_443), .B(n_364), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_383), .B(n_364), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_446), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_429), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_429), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_383), .B(n_366), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_384), .B(n_366), .Y(n_513) );
INVxp33_ASAP7_75t_L g514 ( .A(n_385), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_444), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_405), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_436), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_384), .B(n_366), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_387), .A2(n_349), .B1(n_366), .B2(n_343), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_387), .B(n_353), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_390), .B(n_370), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_436), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_414), .B(n_370), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_390), .B(n_370), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_394), .B(n_343), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_394), .B(n_323), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_441), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_414), .B(n_12), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_441), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_474), .Y(n_530) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_498), .B(n_388), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_483), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_448), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_489), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_452), .B(n_411), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
INVxp67_ASAP7_75t_L g537 ( .A(n_465), .Y(n_537) );
NOR2x1p5_ASAP7_75t_SL g538 ( .A(n_454), .B(n_421), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_513), .B(n_418), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_452), .B(n_418), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_466), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_475), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_513), .B(n_423), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_497), .A2(n_421), .B1(n_410), .B2(n_440), .Y(n_545) );
NOR2x1_ASAP7_75t_L g546 ( .A(n_498), .B(n_431), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_448), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_499), .B(n_423), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_472), .B(n_425), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_492), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
OAI221xp5_ASAP7_75t_SL g552 ( .A1(n_519), .A2(n_439), .B1(n_427), .B2(n_435), .C(n_425), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_465), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_516), .B(n_424), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_467), .B(n_424), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_475), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_496), .B(n_294), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_461), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_503), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_473), .B(n_431), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_467), .B(n_432), .Y(n_561) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_485), .B(n_432), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_468), .B(n_437), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_462), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_468), .B(n_437), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_471), .B(n_406), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_471), .B(n_427), .Y(n_568) );
AOI32xp33_ASAP7_75t_L g569 ( .A1(n_497), .A2(n_439), .A3(n_435), .B1(n_305), .B2(n_323), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_447), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_455), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_470), .B(n_430), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_486), .B(n_406), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_487), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_456), .Y(n_575) );
INVx2_ASAP7_75t_SL g576 ( .A(n_478), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_507), .B(n_430), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_450), .B(n_406), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_454), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_451), .B(n_406), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_463), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_523), .B(n_406), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_512), .B(n_294), .Y(n_583) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_480), .Y(n_584) );
OAI33xp33_ASAP7_75t_L g585 ( .A1(n_504), .A2(n_13), .A3(n_14), .B1(n_15), .B2(n_17), .B3(n_18), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_457), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_520), .B(n_294), .C(n_290), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_476), .B(n_303), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_464), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_SL g590 ( .A1(n_514), .A2(n_13), .B(n_14), .C(n_15), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_518), .B(n_294), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_488), .B(n_305), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_480), .Y(n_593) );
INVxp67_ASAP7_75t_L g594 ( .A(n_528), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_525), .B(n_295), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_469), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_449), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_490), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_490), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_525), .B(n_296), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_453), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_515), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_500), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_509), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_458), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_581), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_541), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_562), .A2(n_459), .B1(n_524), .B2(n_521), .Y(n_609) );
OAI22xp33_ASAP7_75t_SL g610 ( .A1(n_546), .A2(n_485), .B1(n_505), .B2(n_508), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_540), .B(n_477), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_533), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_554), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_577), .B(n_521), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_547), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_554), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_535), .B(n_477), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_539), .B(n_524), .Y(n_618) );
OAI22xp33_ASAP7_75t_SL g619 ( .A1(n_552), .A2(n_485), .B1(n_505), .B2(n_477), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_576), .A2(n_514), .B1(n_459), .B2(n_479), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_559), .Y(n_621) );
OR2x6_ASAP7_75t_L g622 ( .A(n_538), .B(n_505), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_590), .A2(n_481), .B(n_460), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_555), .B(n_479), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_552), .A2(n_482), .B1(n_484), .B2(n_526), .C(n_494), .Y(n_625) );
INVxp67_ASAP7_75t_L g626 ( .A(n_605), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g627 ( .A1(n_565), .A2(n_479), .B1(n_493), .B2(n_501), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_585), .A2(n_526), .B1(n_502), .B2(n_506), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_585), .A2(n_527), .B1(n_529), .B2(n_522), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_569), .A2(n_529), .B(n_522), .C(n_517), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_594), .A2(n_517), .B(n_511), .Y(n_631) );
OAI21xp33_ASAP7_75t_L g632 ( .A1(n_577), .A2(n_511), .B(n_510), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_584), .Y(n_633) );
INVxp33_ASAP7_75t_L g634 ( .A(n_531), .Y(n_634) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_594), .A2(n_510), .B(n_18), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_558), .Y(n_636) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_537), .A2(n_296), .B(n_290), .Y(n_637) );
AOI322xp5_ASAP7_75t_L g638 ( .A1(n_539), .A2(n_286), .A3(n_273), .B1(n_290), .B2(n_276), .C1(n_131), .C2(n_133), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_572), .B(n_290), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_537), .A2(n_296), .B(n_290), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_545), .A2(n_290), .B(n_273), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
OAI21xp5_ASAP7_75t_L g643 ( .A1(n_553), .A2(n_296), .B(n_285), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_572), .B(n_268), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_544), .A2(n_23), .B(n_28), .Y(n_645) );
INVx1_ASAP7_75t_SL g646 ( .A(n_548), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_564), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_553), .B(n_268), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_571), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_570), .B(n_265), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_595), .A2(n_265), .B1(n_268), .B2(n_32), .Y(n_651) );
OAI21xp5_ASAP7_75t_SL g652 ( .A1(n_588), .A2(n_265), .B(n_31), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_559), .A2(n_268), .B(n_265), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_575), .A2(n_29), .B1(n_36), .B2(n_37), .C(n_38), .Y(n_654) );
OAI21xp5_ASAP7_75t_L g655 ( .A1(n_557), .A2(n_39), .B(n_40), .Y(n_655) );
O2A1O1Ixp33_ASAP7_75t_L g656 ( .A1(n_619), .A2(n_589), .B(n_586), .C(n_596), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_652), .A2(n_557), .B(n_592), .Y(n_657) );
CKINVDCx14_ASAP7_75t_R g658 ( .A(n_621), .Y(n_658) );
OR2x2_ASAP7_75t_L g659 ( .A(n_618), .B(n_544), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_625), .A2(n_582), .B1(n_580), .B2(n_578), .C(n_534), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_609), .A2(n_568), .B1(n_560), .B2(n_549), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_630), .A2(n_582), .B1(n_580), .B2(n_578), .C(n_551), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_610), .A2(n_584), .B(n_556), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g664 ( .A1(n_634), .A2(n_574), .B(n_567), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_612), .A2(n_563), .B(n_561), .C(n_530), .Y(n_665) );
OAI222xp33_ASAP7_75t_L g666 ( .A1(n_622), .A2(n_542), .B1(n_550), .B2(n_532), .C1(n_583), .C2(n_591), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_626), .A2(n_601), .B1(n_597), .B2(n_604), .C(n_603), .Y(n_667) );
NAND3xp33_ASAP7_75t_L g668 ( .A(n_629), .B(n_587), .C(n_543), .Y(n_668) );
OAI21xp33_ASAP7_75t_SL g669 ( .A1(n_622), .A2(n_536), .B(n_566), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_628), .B(n_591), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_620), .A2(n_600), .B(n_583), .C(n_573), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_615), .B(n_623), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_631), .A2(n_599), .B1(n_598), .B2(n_593), .C(n_579), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_636), .B(n_41), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_622), .A2(n_268), .B(n_44), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_646), .A2(n_43), .B1(n_45), .B2(n_47), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_635), .A2(n_606), .B(n_648), .Y(n_677) );
XNOR2x1_ASAP7_75t_L g678 ( .A(n_627), .B(n_48), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_628), .A2(n_49), .B1(n_50), .B2(n_51), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_613), .A2(n_54), .B1(n_56), .B2(n_59), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_614), .A2(n_61), .B1(n_64), .B2(n_68), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_616), .A2(n_69), .B1(n_71), .B2(n_72), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g683 ( .A1(n_632), .A2(n_73), .B1(n_74), .B2(n_75), .C(n_78), .Y(n_683) );
AOI221x1_ASAP7_75t_L g684 ( .A1(n_670), .A2(n_645), .B1(n_649), .B2(n_647), .C(n_642), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_656), .A2(n_641), .B(n_643), .C(n_653), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_658), .B(n_617), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_659), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_672), .A2(n_655), .B(n_644), .C(n_654), .Y(n_688) );
AOI221x1_ASAP7_75t_L g689 ( .A1(n_677), .A2(n_607), .B1(n_608), .B2(n_633), .C(n_639), .Y(n_689) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_669), .A2(n_624), .A3(n_611), .B1(n_651), .B2(n_650), .C1(n_638), .C2(n_640), .Y(n_690) );
NAND4xp25_ASAP7_75t_SL g691 ( .A(n_679), .B(n_651), .C(n_637), .D(n_82), .Y(n_691) );
AOI31xp33_ASAP7_75t_L g692 ( .A1(n_678), .A2(n_80), .A3(n_81), .B(n_83), .Y(n_692) );
NAND4xp75_ASAP7_75t_L g693 ( .A(n_663), .B(n_84), .C(n_85), .D(n_87), .Y(n_693) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_668), .A2(n_90), .B(n_91), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_665), .B(n_92), .Y(n_695) );
OA21x2_ASAP7_75t_L g696 ( .A1(n_664), .A2(n_94), .B(n_95), .Y(n_696) );
OAI211xp5_ASAP7_75t_L g697 ( .A1(n_657), .A2(n_96), .B(n_99), .C(n_100), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_690), .A2(n_660), .B(n_671), .C(n_662), .Y(n_698) );
AND4x1_ASAP7_75t_L g699 ( .A(n_684), .B(n_674), .C(n_675), .D(n_667), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_692), .A2(n_666), .B(n_675), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_687), .B(n_673), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_696), .A2(n_661), .B(n_683), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_686), .B(n_676), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g704 ( .A1(n_691), .A2(n_681), .B(n_680), .C(n_682), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_701), .B(n_690), .Y(n_705) );
NAND4xp75_ASAP7_75t_L g706 ( .A(n_702), .B(n_689), .C(n_695), .D(n_694), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_699), .B(n_697), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g708 ( .A(n_698), .B(n_693), .C(n_685), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_708), .B(n_703), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_705), .Y(n_710) );
NAND3xp33_ASAP7_75t_L g711 ( .A(n_707), .B(n_700), .C(n_704), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_709), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_713), .B(n_710), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_714), .B(n_706), .Y(n_716) );
OA21x2_ASAP7_75t_L g717 ( .A1(n_715), .A2(n_688), .B(n_696), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_716), .A2(n_715), .B(n_106), .Y(n_718) );
OA21x2_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_716), .B(n_717), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_719), .B(n_716), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_720), .B(n_717), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_102), .B1(n_213), .B2(n_717), .C(n_713), .Y(n_722) );
endmodule