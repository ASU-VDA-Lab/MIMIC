module real_jpeg_26040_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_344, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_344;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_1),
.A2(n_69),
.B(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_1),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_1),
.B(n_61),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_122),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_1),
.B(n_43),
.C(n_48),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_1),
.B(n_29),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_1),
.A2(n_98),
.B1(n_215),
.B2(n_222),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_54),
.B1(n_75),
.B2(n_113),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_113),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_113),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_27),
.B1(n_69),
.B2(n_75),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_6),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_8),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_67),
.Y(n_299)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_10),
.A2(n_56),
.B1(n_75),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_10),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_125),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_125),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_125),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_11),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_11),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_57),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_13),
.A2(n_25),
.B1(n_28),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_13),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_115),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_115),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_13),
.A2(n_54),
.B1(n_68),
.B2(n_115),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_38),
.B1(n_56),
.B2(n_75),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_14),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_105)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_15),
.Y(n_143)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_15),
.Y(n_216)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_15),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_83),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_71),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_20),
.B(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_39),
.C(n_51),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_21),
.A2(n_22),
.B1(n_39),
.B2(n_323),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_23),
.A2(n_111),
.B(n_114),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_24),
.A2(n_29),
.B(n_35),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_24),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_28),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_25),
.A2(n_63),
.B(n_121),
.C(n_137),
.Y(n_136)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_25),
.B(n_122),
.CON(n_167),
.SN(n_167)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_28),
.B(n_55),
.C(n_62),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_28),
.A2(n_30),
.A3(n_32),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_29),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_29),
.A2(n_35),
.B1(n_158),
.B2(n_167),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_29),
.B(n_37),
.Y(n_264)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_32),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_31),
.B(n_33),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_32),
.B(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_34),
.A2(n_116),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_35),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_39),
.A2(n_319),
.B1(n_320),
.B2(n_323),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_39),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_41),
.A2(n_50),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_41),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_41),
.A2(n_176),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_41),
.A2(n_175),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_41),
.A2(n_174),
.B1(n_175),
.B2(n_195),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_41),
.A2(n_175),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_41),
.A2(n_109),
.B(n_254),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_46),
.B(n_96),
.Y(n_109)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_46),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_46),
.B(n_49),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_46),
.B(n_122),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_47),
.B(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_51),
.B(n_328),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_59),
.B1(n_61),
.B2(n_66),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_53),
.A2(n_60),
.B(n_77),
.Y(n_316)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_66),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_59),
.A2(n_61),
.B1(n_124),
.B2(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_59),
.A2(n_61),
.B1(n_132),
.B2(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_59),
.A2(n_80),
.B(n_260),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_59),
.A2(n_73),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_60),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_117)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_65),
.B(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_340),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_70),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_81),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_336),
.B(n_341),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_312),
.A3(n_331),
.B1(n_334),
.B2(n_335),
.C(n_344),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_290),
.B(n_311),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_269),
.B(n_289),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_159),
.B(n_244),
.C(n_268),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_144),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_128),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_106),
.B1(n_126),
.B2(n_127),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_91),
.B(n_127),
.C(n_128),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_92),
.B(n_97),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_93),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_94),
.B(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B(n_104),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_98),
.A2(n_104),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_98),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_98),
.A2(n_212),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_98),
.A2(n_170),
.B(n_223),
.Y(n_277)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_103),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_99),
.B(n_105),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_99),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_101),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_117),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_111),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_111),
.A2(n_116),
.B1(n_285),
.B2(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_122),
.B(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_131),
.B(n_133),
.C(n_135),
.Y(n_266)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_138),
.B1(n_139),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_150),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_145),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_148),
.B(n_150),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_156),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_154),
.B1(n_155),
.B2(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_151),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_153),
.B(n_206),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_239),
.B(n_243),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_189),
.B(n_238),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_177),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_164),
.B(n_177),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_172),
.C(n_173),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_165),
.B(n_236),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_172),
.B(n_173),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_185),
.C(n_188),
.Y(n_240)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_187),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_233),
.B(n_237),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_208),
.B(n_232),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_192),
.B(n_198),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_196),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_203),
.C(n_204),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_202),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_218),
.B(n_231),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_217),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_217),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_225),
.B(n_230),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_220),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_240),
.B(n_241),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_246),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_266),
.B2(n_267),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_256),
.C(n_267),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_255),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_252),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_261),
.C(n_265),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_266),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_270),
.B(n_271),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_288),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_278),
.B1(n_286),
.B2(n_287),
.Y(n_272)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_287),
.C(n_288),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_276),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_276),
.A2(n_277),
.B1(n_303),
.B2(n_305),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_305),
.B(n_306),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_292),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_309),
.B2(n_310),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_301),
.B1(n_307),
.B2(n_308),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_295),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_308),
.C(n_310),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_298),
.B(n_300),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_298),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_314),
.C(n_324),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_314),
.CI(n_324),
.CON(n_333),
.SN(n_333)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_303),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_325),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_313),
.B(n_325),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_316),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_320),
.C(n_323),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_329),
.C(n_330),
.Y(n_337)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_327),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_333),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_338),
.Y(n_341)
);


endmodule