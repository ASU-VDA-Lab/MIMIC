module fake_jpeg_28353_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_46),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_54),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_39),
.B(n_37),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_9),
.B(n_10),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_43),
.B1(n_44),
.B2(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_1),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_42),
.B1(n_47),
.B2(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_5),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_16),
.B1(n_17),
.B2(n_22),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_7),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_61),
.B(n_66),
.Y(n_75)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_79),
.B(n_15),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_12),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_13),
.B(n_14),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_26),
.B(n_27),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_79),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_24),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_70),
.B1(n_75),
.B2(n_78),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_88),
.A2(n_90),
.B(n_91),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_84),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_83),
.B(n_80),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_94),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_28),
.B(n_29),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_30),
.C(n_32),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_33),
.Y(n_102)
);


endmodule