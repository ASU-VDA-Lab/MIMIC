module fake_netlist_1_4384_n_20 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_20);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
INVx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
NAND2xp5_ASAP7_75t_SL g10 ( .A(n_4), .B(n_5), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_1), .B(n_5), .Y(n_12) );
NOR2xp67_ASAP7_75t_L g13 ( .A(n_11), .B(n_0), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_9), .B(n_0), .Y(n_14) );
BUFx2_ASAP7_75t_L g15 ( .A(n_14), .Y(n_15) );
NOR2xp33_ASAP7_75t_L g16 ( .A(n_15), .B(n_13), .Y(n_16) );
OAI21xp5_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_15), .B(n_12), .Y(n_17) );
NAND4xp75_ASAP7_75t_L g18 ( .A(n_17), .B(n_10), .C(n_3), .D(n_4), .Y(n_18) );
OAI22xp5_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_2), .B1(n_3), .B2(n_6), .Y(n_19) );
AOI22xp33_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_2), .B1(n_6), .B2(n_7), .Y(n_20) );
endmodule