module fake_aes_7115_n_1269 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1269);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1269;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_283;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_281;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_280;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_282;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVx2_ASAP7_75t_L g277 ( .A(n_224), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_252), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_227), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_239), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_207), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_86), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_143), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_150), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_6), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_221), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_52), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_263), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_17), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_171), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_194), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_62), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_179), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_265), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_113), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_20), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_152), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_39), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_111), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_202), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_6), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_225), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_147), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_4), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_236), .Y(n_306) );
INVxp67_ASAP7_75t_SL g307 ( .A(n_134), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_185), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_20), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_174), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_248), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_71), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_89), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_222), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_178), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_216), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_156), .Y(n_317) );
BUFx5_ASAP7_75t_L g318 ( .A(n_23), .Y(n_318) );
BUFx10_ASAP7_75t_L g319 ( .A(n_23), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_51), .Y(n_320) );
INVxp33_ASAP7_75t_L g321 ( .A(n_241), .Y(n_321) );
CKINVDCx14_ASAP7_75t_R g322 ( .A(n_71), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_127), .Y(n_323) );
CKINVDCx14_ASAP7_75t_R g324 ( .A(n_189), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_217), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_155), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_160), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_212), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_80), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_269), .Y(n_330) );
NOR2xp67_ASAP7_75t_L g331 ( .A(n_235), .B(n_146), .Y(n_331) );
CKINVDCx14_ASAP7_75t_R g332 ( .A(n_11), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_131), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_21), .Y(n_334) );
CKINVDCx16_ASAP7_75t_R g335 ( .A(n_97), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_165), .Y(n_336) );
CKINVDCx16_ASAP7_75t_R g337 ( .A(n_45), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_242), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_128), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_149), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_211), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_264), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_123), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_130), .Y(n_344) );
BUFx6f_ASAP7_75t_L g345 ( .A(n_35), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_176), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_177), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_191), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_254), .B(n_270), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_62), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_108), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_168), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_120), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_186), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_46), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_157), .Y(n_356) );
INVx2_ASAP7_75t_SL g357 ( .A(n_209), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_54), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_55), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_243), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_249), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_173), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_91), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_63), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_210), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_139), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_19), .B(n_151), .Y(n_367) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_76), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_198), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_162), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_142), .Y(n_371) );
INVxp67_ASAP7_75t_SL g372 ( .A(n_145), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g373 ( .A(n_136), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_244), .Y(n_374) );
CKINVDCx14_ASAP7_75t_R g375 ( .A(n_274), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_110), .Y(n_376) );
NOR2xp67_ASAP7_75t_L g377 ( .A(n_27), .B(n_163), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_90), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_208), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_1), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_167), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_154), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_39), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_43), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_17), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_40), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_268), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_273), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_44), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_73), .Y(n_390) );
CKINVDCx16_ASAP7_75t_R g391 ( .A(n_144), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_153), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_201), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_97), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_148), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_67), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g397 ( .A(n_245), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_138), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_57), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_7), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_205), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_199), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_255), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_26), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_82), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_64), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_89), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_81), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_37), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_5), .Y(n_410) );
CKINVDCx5p33_ASAP7_75t_R g411 ( .A(n_64), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_272), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_258), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_87), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_31), .Y(n_415) );
NOR2xp67_ASAP7_75t_L g416 ( .A(n_246), .B(n_80), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_44), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_135), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_111), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_261), .B(n_187), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_33), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_96), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_41), .Y(n_423) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_226), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_122), .Y(n_425) );
BUFx3_ASAP7_75t_L g426 ( .A(n_50), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_159), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_113), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_16), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_166), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_251), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_196), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_158), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_220), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_29), .Y(n_435) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_50), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_193), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_49), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_12), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_27), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_81), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_237), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_85), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_279), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_318), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_279), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_321), .B(n_322), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_318), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_312), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_383), .B(n_386), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_383), .Y(n_451) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_279), .Y(n_452) );
INVx6_ASAP7_75t_L g453 ( .A(n_279), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_318), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_311), .B(n_0), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_386), .B(n_0), .Y(n_456) );
OAI21x1_ASAP7_75t_L g457 ( .A1(n_277), .A2(n_125), .B(n_124), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_318), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_318), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_295), .B(n_1), .Y(n_460) );
INVx3_ASAP7_75t_L g461 ( .A(n_423), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_423), .B(n_2), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
CKINVDCx6p67_ASAP7_75t_R g464 ( .A(n_346), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_330), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_322), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_466) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_277), .A2(n_129), .B(n_126), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_330), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_287), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_287), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_292), .Y(n_471) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_332), .A2(n_7), .B1(n_3), .B2(n_5), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_292), .Y(n_473) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_325), .A2(n_133), .B(n_132), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_390), .B(n_8), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_359), .Y(n_476) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_330), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_330), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_278), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_332), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_359), .B(n_9), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_321), .B(n_10), .Y(n_482) );
INVx4_ASAP7_75t_L g483 ( .A(n_456), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_447), .B(n_391), .Y(n_486) );
OR2x6_ASAP7_75t_L g487 ( .A(n_480), .B(n_394), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_444), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_445), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_448), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_447), .B(n_357), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_448), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_481), .A2(n_296), .B1(n_299), .B2(n_282), .Y(n_494) );
INVx4_ASAP7_75t_L g495 ( .A(n_456), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_481), .A2(n_309), .B1(n_313), .B2(n_305), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_454), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_464), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_464), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_481), .A2(n_320), .B1(n_334), .B2(n_329), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_482), .B(n_324), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_450), .B(n_397), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_482), .B(n_324), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_449), .B(n_375), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_466), .A2(n_335), .B1(n_337), .B2(n_301), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_454), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_450), .B(n_424), .Y(n_507) );
AND3x2_ASAP7_75t_L g508 ( .A(n_456), .B(n_355), .C(n_307), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_458), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_472), .A2(n_385), .B1(n_408), .B2(n_363), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_461), .B(n_325), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g512 ( .A(n_462), .B(n_315), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_479), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_444), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_444), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_461), .B(n_333), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_462), .A2(n_404), .B1(n_300), .B2(n_316), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_449), .B(n_394), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_461), .B(n_333), .Y(n_520) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_460), .A2(n_385), .B1(n_408), .B2(n_363), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_458), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_519), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_494), .B(n_455), .C(n_475), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_501), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_513), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_501), .B(n_459), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_503), .A2(n_300), .B1(n_316), .B2(n_291), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_519), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_504), .B(n_459), .Y(n_530) );
INVx2_ASAP7_75t_SL g531 ( .A(n_504), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_486), .A2(n_369), .B1(n_373), .B2(n_291), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_492), .B(n_451), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_519), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_513), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_521), .B(n_350), .Y(n_537) );
OR2x6_ASAP7_75t_L g538 ( .A(n_498), .B(n_457), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_492), .B(n_463), .Y(n_539) );
INVx2_ASAP7_75t_SL g540 ( .A(n_508), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_517), .A2(n_516), .B(n_520), .C(n_511), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_518), .B(n_364), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_502), .A2(n_373), .B1(n_402), .B2(n_369), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_507), .A2(n_402), .B1(n_289), .B2(n_298), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_499), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_483), .B(n_434), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_517), .B(n_457), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_513), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_487), .A2(n_378), .B1(n_389), .B2(n_353), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_517), .B(n_304), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_505), .A2(n_351), .B1(n_358), .B2(n_285), .Y(n_551) );
AND2x4_ASAP7_75t_SL g552 ( .A(n_518), .B(n_319), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_519), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_512), .B(n_469), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g555 ( .A1(n_485), .A2(n_474), .B(n_467), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_508), .B(n_495), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_496), .A2(n_406), .B1(n_409), .B2(n_399), .C(n_396), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_505), .A2(n_380), .B1(n_407), .B2(n_384), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_495), .B(n_469), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_495), .B(n_470), .Y(n_560) );
INVx6_ASAP7_75t_L g561 ( .A(n_487), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_487), .A2(n_414), .B1(n_419), .B2(n_411), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_511), .Y(n_563) );
O2A1O1Ixp33_ASAP7_75t_L g564 ( .A1(n_510), .A2(n_473), .B(n_476), .C(n_471), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_510), .B(n_421), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_500), .B(n_516), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_520), .B(n_471), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_485), .B(n_361), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_489), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_490), .B(n_476), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_490), .B(n_372), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_493), .A2(n_417), .B(n_410), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_493), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_497), .B(n_413), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_506), .A2(n_422), .B1(n_440), .B2(n_425), .Y(n_575) );
XOR2xp5_ASAP7_75t_L g576 ( .A(n_506), .B(n_443), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_509), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_509), .B(n_467), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_522), .A2(n_319), .B1(n_429), .B2(n_428), .Y(n_579) );
AO22x1_ASAP7_75t_L g580 ( .A1(n_484), .A2(n_280), .B1(n_288), .B2(n_284), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_484), .B(n_306), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_488), .B(n_467), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_488), .A2(n_438), .B1(n_439), .B2(n_435), .Y(n_583) );
OR2x6_ASAP7_75t_L g584 ( .A(n_488), .B(n_400), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_491), .B(n_338), .Y(n_585) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_491), .A2(n_441), .B1(n_405), .B2(n_415), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_491), .B(n_381), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_514), .B(n_297), .Y(n_588) );
BUFx3_ASAP7_75t_L g589 ( .A(n_514), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_515), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_501), .B(n_302), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_569), .Y(n_592) );
INVx3_ASAP7_75t_L g593 ( .A(n_523), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_564), .A2(n_400), .B(n_415), .C(n_405), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_547), .A2(n_474), .B(n_367), .Y(n_595) );
NOR2xp33_ASAP7_75t_SL g596 ( .A(n_563), .B(n_420), .Y(n_596) );
NOR2xp67_ASAP7_75t_L g597 ( .A(n_535), .B(n_540), .Y(n_597) );
INVx3_ASAP7_75t_L g598 ( .A(n_529), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_547), .A2(n_474), .B(n_283), .Y(n_599) );
INVx4_ASAP7_75t_L g600 ( .A(n_556), .Y(n_600) );
AOI21xp33_ASAP7_75t_L g601 ( .A1(n_556), .A2(n_326), .B(n_314), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_578), .A2(n_474), .B(n_286), .Y(n_602) );
NOR2xp67_ASAP7_75t_SL g603 ( .A(n_561), .B(n_339), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_560), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_528), .B(n_345), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_578), .A2(n_290), .B(n_281), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_555), .A2(n_294), .B(n_293), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_565), .B(n_345), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_531), .B(n_352), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_525), .B(n_354), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_567), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_534), .B(n_377), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_561), .A2(n_416), .B1(n_303), .B2(n_310), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_544), .B(n_360), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_555), .A2(n_317), .B(n_308), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_561), .A2(n_368), .B1(n_376), .B2(n_345), .Y(n_617) );
INVx3_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
O2A1O1Ixp33_ASAP7_75t_SL g619 ( .A1(n_541), .A2(n_327), .B(n_328), .C(n_323), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_577), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_566), .B(n_388), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_559), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_562), .B(n_393), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_549), .A2(n_345), .B1(n_376), .B2(n_368), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_527), .Y(n_625) );
AOI21x1_ASAP7_75t_L g626 ( .A1(n_538), .A2(n_331), .B(n_343), .Y(n_626) );
AO21x1_ASAP7_75t_L g627 ( .A1(n_582), .A2(n_348), .B(n_347), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_584), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_552), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_530), .A2(n_365), .B(n_362), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_524), .A2(n_368), .B1(n_436), .B2(n_376), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_530), .A2(n_370), .B(n_366), .Y(n_632) );
AND2x4_ASAP7_75t_L g633 ( .A(n_533), .B(n_374), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_539), .B(n_379), .Y(n_634) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_545), .B(n_382), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_584), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_550), .A2(n_395), .B(n_392), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_557), .A2(n_401), .B(n_403), .C(n_398), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_570), .Y(n_639) );
BUFx2_ASAP7_75t_SL g640 ( .A(n_543), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_554), .A2(n_376), .B1(n_436), .B2(n_368), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_591), .B(n_418), .Y(n_642) );
BUFx4f_ASAP7_75t_L g643 ( .A(n_542), .Y(n_643) );
INVx2_ASAP7_75t_SL g644 ( .A(n_576), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_568), .Y(n_645) );
BUFx2_ASAP7_75t_L g646 ( .A(n_532), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_575), .B(n_430), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_568), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_537), .B(n_436), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_571), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_546), .A2(n_432), .B(n_427), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_551), .A2(n_433), .B1(n_437), .B2(n_431), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_586), .B(n_436), .C(n_340), .Y(n_653) );
BUFx8_ASAP7_75t_L g654 ( .A(n_526), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_584), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_579), .B(n_349), .C(n_340), .Y(n_656) );
NOR2xp33_ASAP7_75t_SL g657 ( .A(n_572), .B(n_349), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_571), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_574), .Y(n_659) );
BUFx10_ASAP7_75t_L g660 ( .A(n_581), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_536), .A2(n_341), .B(n_336), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_548), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g663 ( .A1(n_574), .A2(n_336), .B1(n_371), .B2(n_341), .Y(n_663) );
OR2x2_ASAP7_75t_L g664 ( .A(n_558), .B(n_11), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_580), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_583), .B(n_387), .Y(n_666) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_589), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_585), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_588), .A2(n_342), .B(n_278), .Y(n_669) );
CKINVDCx8_ASAP7_75t_R g670 ( .A(n_587), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_590), .A2(n_442), .B(n_412), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_524), .B(n_356), .C(n_344), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_SL g673 ( .A1(n_541), .A2(n_140), .B(n_141), .C(n_137), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_563), .A2(n_453), .B1(n_356), .B2(n_344), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_563), .B(n_13), .Y(n_675) );
BUFx6f_ASAP7_75t_L g676 ( .A(n_584), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_564), .A2(n_16), .B(n_14), .C(n_15), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_563), .B(n_15), .Y(n_678) );
CKINVDCx11_ASAP7_75t_R g679 ( .A(n_545), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_563), .B(n_18), .Y(n_680) );
NAND2x1p5_ASAP7_75t_L g681 ( .A(n_563), .B(n_344), .Y(n_681) );
NOR3xp33_ASAP7_75t_L g682 ( .A(n_564), .B(n_18), .C(n_19), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_563), .B(n_21), .Y(n_683) );
BUFx3_ASAP7_75t_L g684 ( .A(n_545), .Y(n_684) );
INVx1_ASAP7_75t_SL g685 ( .A(n_563), .Y(n_685) );
BUFx8_ASAP7_75t_L g686 ( .A(n_545), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_540), .B(n_22), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_560), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_563), .A2(n_452), .B1(n_465), .B2(n_446), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_563), .B(n_24), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_547), .A2(n_468), .B(n_465), .Y(n_691) );
BUFx12f_ASAP7_75t_L g692 ( .A(n_545), .Y(n_692) );
INVx5_ASAP7_75t_L g693 ( .A(n_676), .Y(n_693) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_595), .A2(n_468), .B(n_465), .Y(n_694) );
AOI221x1_ASAP7_75t_L g695 ( .A1(n_672), .A2(n_478), .B1(n_477), .B2(n_468), .C(n_29), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_602), .A2(n_477), .B(n_468), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_685), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_685), .Y(n_698) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_679), .Y(n_699) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_596), .A2(n_478), .B1(n_477), .B2(n_28), .Y(n_700) );
BUFx3_ASAP7_75t_L g701 ( .A(n_654), .Y(n_701) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_692), .B(n_25), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g703 ( .A1(n_599), .A2(n_478), .B(n_477), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_611), .B(n_26), .Y(n_704) );
AO31x2_ASAP7_75t_L g705 ( .A1(n_627), .A2(n_31), .A3(n_28), .B(n_30), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_611), .Y(n_706) );
BUFx12f_ASAP7_75t_L g707 ( .A(n_686), .Y(n_707) );
NAND3x1_ASAP7_75t_L g708 ( .A(n_635), .B(n_30), .C(n_32), .Y(n_708) );
AO31x2_ASAP7_75t_L g709 ( .A1(n_607), .A2(n_34), .A3(n_32), .B(n_33), .Y(n_709) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_645), .A2(n_650), .B(n_658), .C(n_648), .Y(n_710) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_667), .Y(n_711) );
AO31x2_ASAP7_75t_L g712 ( .A1(n_616), .A2(n_38), .A3(n_36), .B(n_37), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_659), .B(n_36), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_654), .Y(n_714) );
INVxp67_ASAP7_75t_L g715 ( .A(n_596), .Y(n_715) );
INVx2_ASAP7_75t_SL g716 ( .A(n_686), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g717 ( .A1(n_606), .A2(n_164), .B(n_161), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_643), .A2(n_42), .B1(n_40), .B2(n_41), .Y(n_718) );
AOI221xp5_ASAP7_75t_SL g719 ( .A1(n_613), .A2(n_42), .B1(n_43), .B2(n_45), .C(n_46), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_620), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_639), .B(n_47), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_630), .A2(n_49), .B(n_47), .C(n_48), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_640), .B(n_48), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_629), .B(n_52), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_684), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_600), .B(n_53), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_649), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_604), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_644), .B(n_56), .Y(n_729) );
INVxp67_ASAP7_75t_L g730 ( .A(n_597), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_632), .A2(n_170), .B(n_169), .Y(n_731) );
OAI21xp5_ASAP7_75t_L g732 ( .A1(n_672), .A2(n_175), .B(n_172), .Y(n_732) );
AO31x2_ASAP7_75t_L g733 ( .A1(n_691), .A2(n_57), .A3(n_58), .B(n_59), .Y(n_733) );
O2A1O1Ixp33_ASAP7_75t_SL g734 ( .A1(n_621), .A2(n_197), .B(n_276), .C(n_275), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_618), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_633), .B(n_58), .Y(n_736) );
AOI221xp5_ASAP7_75t_SL g737 ( .A1(n_613), .A2(n_60), .B1(n_61), .B2(n_63), .C(n_65), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_615), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_623), .A2(n_60), .B1(n_65), .B2(n_66), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_634), .B(n_66), .Y(n_740) );
BUFx10_ASAP7_75t_L g741 ( .A(n_676), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_600), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_614), .B(n_67), .Y(n_743) );
NAND3x1_ASAP7_75t_L g744 ( .A(n_682), .B(n_68), .C(n_69), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_688), .A2(n_70), .B1(n_72), .B2(n_73), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_622), .A2(n_72), .B1(n_74), .B2(n_75), .Y(n_746) );
INVx5_ASAP7_75t_L g747 ( .A(n_676), .Y(n_747) );
CKINVDCx11_ASAP7_75t_R g748 ( .A(n_670), .Y(n_748) );
AO21x1_ASAP7_75t_L g749 ( .A1(n_669), .A2(n_181), .B(n_180), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_L g750 ( .A1(n_594), .A2(n_77), .B(n_78), .C(n_79), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_608), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_675), .Y(n_752) );
BUFx2_ASAP7_75t_L g753 ( .A(n_628), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_628), .B(n_77), .Y(n_754) );
AO31x2_ASAP7_75t_L g755 ( .A1(n_674), .A2(n_78), .A3(n_79), .B(n_82), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_636), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_619), .A2(n_183), .B(n_182), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_638), .A2(n_83), .B1(n_84), .B2(n_85), .C(n_86), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g759 ( .A1(n_637), .A2(n_83), .B(n_84), .C(n_87), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_678), .A2(n_683), .B1(n_690), .B2(n_680), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_677), .A2(n_88), .B(n_90), .C(n_91), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_605), .B(n_88), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_592), .Y(n_763) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_667), .B(n_92), .Y(n_764) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_668), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_765) );
A2O1A1Ixp33_ASAP7_75t_L g766 ( .A1(n_661), .A2(n_93), .B(n_94), .C(n_95), .Y(n_766) );
O2A1O1Ixp33_ASAP7_75t_L g767 ( .A1(n_664), .A2(n_96), .B(n_98), .C(n_99), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_665), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_601), .Y(n_769) );
AOI221x1_ASAP7_75t_L g770 ( .A1(n_656), .A2(n_98), .B1(n_99), .B2(n_100), .C(n_101), .Y(n_770) );
BUFx2_ASAP7_75t_L g771 ( .A(n_636), .Y(n_771) );
INVx2_ASAP7_75t_SL g772 ( .A(n_647), .Y(n_772) );
OA21x2_ASAP7_75t_L g773 ( .A1(n_671), .A2(n_223), .B(n_271), .Y(n_773) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_667), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_655), .Y(n_775) );
INVx2_ASAP7_75t_L g776 ( .A(n_593), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_652), .B(n_101), .Y(n_777) );
NAND2x1p5_ASAP7_75t_L g778 ( .A(n_603), .B(n_102), .Y(n_778) );
AND2x4_ASAP7_75t_L g779 ( .A(n_598), .B(n_102), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_598), .B(n_103), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_651), .A2(n_104), .B(n_105), .C(n_106), .Y(n_781) );
AO31x2_ASAP7_75t_L g782 ( .A1(n_663), .A2(n_105), .A3(n_106), .B(n_107), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_660), .B(n_107), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_662), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_642), .B(n_108), .Y(n_785) );
BUFx6f_ASAP7_75t_L g786 ( .A(n_660), .Y(n_786) );
BUFx12f_ASAP7_75t_L g787 ( .A(n_612), .Y(n_787) );
O2A1O1Ixp33_ASAP7_75t_SL g788 ( .A1(n_666), .A2(n_219), .B(n_267), .C(n_266), .Y(n_788) );
NAND3xp33_ASAP7_75t_SL g789 ( .A(n_612), .B(n_109), .C(n_110), .Y(n_789) );
INVx3_ASAP7_75t_L g790 ( .A(n_609), .Y(n_790) );
O2A1O1Ixp33_ASAP7_75t_L g791 ( .A1(n_624), .A2(n_109), .B(n_112), .C(n_114), .Y(n_791) );
OAI21x1_ASAP7_75t_L g792 ( .A1(n_689), .A2(n_228), .B(n_262), .Y(n_792) );
OA21x2_ASAP7_75t_L g793 ( .A1(n_631), .A2(n_653), .B(n_641), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_687), .B(n_112), .Y(n_794) );
AO31x2_ASAP7_75t_L g795 ( .A1(n_617), .A2(n_114), .A3(n_115), .B(n_116), .Y(n_795) );
OAI21x1_ASAP7_75t_L g796 ( .A1(n_653), .A2(n_229), .B(n_260), .Y(n_796) );
AO31x2_ASAP7_75t_L g797 ( .A1(n_673), .A2(n_115), .A3(n_116), .B(n_117), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_610), .A2(n_215), .B(n_259), .Y(n_798) );
AO21x2_ASAP7_75t_L g799 ( .A1(n_657), .A2(n_214), .B(n_257), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_657), .Y(n_800) );
AO21x1_ASAP7_75t_L g801 ( .A1(n_607), .A2(n_213), .B(n_256), .Y(n_801) );
BUFx10_ASAP7_75t_L g802 ( .A(n_676), .Y(n_802) );
AO31x2_ASAP7_75t_L g803 ( .A1(n_627), .A2(n_117), .A3(n_118), .B(n_119), .Y(n_803) );
A2O1A1Ixp33_ASAP7_75t_L g804 ( .A1(n_645), .A2(n_118), .B(n_119), .C(n_120), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_595), .A2(n_230), .B(n_253), .Y(n_805) );
A2O1A1Ixp33_ASAP7_75t_L g806 ( .A1(n_645), .A2(n_121), .B(n_122), .C(n_184), .Y(n_806) );
BUFx2_ASAP7_75t_L g807 ( .A(n_685), .Y(n_807) );
INVx2_ASAP7_75t_SL g808 ( .A(n_654), .Y(n_808) );
AO31x2_ASAP7_75t_L g809 ( .A1(n_627), .A2(n_188), .A3(n_190), .B(n_192), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_644), .B(n_195), .Y(n_810) );
BUFx24_ASAP7_75t_L g811 ( .A(n_686), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_685), .Y(n_812) );
AOI31xp67_ASAP7_75t_L g813 ( .A1(n_689), .A2(n_200), .A3(n_203), .B(n_204), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_685), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_706), .B(n_206), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_720), .Y(n_816) );
OR2x2_ASAP7_75t_L g817 ( .A(n_807), .B(n_231), .Y(n_817) );
AO31x2_ASAP7_75t_L g818 ( .A1(n_801), .A2(n_232), .A3(n_233), .B(n_234), .Y(n_818) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_711), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_814), .B(n_238), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_710), .B(n_240), .Y(n_821) );
BUFx2_ASAP7_75t_L g822 ( .A(n_714), .Y(n_822) );
NAND2x1p5_ASAP7_75t_L g823 ( .A(n_701), .B(n_250), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_763), .Y(n_824) );
INVx4_ASAP7_75t_L g825 ( .A(n_707), .Y(n_825) );
AND2x4_ASAP7_75t_L g826 ( .A(n_786), .B(n_247), .Y(n_826) );
INVx3_ASAP7_75t_L g827 ( .A(n_741), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_697), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_698), .Y(n_829) );
BUFx2_ASAP7_75t_R g830 ( .A(n_699), .Y(n_830) );
INVx4_ASAP7_75t_L g831 ( .A(n_693), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_812), .Y(n_832) );
AO31x2_ASAP7_75t_L g833 ( .A1(n_800), .A2(n_749), .A3(n_770), .B(n_757), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_738), .Y(n_834) );
INVx4_ASAP7_75t_L g835 ( .A(n_693), .Y(n_835) );
AO31x2_ASAP7_75t_L g836 ( .A1(n_805), .A2(n_761), .A3(n_806), .B(n_750), .Y(n_836) );
OAI21x1_ASAP7_75t_SL g837 ( .A1(n_798), .A2(n_731), .B(n_717), .Y(n_837) );
OA21x2_ASAP7_75t_L g838 ( .A1(n_796), .A2(n_732), .B(n_792), .Y(n_838) );
CKINVDCx16_ASAP7_75t_R g839 ( .A(n_811), .Y(n_839) );
HB1xp67_ASAP7_75t_L g840 ( .A(n_725), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_715), .B(n_769), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_786), .B(n_790), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_721), .A2(n_713), .B(n_780), .Y(n_843) );
NAND2x1p5_ASAP7_75t_L g844 ( .A(n_808), .B(n_693), .Y(n_844) );
INVx2_ASAP7_75t_SL g845 ( .A(n_742), .Y(n_845) );
BUFx4_ASAP7_75t_SL g846 ( .A(n_768), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_751), .B(n_727), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_754), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_784), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_741), .Y(n_850) );
A2O1A1Ixp33_ASAP7_75t_L g851 ( .A1(n_743), .A2(n_723), .B(n_767), .C(n_791), .Y(n_851) );
BUFx3_ASAP7_75t_L g852 ( .A(n_716), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_772), .B(n_729), .Y(n_853) );
NAND2xp5_ASAP7_75t_SL g854 ( .A(n_779), .B(n_747), .Y(n_854) );
OR2x2_ASAP7_75t_L g855 ( .A(n_736), .B(n_740), .Y(n_855) );
BUFx3_ASAP7_75t_L g856 ( .A(n_787), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_704), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_752), .A2(n_773), .B(n_734), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_728), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_733), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_745), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_810), .B(n_724), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_733), .Y(n_863) );
INVx2_ASAP7_75t_L g864 ( .A(n_733), .Y(n_864) );
INVx2_ASAP7_75t_SL g865 ( .A(n_802), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_782), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_747), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_775), .B(n_777), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_782), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_744), .A2(n_700), .B1(n_778), .B2(n_739), .Y(n_870) );
INVx1_ASAP7_75t_SL g871 ( .A(n_802), .Y(n_871) );
AOI21xp5_ASAP7_75t_L g872 ( .A1(n_794), .A2(n_793), .B(n_788), .Y(n_872) );
AOI21xp5_ASAP7_75t_L g873 ( .A1(n_793), .A2(n_762), .B(n_776), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_726), .A2(n_783), .B1(n_789), .B2(n_758), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_782), .Y(n_875) );
BUFx3_ASAP7_75t_L g876 ( .A(n_748), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_747), .Y(n_877) );
AOI21xp5_ASAP7_75t_L g878 ( .A1(n_735), .A2(n_785), .B(n_764), .Y(n_878) );
NAND2xp5_ASAP7_75t_SL g879 ( .A(n_702), .B(n_730), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_756), .B(n_753), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_709), .Y(n_881) );
NAND2x1p5_ASAP7_75t_L g882 ( .A(n_771), .B(n_718), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_719), .B(n_737), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_709), .Y(n_884) );
INVxp67_ASAP7_75t_SL g885 ( .A(n_774), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_722), .B(n_759), .Y(n_886) );
NAND2x1p5_ASAP7_75t_L g887 ( .A(n_765), .B(n_746), .Y(n_887) );
NAND2x1p5_ASAP7_75t_L g888 ( .A(n_708), .B(n_804), .Y(n_888) );
AOI21x1_ASAP7_75t_L g889 ( .A1(n_813), .A2(n_797), .B(n_809), .Y(n_889) );
OAI21x1_ASAP7_75t_L g890 ( .A1(n_799), .A2(n_797), .B(n_809), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_781), .B(n_705), .Y(n_891) );
INVx6_ASAP7_75t_L g892 ( .A(n_766), .Y(n_892) );
AO31x2_ASAP7_75t_L g893 ( .A1(n_797), .A2(n_809), .A3(n_803), .B(n_705), .Y(n_893) );
OR2x6_ASAP7_75t_L g894 ( .A(n_795), .B(n_709), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_803), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_705), .B(n_803), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_712), .B(n_795), .Y(n_897) );
OAI21x1_ASAP7_75t_L g898 ( .A1(n_712), .A2(n_755), .B(n_795), .Y(n_898) );
OA21x2_ASAP7_75t_L g899 ( .A1(n_755), .A2(n_694), .B(n_696), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_755), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_699), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_706), .Y(n_902) );
BUFx3_ASAP7_75t_L g903 ( .A(n_701), .Y(n_903) );
AOI21x1_ASAP7_75t_L g904 ( .A1(n_694), .A2(n_626), .B(n_696), .Y(n_904) );
OAI21x1_ASAP7_75t_SL g905 ( .A1(n_798), .A2(n_731), .B(n_717), .Y(n_905) );
BUFx4f_ASAP7_75t_L g906 ( .A(n_707), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_710), .B(n_625), .Y(n_907) );
AOI21xp33_ASAP7_75t_SL g908 ( .A1(n_715), .A2(n_811), .B(n_808), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_706), .B(n_685), .Y(n_909) );
OAI21x1_ASAP7_75t_L g910 ( .A1(n_694), .A2(n_696), .B(n_703), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_710), .B(n_625), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_720), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_720), .Y(n_913) );
INVx4_ASAP7_75t_L g914 ( .A(n_707), .Y(n_914) );
NAND2x1p5_ASAP7_75t_L g915 ( .A(n_701), .B(n_714), .Y(n_915) );
BUFx2_ASAP7_75t_L g916 ( .A(n_714), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g917 ( .A(n_710), .B(n_625), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_706), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_706), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_720), .Y(n_920) );
AO21x1_ASAP7_75t_L g921 ( .A1(n_760), .A2(n_800), .B(n_681), .Y(n_921) );
NAND2xp5_ASAP7_75t_SL g922 ( .A(n_715), .B(n_685), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_710), .B(n_625), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_706), .Y(n_924) );
BUFx2_ASAP7_75t_L g925 ( .A(n_714), .Y(n_925) );
AO31x2_ASAP7_75t_L g926 ( .A1(n_801), .A2(n_627), .A3(n_695), .B(n_800), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_706), .B(n_685), .Y(n_927) );
NAND3xp33_ASAP7_75t_L g928 ( .A(n_770), .B(n_737), .C(n_719), .Y(n_928) );
CKINVDCx11_ASAP7_75t_R g929 ( .A(n_707), .Y(n_929) );
OAI21x1_ASAP7_75t_SL g930 ( .A1(n_798), .A2(n_731), .B(n_717), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_706), .Y(n_931) );
AO31x2_ASAP7_75t_L g932 ( .A1(n_801), .A2(n_627), .A3(n_695), .B(n_800), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_694), .A2(n_595), .B(n_696), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_710), .B(n_625), .Y(n_934) );
OAI21x1_ASAP7_75t_SL g935 ( .A1(n_798), .A2(n_731), .B(n_717), .Y(n_935) );
INVx6_ASAP7_75t_L g936 ( .A(n_707), .Y(n_936) );
CKINVDCx11_ASAP7_75t_R g937 ( .A(n_707), .Y(n_937) );
INVx4_ASAP7_75t_SL g938 ( .A(n_707), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_706), .B(n_685), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_706), .Y(n_940) );
AOI21x1_ASAP7_75t_L g941 ( .A1(n_694), .A2(n_626), .B(n_696), .Y(n_941) );
BUFx2_ASAP7_75t_SL g942 ( .A(n_856), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_909), .B(n_927), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_834), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_939), .B(n_912), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_840), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_913), .B(n_920), .Y(n_947) );
OR2x6_ASAP7_75t_L g948 ( .A(n_854), .B(n_823), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_816), .Y(n_949) );
BUFx6f_ASAP7_75t_L g950 ( .A(n_819), .Y(n_950) );
BUFx2_ASAP7_75t_L g951 ( .A(n_839), .Y(n_951) );
INVx1_ASAP7_75t_L g952 ( .A(n_902), .Y(n_952) );
AO21x2_ASAP7_75t_L g953 ( .A1(n_889), .A2(n_897), .B(n_837), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_822), .B(n_916), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_918), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_824), .B(n_849), .Y(n_956) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_925), .B(n_868), .Y(n_957) );
BUFx3_ASAP7_75t_L g958 ( .A(n_915), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_896), .B(n_866), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_919), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_924), .B(n_931), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_940), .Y(n_962) );
AO21x2_ASAP7_75t_L g963 ( .A1(n_897), .A2(n_930), .B(n_905), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g964 ( .A1(n_839), .A2(n_870), .B1(n_892), .B2(n_888), .Y(n_964) );
BUFx2_ASAP7_75t_L g965 ( .A(n_844), .Y(n_965) );
AO21x2_ASAP7_75t_L g966 ( .A1(n_935), .A2(n_872), .B(n_891), .Y(n_966) );
OA21x2_ASAP7_75t_L g967 ( .A1(n_890), .A2(n_898), .B(n_873), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_859), .B(n_861), .Y(n_968) );
INVx2_ASAP7_75t_SL g969 ( .A(n_842), .Y(n_969) );
AO21x2_ASAP7_75t_L g970 ( .A1(n_891), .A2(n_933), .B(n_869), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_828), .Y(n_971) );
CKINVDCx10_ASAP7_75t_R g972 ( .A(n_906), .Y(n_972) );
INVxp67_ASAP7_75t_SL g973 ( .A(n_880), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_887), .A2(n_870), .B1(n_874), .B2(n_892), .Y(n_974) );
BUFx3_ASAP7_75t_L g975 ( .A(n_903), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_829), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_832), .B(n_857), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_847), .B(n_895), .Y(n_978) );
BUFx12f_ASAP7_75t_L g979 ( .A(n_929), .Y(n_979) );
OR2x6_ASAP7_75t_L g980 ( .A(n_882), .B(n_831), .Y(n_980) );
INVx6_ASAP7_75t_L g981 ( .A(n_938), .Y(n_981) );
INVx3_ASAP7_75t_L g982 ( .A(n_831), .Y(n_982) );
INVxp67_ASAP7_75t_SL g983 ( .A(n_880), .Y(n_983) );
INVx3_ASAP7_75t_L g984 ( .A(n_835), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_894), .B(n_907), .Y(n_985) );
OA21x2_ASAP7_75t_L g986 ( .A1(n_860), .A2(n_863), .B(n_864), .Y(n_986) );
OA21x2_ASAP7_75t_L g987 ( .A1(n_881), .A2(n_884), .B(n_875), .Y(n_987) );
BUFx3_ASAP7_75t_L g988 ( .A(n_906), .Y(n_988) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_900), .A2(n_921), .B(n_858), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_894), .B(n_907), .Y(n_990) );
BUFx4f_ASAP7_75t_SL g991 ( .A(n_825), .Y(n_991) );
INVx2_ASAP7_75t_SL g992 ( .A(n_835), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_848), .Y(n_993) );
BUFx6f_ASAP7_75t_L g994 ( .A(n_910), .Y(n_994) );
OR2x6_ASAP7_75t_L g995 ( .A(n_911), .B(n_917), .Y(n_995) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_867), .Y(n_996) );
OR2x2_ASAP7_75t_L g997 ( .A(n_894), .B(n_883), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_922), .Y(n_998) );
AND2x2_ASAP7_75t_L g999 ( .A(n_923), .B(n_934), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_817), .Y(n_1000) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_885), .Y(n_1001) );
AND2x4_ASAP7_75t_L g1002 ( .A(n_877), .B(n_923), .Y(n_1002) );
INVx4_ASAP7_75t_L g1003 ( .A(n_827), .Y(n_1003) );
OAI21xp5_ASAP7_75t_L g1004 ( .A1(n_851), .A2(n_928), .B(n_843), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_871), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1006 ( .A(n_883), .B(n_855), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_934), .B(n_893), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_826), .Y(n_1008) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_852), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_862), .A2(n_908), .B1(n_928), .B2(n_886), .Y(n_1010) );
AO21x2_ASAP7_75t_L g1011 ( .A1(n_843), .A2(n_941), .B(n_904), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_871), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_899), .Y(n_1013) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_827), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_826), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1016 ( .A(n_937), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_820), .Y(n_1017) );
AND2x4_ASAP7_75t_L g1018 ( .A(n_815), .B(n_878), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_893), .B(n_886), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_893), .B(n_836), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_850), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_865), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_836), .B(n_899), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_938), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_836), .B(n_821), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_846), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_845), .Y(n_1027) );
HB1xp67_ASAP7_75t_L g1028 ( .A(n_853), .Y(n_1028) );
OR2x6_ASAP7_75t_L g1029 ( .A(n_879), .B(n_841), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_833), .B(n_932), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_818), .Y(n_1031) );
AO21x2_ASAP7_75t_L g1032 ( .A1(n_833), .A2(n_926), .B(n_838), .Y(n_1032) );
INVx2_ASAP7_75t_L g1033 ( .A(n_833), .Y(n_1033) );
INVx2_ASAP7_75t_L g1034 ( .A(n_936), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_825), .B(n_914), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_936), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_876), .Y(n_1037) );
AND2x4_ASAP7_75t_L g1038 ( .A(n_914), .B(n_901), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_830), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_830), .B(n_646), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_909), .B(n_939), .Y(n_1041) );
BUFx3_ASAP7_75t_L g1042 ( .A(n_965), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_959), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_978), .B(n_968), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_1001), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_959), .Y(n_1046) );
OR2x2_ASAP7_75t_L g1047 ( .A(n_973), .B(n_983), .Y(n_1047) );
INVx4_ASAP7_75t_L g1048 ( .A(n_980), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_943), .B(n_1041), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_987), .Y(n_1050) );
INVxp67_ASAP7_75t_L g1051 ( .A(n_942), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_943), .B(n_1041), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_946), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_985), .B(n_990), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_997), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_1005), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_1013), .Y(n_1057) );
AND2x2_ASAP7_75t_L g1058 ( .A(n_990), .B(n_1019), .Y(n_1058) );
AND2x2_ASAP7_75t_SL g1059 ( .A(n_951), .B(n_1024), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_945), .B(n_1020), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_986), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1020), .B(n_1007), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_1007), .B(n_1004), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1023), .B(n_999), .Y(n_1064) );
BUFx3_ASAP7_75t_L g1065 ( .A(n_958), .Y(n_1065) );
INVx1_ASAP7_75t_L g1066 ( .A(n_944), .Y(n_1066) );
NOR2x1_ASAP7_75t_L g1067 ( .A(n_1003), .B(n_982), .Y(n_1067) );
INVxp67_ASAP7_75t_L g1068 ( .A(n_996), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1023), .B(n_999), .Y(n_1069) );
INVx1_ASAP7_75t_SL g1070 ( .A(n_975), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1071 ( .A(n_1012), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_947), .B(n_961), .Y(n_1072) );
INVx6_ASAP7_75t_L g1073 ( .A(n_981), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_949), .Y(n_1074) );
INVx5_ASAP7_75t_L g1075 ( .A(n_980), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_1002), .B(n_1018), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_952), .Y(n_1077) );
CKINVDCx11_ASAP7_75t_R g1078 ( .A(n_979), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_955), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_970), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_956), .B(n_977), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_974), .A2(n_964), .B1(n_1010), .B2(n_1028), .Y(n_1082) );
CKINVDCx6p67_ASAP7_75t_R g1083 ( .A(n_972), .Y(n_1083) );
INVxp33_ASAP7_75t_L g1084 ( .A(n_1026), .Y(n_1084) );
AND2x4_ASAP7_75t_L g1085 ( .A(n_1002), .B(n_1018), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_995), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1087 ( .A(n_1014), .Y(n_1087) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_950), .Y(n_1088) );
INVxp67_ASAP7_75t_L g1089 ( .A(n_954), .Y(n_1089) );
INVxp67_ASAP7_75t_L g1090 ( .A(n_1009), .Y(n_1090) );
INVx4_ASAP7_75t_L g1091 ( .A(n_980), .Y(n_1091) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_1018), .B(n_1008), .Y(n_1092) );
NOR2xp67_ASAP7_75t_L g1093 ( .A(n_1003), .B(n_992), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1006), .B(n_995), .Y(n_1094) );
AND2x2_ASAP7_75t_L g1095 ( .A(n_995), .B(n_1030), .Y(n_1095) );
BUFx3_ASAP7_75t_L g1096 ( .A(n_958), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1030), .B(n_1025), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1025), .B(n_960), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1049), .B(n_962), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1100 ( .A(n_1045), .Y(n_1100) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1050), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_1057), .Y(n_1102) );
AND2x4_ASAP7_75t_L g1103 ( .A(n_1076), .B(n_963), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1066), .Y(n_1104) );
NAND2x1p5_ASAP7_75t_L g1105 ( .A(n_1075), .B(n_984), .Y(n_1105) );
INVx1_ASAP7_75t_L g1106 ( .A(n_1074), .Y(n_1106) );
INVxp67_ASAP7_75t_L g1107 ( .A(n_1053), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1062), .B(n_963), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1097), .B(n_953), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1077), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1097), .B(n_953), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1079), .Y(n_1112) );
INVxp67_ASAP7_75t_L g1113 ( .A(n_1087), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_1064), .B(n_953), .Y(n_1114) );
AOI22xp5_ASAP7_75t_SL g1115 ( .A1(n_1051), .A2(n_1016), .B1(n_1038), .B2(n_988), .Y(n_1115) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_1067), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1064), .B(n_1011), .Y(n_1117) );
NAND3xp33_ASAP7_75t_L g1118 ( .A(n_1082), .B(n_957), .C(n_998), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1049), .B(n_971), .Y(n_1119) );
AND2x4_ASAP7_75t_L g1120 ( .A(n_1076), .B(n_1011), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1060), .B(n_1033), .Y(n_1121) );
NOR2xp33_ASAP7_75t_L g1122 ( .A(n_1084), .B(n_1036), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1069), .B(n_966), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1058), .B(n_966), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1063), .B(n_1032), .Y(n_1125) );
AND2x4_ASAP7_75t_L g1126 ( .A(n_1076), .B(n_994), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1093), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1063), .B(n_1032), .Y(n_1128) );
INVx1_ASAP7_75t_SL g1129 ( .A(n_1070), .Y(n_1129) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_1052), .B(n_976), .Y(n_1130) );
INVxp67_ASAP7_75t_L g1131 ( .A(n_1056), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1098), .B(n_1032), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1044), .B(n_1031), .Y(n_1133) );
AND3x1_ASAP7_75t_L g1134 ( .A(n_1078), .B(n_1039), .C(n_1035), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1054), .B(n_967), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1095), .B(n_967), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1095), .B(n_967), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g1138 ( .A(n_1047), .Y(n_1138) );
BUFx2_ASAP7_75t_SL g1139 ( .A(n_1075), .Y(n_1139) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1072), .B(n_989), .Y(n_1140) );
BUFx2_ASAP7_75t_L g1141 ( .A(n_1088), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1072), .B(n_989), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_1071), .Y(n_1143) );
INVx3_ASAP7_75t_L g1144 ( .A(n_1048), .Y(n_1144) );
INVx4_ASAP7_75t_L g1145 ( .A(n_1105), .Y(n_1145) );
INVxp67_ASAP7_75t_L g1146 ( .A(n_1100), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1101), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1121), .B(n_1055), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1117), .B(n_1085), .Y(n_1149) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1102), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1101), .Y(n_1151) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1102), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1117), .B(n_1085), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1154 ( .A(n_1120), .B(n_1085), .Y(n_1154) );
OR2x6_ASAP7_75t_L g1155 ( .A(n_1139), .B(n_1048), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1109), .B(n_1086), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1111), .B(n_1086), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1111), .B(n_1092), .Y(n_1158) );
NOR2xp33_ASAP7_75t_L g1159 ( .A(n_1129), .B(n_1034), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1125), .B(n_1043), .Y(n_1160) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_1138), .Y(n_1161) );
INVx1_ASAP7_75t_SL g1162 ( .A(n_1141), .Y(n_1162) );
INVx2_ASAP7_75t_SL g1163 ( .A(n_1127), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1128), .B(n_1046), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1165 ( .A(n_1120), .B(n_1080), .Y(n_1165) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1115), .B(n_1034), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1124), .B(n_1081), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1123), .B(n_1061), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1128), .B(n_1094), .Y(n_1169) );
HB1xp67_ASAP7_75t_L g1170 ( .A(n_1143), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1171 ( .A(n_1107), .B(n_1037), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1167), .B(n_1168), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1147), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1150), .Y(n_1174) );
INVx3_ASAP7_75t_L g1175 ( .A(n_1145), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1147), .Y(n_1176) );
BUFx2_ASAP7_75t_L g1177 ( .A(n_1145), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1161), .Y(n_1178) );
NOR2x1_ASAP7_75t_L g1179 ( .A(n_1145), .B(n_1139), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1151), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1168), .B(n_1136), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1151), .Y(n_1182) );
INVx1_ASAP7_75t_SL g1183 ( .A(n_1170), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1156), .B(n_1136), .Y(n_1184) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1150), .Y(n_1185) );
AOI22xp5_ASAP7_75t_L g1186 ( .A1(n_1166), .A2(n_1118), .B1(n_1140), .B2(n_1142), .Y(n_1186) );
AOI221xp5_ASAP7_75t_L g1187 ( .A1(n_1146), .A2(n_1131), .B1(n_1113), .B2(n_1068), .C(n_1089), .Y(n_1187) );
AO21x1_ASAP7_75t_L g1188 ( .A1(n_1171), .A2(n_1106), .B(n_1104), .Y(n_1188) );
AND2x2_ASAP7_75t_SL g1189 ( .A(n_1154), .B(n_1059), .Y(n_1189) );
AO21x1_ASAP7_75t_L g1190 ( .A1(n_1159), .A2(n_1112), .B(n_1110), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1156), .B(n_1137), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1157), .B(n_1137), .Y(n_1192) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1169), .B(n_1132), .Y(n_1193) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1150), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1152), .Y(n_1195) );
NOR2x1_ASAP7_75t_L g1196 ( .A(n_1155), .B(n_1116), .Y(n_1196) );
AND2x4_ASAP7_75t_L g1197 ( .A(n_1165), .B(n_1120), .Y(n_1197) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_1162), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1152), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1172), .B(n_1157), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1173), .Y(n_1201) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1193), .B(n_1160), .Y(n_1202) );
OAI21xp5_ASAP7_75t_SL g1203 ( .A1(n_1177), .A2(n_1105), .B(n_1116), .Y(n_1203) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_1189), .A2(n_1155), .B1(n_1163), .B2(n_1091), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g1205 ( .A1(n_1189), .A2(n_1155), .B1(n_1163), .B2(n_1091), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1176), .Y(n_1206) );
INVx1_ASAP7_75t_SL g1207 ( .A(n_1183), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1180), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1180), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1182), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1186), .B(n_1164), .Y(n_1211) );
OAI211xp5_ASAP7_75t_L g1212 ( .A1(n_1177), .A2(n_1040), .B(n_1162), .C(n_1122), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1178), .B(n_1164), .Y(n_1213) );
OAI22xp33_ASAP7_75t_SL g1214 ( .A1(n_1175), .A2(n_1155), .B1(n_981), .B2(n_1105), .Y(n_1214) );
AOI222xp33_ASAP7_75t_L g1215 ( .A1(n_1187), .A2(n_1119), .B1(n_1130), .B2(n_1099), .C1(n_1090), .C2(n_1108), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1193), .B(n_1148), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1182), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_1188), .A2(n_1154), .B1(n_1165), .B2(n_1134), .Y(n_1218) );
INVx1_ASAP7_75t_SL g1219 ( .A(n_1175), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1211), .B(n_1181), .Y(n_1220) );
OAI211xp5_ASAP7_75t_L g1221 ( .A1(n_1218), .A2(n_1179), .B(n_1175), .C(n_1196), .Y(n_1221) );
AOI222xp33_ASAP7_75t_L g1222 ( .A1(n_1207), .A2(n_1198), .B1(n_1181), .B2(n_1184), .C1(n_1192), .C2(n_1191), .Y(n_1222) );
NAND2xp5_ASAP7_75t_SL g1223 ( .A(n_1214), .B(n_1190), .Y(n_1223) );
NOR2xp33_ASAP7_75t_L g1224 ( .A(n_1213), .B(n_1083), .Y(n_1224) );
AOI21xp5_ASAP7_75t_L g1225 ( .A1(n_1203), .A2(n_1212), .B(n_1205), .Y(n_1225) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_1215), .A2(n_1197), .B1(n_1103), .B2(n_1154), .Y(n_1226) );
O2A1O1Ixp33_ASAP7_75t_L g1227 ( .A1(n_1204), .A2(n_1038), .B(n_1027), .C(n_988), .Y(n_1227) );
AOI321xp33_ASAP7_75t_L g1228 ( .A1(n_1216), .A2(n_1108), .A3(n_1165), .B1(n_1123), .B2(n_1114), .C(n_1133), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1202), .B(n_1149), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1200), .B(n_1153), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_1219), .A2(n_1154), .B1(n_1048), .B2(n_1075), .Y(n_1231) );
O2A1O1Ixp33_ASAP7_75t_L g1232 ( .A1(n_1216), .A2(n_1038), .B(n_1022), .C(n_1021), .Y(n_1232) );
A2O1A1Ixp33_ASAP7_75t_L g1233 ( .A1(n_1201), .A2(n_1042), .B(n_1096), .C(n_1065), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_1206), .A2(n_1103), .B1(n_1165), .B2(n_1114), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1208), .Y(n_1235) );
OA21x2_ASAP7_75t_L g1236 ( .A1(n_1209), .A2(n_1185), .B(n_1174), .Y(n_1236) );
O2A1O1Ixp5_ASAP7_75t_L g1237 ( .A1(n_1210), .A2(n_1199), .B(n_1174), .C(n_1195), .Y(n_1237) );
NAND4xp25_ASAP7_75t_L g1238 ( .A(n_1217), .B(n_1096), .C(n_1065), .D(n_975), .Y(n_1238) );
A2O1A1Ixp33_ASAP7_75t_L g1239 ( .A1(n_1203), .A2(n_1042), .B(n_1144), .C(n_1075), .Y(n_1239) );
AOI22xp5_ASAP7_75t_L g1240 ( .A1(n_1215), .A2(n_1158), .B1(n_1133), .B2(n_1103), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1216), .Y(n_1241) );
NOR2x1_ASAP7_75t_L g1242 ( .A(n_1221), .B(n_1223), .Y(n_1242) );
INVxp33_ASAP7_75t_L g1243 ( .A(n_1224), .Y(n_1243) );
NAND4xp25_ASAP7_75t_SL g1244 ( .A(n_1226), .B(n_1225), .C(n_1240), .D(n_1222), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1241), .B(n_1229), .Y(n_1245) );
NAND3xp33_ASAP7_75t_SL g1246 ( .A(n_1016), .B(n_1232), .C(n_1227), .Y(n_1246) );
NOR2xp67_ASAP7_75t_L g1247 ( .A(n_979), .B(n_1231), .Y(n_1247) );
NOR3x1_ASAP7_75t_L g1248 ( .A(n_1238), .B(n_1220), .C(n_991), .Y(n_1248) );
OAI211xp5_ASAP7_75t_L g1249 ( .A1(n_1239), .A2(n_1228), .B(n_1234), .C(n_1233), .Y(n_1249) );
INVx2_ASAP7_75t_L g1250 ( .A(n_1248), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1243), .B(n_1230), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1252 ( .A(n_1244), .B(n_1235), .Y(n_1252) );
NAND3xp33_ASAP7_75t_SL g1253 ( .A(n_1249), .B(n_1237), .C(n_981), .Y(n_1253) );
NAND5xp2_ASAP7_75t_L g1254 ( .A(n_1242), .B(n_1000), .C(n_1017), .D(n_1015), .E(n_1073), .Y(n_1254) );
AOI21xp5_ASAP7_75t_SL g1255 ( .A1(n_1253), .A2(n_1246), .B(n_1247), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1251), .B(n_1245), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1250), .B(n_1236), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1252), .B(n_1029), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1257), .Y(n_1259) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1256), .Y(n_1260) );
XOR2xp5_ASAP7_75t_L g1261 ( .A(n_1258), .B(n_1254), .Y(n_1261) );
AOI22xp5_ASAP7_75t_L g1262 ( .A1(n_1259), .A2(n_1255), .B1(n_1073), .B2(n_1029), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1260), .Y(n_1263) );
AOI22x1_ASAP7_75t_SL g1264 ( .A1(n_1263), .A2(n_1261), .B1(n_984), .B2(n_993), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g1265 ( .A1(n_1262), .A2(n_1029), .B1(n_948), .B2(n_1075), .Y(n_1265) );
XNOR2xp5_ASAP7_75t_L g1266 ( .A(n_1264), .B(n_948), .Y(n_1266) );
NAND2xp5_ASAP7_75t_SL g1267 ( .A(n_1266), .B(n_1265), .Y(n_1267) );
AO221x2_ASAP7_75t_L g1268 ( .A1(n_1267), .A2(n_1199), .B1(n_1195), .B2(n_1194), .C(n_1185), .Y(n_1268) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_1268), .A2(n_969), .B1(n_1126), .B2(n_1135), .Y(n_1269) );
endmodule