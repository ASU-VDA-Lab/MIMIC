module fake_jpeg_32090_n_543 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_543);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_543;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_54),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_69),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_70),
.B(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_72),
.Y(n_156)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_100),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_94),
.Y(n_162)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_19),
.B(n_1),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_20),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_96),
.B(n_101),
.Y(n_166)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_98),
.Y(n_157)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_20),
.B(n_1),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_61),
.A2(n_75),
.B1(n_69),
.B2(n_58),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_107),
.A2(n_148),
.B1(n_165),
.B2(n_84),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_62),
.A2(n_49),
.B1(n_36),
.B2(n_33),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_124),
.A2(n_23),
.B1(n_36),
.B2(n_33),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_53),
.B(n_21),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_22),
.Y(n_168)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_151),
.Y(n_173)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_91),
.Y(n_137)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_52),
.A2(n_47),
.B1(n_49),
.B2(n_24),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_21),
.B1(n_50),
.B2(n_39),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_35),
.B1(n_22),
.B2(n_50),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_154),
.Y(n_216)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_59),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_164),
.Y(n_190)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_60),
.Y(n_161)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_85),
.A2(n_47),
.B1(n_33),
.B2(n_49),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_104),
.A2(n_85),
.B1(n_82),
.B2(n_83),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_168),
.B(n_185),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_169),
.A2(n_179),
.B1(n_202),
.B2(n_221),
.Y(n_276)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_80),
.B1(n_83),
.B2(n_68),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_177),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_111),
.A2(n_57),
.B1(n_68),
.B2(n_27),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_171),
.Y(n_272)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_172),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_105),
.A2(n_27),
.B(n_29),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_4),
.Y(n_237)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_178),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_136),
.A2(n_57),
.B1(n_25),
.B2(n_51),
.Y(n_179)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_181),
.Y(n_280)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_140),
.Y(n_182)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_121),
.Y(n_184)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_39),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_35),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_194),
.Y(n_251)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_80),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_217),
.Y(n_246)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_25),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_193),
.Y(n_241)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_29),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_133),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_64),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_195),
.B(n_203),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_196),
.Y(n_242)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_132),
.A2(n_81),
.B1(n_79),
.B2(n_78),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_200),
.A2(n_226),
.B1(n_134),
.B2(n_147),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_123),
.A2(n_51),
.B1(n_30),
.B2(n_49),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_30),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_113),
.A2(n_2),
.B(n_3),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_204),
.A2(n_4),
.B(n_5),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_113),
.B(n_49),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_205),
.B(n_211),
.Y(n_278)
);

INVx5_ASAP7_75t_SL g206 ( 
.A(n_117),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_206),
.Y(n_258)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_158),
.A2(n_72),
.B1(n_23),
.B2(n_33),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_215),
.B1(n_223),
.B2(n_115),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_36),
.Y(n_211)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_159),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_105),
.B(n_36),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_225),
.Y(n_257)
);

NAND2xp33_ASAP7_75t_SL g217 ( 
.A(n_114),
.B(n_36),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_112),
.B(n_33),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_107),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_115),
.A2(n_116),
.B1(n_125),
.B2(n_156),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_124),
.A2(n_23),
.B1(n_3),
.B2(n_4),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_224),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_122),
.B(n_2),
.Y(n_225)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_165),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_232),
.A2(n_226),
.B(n_174),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_233),
.B(n_226),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_237),
.B(n_252),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_157),
.B(n_127),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_244),
.A2(n_268),
.B(n_215),
.Y(n_312)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_245),
.A2(n_265),
.B1(n_208),
.B2(n_172),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_157),
.C(n_139),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_248),
.B(n_233),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_206),
.A2(n_134),
.B1(n_116),
.B2(n_125),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_249),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_190),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_255),
.B(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_256),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_169),
.A2(n_139),
.B1(n_147),
.B2(n_145),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_259),
.A2(n_263),
.B1(n_279),
.B2(n_210),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_156),
.B1(n_145),
.B2(n_138),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_264),
.A2(n_174),
.B1(n_186),
.B2(n_227),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_188),
.A2(n_138),
.B(n_120),
.C(n_7),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_173),
.B(n_5),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_269),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_220),
.A2(n_5),
.B(n_6),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_220),
.B(n_7),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_170),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_218),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_181),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_281),
.B(n_282),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g282 ( 
.A(n_258),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_247),
.A2(n_192),
.B1(n_182),
.B2(n_213),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g340 ( 
.A1(n_283),
.A2(n_310),
.B1(n_328),
.B2(n_253),
.Y(n_340)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_240),
.Y(n_284)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

CKINVDCx10_ASAP7_75t_R g285 ( 
.A(n_238),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_285),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_309),
.B1(n_246),
.B2(n_265),
.Y(n_333)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_228),
.B(n_217),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_287),
.B(n_291),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_242),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_240),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_289),
.Y(n_360)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_290),
.B(n_292),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g291 ( 
.A(n_228),
.B(n_170),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_254),
.B(n_197),
.Y(n_292)
);

AND2x6_ASAP7_75t_L g293 ( 
.A(n_228),
.B(n_170),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_293),
.B(n_299),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_295),
.A2(n_8),
.B(n_10),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_175),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_241),
.B(n_262),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_230),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_300),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_230),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_303),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_304),
.A2(n_245),
.B1(n_248),
.B2(n_236),
.Y(n_334)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_305),
.B(n_306),
.Y(n_353)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_212),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_316),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_308),
.B(n_324),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_272),
.A2(n_247),
.B1(n_276),
.B2(n_263),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_272),
.A2(n_183),
.B1(n_198),
.B2(n_199),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_314),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_312),
.A2(n_232),
.B(n_269),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_313),
.Y(n_358)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_315),
.A2(n_318),
.B1(n_327),
.B2(n_243),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_257),
.B(n_212),
.Y(n_316)
);

BUFx4f_ASAP7_75t_SL g317 ( 
.A(n_271),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_231),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_229),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_322),
.Y(n_347)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_241),
.B(n_237),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_244),
.B(n_180),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_325),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_246),
.A2(n_226),
.B1(n_209),
.B2(n_189),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_229),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_326),
.B(n_242),
.Y(n_355)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_239),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_236),
.A2(n_183),
.B1(n_201),
.B2(n_216),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g378 ( 
.A(n_333),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_334),
.A2(n_348),
.B1(n_361),
.B2(n_363),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_337),
.A2(n_356),
.B(n_296),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_340),
.A2(n_352),
.B(n_354),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_267),
.B1(n_235),
.B2(n_250),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_344),
.Y(n_371)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_261),
.C(n_250),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_307),
.C(n_316),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_311),
.A2(n_267),
.B1(n_270),
.B2(n_261),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_311),
.A2(n_270),
.B1(n_274),
.B2(n_207),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_369),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_323),
.A2(n_274),
.B1(n_222),
.B2(n_207),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_295),
.A2(n_243),
.B(n_280),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_297),
.A2(n_280),
.B(n_271),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_355),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_297),
.A2(n_275),
.B(n_253),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_308),
.A2(n_222),
.B1(n_273),
.B2(n_239),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_321),
.A2(n_325),
.B1(n_308),
.B2(n_324),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_362),
.A2(n_365),
.B(n_317),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_304),
.A2(n_219),
.B1(n_268),
.B2(n_273),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_308),
.A2(n_184),
.B(n_178),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_364),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_321),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_368),
.A2(n_286),
.B1(n_300),
.B2(n_17),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_291),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_293),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_370),
.B(n_302),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_374),
.B(n_379),
.Y(n_422)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_301),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_383),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_358),
.B(n_294),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_392),
.C(n_396),
.Y(n_421)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_331),
.B(n_301),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_353),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_384),
.B(n_385),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_355),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_387),
.A2(n_397),
.B1(n_347),
.B2(n_333),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_326),
.Y(n_388)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_388),
.Y(n_416)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_360),
.Y(n_389)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_390),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_404),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_302),
.C(n_287),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_355),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_393),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_347),
.B(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_338),
.B(n_343),
.C(n_335),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_399),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_284),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_329),
.B(n_362),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_402),
.Y(n_418)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_403),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_357),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_289),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_396),
.B(n_335),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_411),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_378),
.A2(n_334),
.B1(n_349),
.B2(n_337),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_410),
.A2(n_419),
.B1(n_427),
.B2(n_386),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_367),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g414 ( 
.A(n_379),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_417),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_377),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_378),
.A2(n_349),
.B1(n_352),
.B2(n_363),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_420),
.A2(n_384),
.B1(n_402),
.B2(n_382),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_329),
.C(n_339),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_430),
.C(n_431),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_382),
.A2(n_348),
.B1(n_356),
.B2(n_364),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_367),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_341),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_394),
.B(n_345),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_432),
.B(n_383),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_344),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g451 ( 
.A(n_434),
.B(n_405),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_386),
.A2(n_370),
.B1(n_369),
.B2(n_340),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_435),
.A2(n_375),
.B1(n_397),
.B2(n_395),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_346),
.C(n_357),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_436),
.B(n_426),
.C(n_421),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_437),
.B(n_440),
.Y(n_473)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_439),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_434),
.A2(n_375),
.B1(n_373),
.B2(n_385),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_416),
.Y(n_442)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_442),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_429),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_445),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_444),
.A2(n_364),
.B1(n_424),
.B2(n_408),
.Y(n_479)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_422),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_423),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_446),
.B(n_454),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_427),
.A2(n_391),
.B1(n_399),
.B2(n_371),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_452),
.B1(n_456),
.B2(n_415),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_453),
.C(n_459),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_450),
.A2(n_461),
.B(n_390),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_448),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_371),
.C(n_399),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_423),
.B(n_388),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_409),
.A2(n_393),
.B1(n_373),
.B2(n_398),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_455),
.B(n_458),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_419),
.A2(n_361),
.B1(n_395),
.B2(n_387),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_425),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_425),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_404),
.C(n_401),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_389),
.C(n_405),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_460),
.B(n_451),
.C(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_433),
.B(n_315),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_462),
.B(n_351),
.Y(n_463)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_464),
.A2(n_479),
.B1(n_437),
.B2(n_440),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_468),
.C(n_469),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_436),
.C(n_415),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_415),
.C(n_431),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_410),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_470),
.B(n_474),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_471),
.B(n_359),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_413),
.C(n_428),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_475),
.B(n_476),
.C(n_477),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_447),
.B(n_430),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_409),
.C(n_412),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_450),
.A2(n_424),
.B(n_390),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_481),
.B(n_336),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_453),
.B(n_408),
.C(n_424),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_336),
.C(n_330),
.Y(n_491)
);

AOI322xp5_ASAP7_75t_SL g485 ( 
.A1(n_484),
.A2(n_438),
.A3(n_443),
.B1(n_456),
.B2(n_444),
.C1(n_445),
.C2(n_368),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_485),
.B(n_305),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_488),
.B1(n_493),
.B2(n_474),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_480),
.A2(n_458),
.B1(n_457),
.B2(n_461),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_487),
.B(n_492),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_479),
.A2(n_455),
.B1(n_364),
.B2(n_365),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_476),
.C(n_468),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_359),
.Y(n_493)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_472),
.B(n_359),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_498),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_473),
.A2(n_354),
.B1(n_376),
.B2(n_374),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_497),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_482),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_467),
.B(n_477),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_500),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_366),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_502),
.B(n_489),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g521 ( 
.A(n_504),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_495),
.A2(n_483),
.B(n_465),
.Y(n_506)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_506),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_486),
.A2(n_478),
.B1(n_470),
.B2(n_469),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_508),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_493),
.A2(n_466),
.B(n_465),
.Y(n_508)
);

INVx11_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_487),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_490),
.B(n_350),
.C(n_320),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_489),
.C(n_490),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_499),
.A2(n_285),
.B(n_306),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g518 ( 
.A(n_512),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_496),
.Y(n_524)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_523),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_514),
.A2(n_491),
.B(n_488),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_520),
.B(n_507),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_524),
.A2(n_525),
.B1(n_509),
.B2(n_503),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_511),
.B(n_327),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_504),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_526),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_514),
.B(n_510),
.Y(n_527)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_527),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_531),
.C(n_518),
.Y(n_535)
);

AOI322xp5_ASAP7_75t_L g532 ( 
.A1(n_528),
.A2(n_521),
.A3(n_516),
.B1(n_520),
.B2(n_505),
.C1(n_510),
.C2(n_512),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_527),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_529),
.Y(n_536)
);

AOI322xp5_ASAP7_75t_L g538 ( 
.A1(n_536),
.A2(n_537),
.A3(n_534),
.B1(n_533),
.B2(n_526),
.C1(n_530),
.C2(n_519),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_508),
.C(n_502),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_539),
.A2(n_515),
.B(n_317),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_515),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_318),
.C(n_290),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_542),
.B(n_17),
.Y(n_543)
);


endmodule