module real_aes_15897_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
OAI22xp33_ASAP7_75t_SL g807 ( .A1(n_0), .A2(n_133), .B1(n_499), .B2(n_513), .Y(n_807) );
OAI22xp33_ASAP7_75t_L g818 ( .A1(n_0), .A2(n_25), .B1(n_398), .B2(n_399), .Y(n_818) );
INVx1_ASAP7_75t_L g591 ( .A(n_1), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_2), .A2(n_26), .B1(n_428), .B2(n_456), .Y(n_847) );
OAI22xp5_ASAP7_75t_SL g856 ( .A1(n_2), .A2(n_139), .B1(n_398), .B2(n_420), .Y(n_856) );
INVx1_ASAP7_75t_L g950 ( .A(n_3), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_4), .A2(n_264), .B1(n_476), .B2(n_480), .Y(n_475) );
INVxp33_ASAP7_75t_SL g543 ( .A(n_4), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_5), .Y(n_850) );
OAI211xp5_ASAP7_75t_L g1070 ( .A1(n_6), .A2(n_438), .B(n_615), .C(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1080 ( .A(n_6), .Y(n_1080) );
INVx1_ASAP7_75t_L g998 ( .A(n_7), .Y(n_998) );
INVx1_ASAP7_75t_L g934 ( .A(n_8), .Y(n_934) );
INVx1_ASAP7_75t_L g1373 ( .A(n_9), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_10), .Y(n_824) );
INVx1_ASAP7_75t_L g295 ( .A(n_11), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_11), .B(n_305), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_12), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_13), .A2(n_238), .B1(n_681), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_13), .A2(n_57), .B1(n_911), .B2(n_912), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_14), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g785 ( .A(n_15), .Y(n_785) );
INVx1_ASAP7_75t_L g1387 ( .A(n_16), .Y(n_1387) );
OAI222xp33_ASAP7_75t_L g870 ( .A1(n_17), .A2(n_220), .B1(n_429), .B2(n_449), .C1(n_871), .C2(n_873), .Y(n_870) );
OAI222xp33_ASAP7_75t_L g900 ( .A1(n_17), .A2(n_160), .B1(n_220), .B2(n_650), .C1(n_901), .C2(n_902), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_18), .A2(n_191), .B1(n_297), .B2(n_499), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_18), .A2(n_191), .B1(n_521), .B2(n_628), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_19), .A2(n_405), .B(n_714), .C(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g727 ( .A(n_19), .Y(n_727) );
INVx1_ASAP7_75t_L g1032 ( .A(n_20), .Y(n_1032) );
INVx1_ASAP7_75t_L g1085 ( .A(n_21), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_22), .B(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_22), .B(n_115), .Y(n_1167) );
INVx2_ASAP7_75t_L g1171 ( .A(n_22), .Y(n_1171) );
OAI22xp33_ASAP7_75t_SL g579 ( .A1(n_23), .A2(n_24), .B1(n_580), .B2(n_581), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_23), .A2(n_24), .B1(n_536), .B2(n_635), .Y(n_634) );
OAI22xp33_ASAP7_75t_SL g804 ( .A1(n_25), .A2(n_248), .B1(n_428), .B2(n_805), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_26), .B(n_419), .Y(n_855) );
OAI22xp33_ASAP7_75t_L g951 ( .A1(n_27), .A2(n_226), .B1(n_398), .B2(n_952), .Y(n_951) );
OAI22xp33_ASAP7_75t_L g962 ( .A1(n_27), .A2(n_273), .B1(n_428), .B2(n_430), .Y(n_962) );
INVx1_ASAP7_75t_L g736 ( .A(n_28), .Y(n_736) );
INVx1_ASAP7_75t_L g606 ( .A(n_29), .Y(n_606) );
INVx1_ASAP7_75t_L g995 ( .A(n_30), .Y(n_995) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_31), .A2(n_196), .B1(n_1172), .B2(n_1177), .Y(n_1176) );
INVx1_ASAP7_75t_L g885 ( .A(n_32), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_32), .A2(n_238), .B1(n_912), .B2(n_920), .Y(n_919) );
XOR2xp5_ASAP7_75t_L g774 ( .A(n_33), .B(n_775), .Y(n_774) );
AOI22xp5_ASAP7_75t_L g1208 ( .A1(n_34), .A2(n_183), .B1(n_1166), .B2(n_1172), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1466 ( .A1(n_35), .A2(n_218), .B1(n_1142), .B2(n_1463), .Y(n_1466) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_35), .A2(n_242), .B1(n_489), .B2(n_1028), .Y(n_1474) );
XNOR2x2_ASAP7_75t_SL g709 ( .A(n_36), .B(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_36), .A2(n_210), .B1(n_1162), .B2(n_1169), .Y(n_1257) );
OAI22xp33_ASAP7_75t_L g975 ( .A1(n_37), .A2(n_151), .B1(n_428), .B2(n_430), .Y(n_975) );
OAI22xp33_ASAP7_75t_SL g977 ( .A1(n_37), .A2(n_151), .B1(n_398), .B2(n_978), .Y(n_977) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_38), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_39), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_40), .Y(n_788) );
INVx1_ASAP7_75t_L g719 ( .A(n_41), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g724 ( .A1(n_41), .A2(n_383), .B(n_725), .C(n_726), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_42), .A2(n_122), .B1(n_488), .B2(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g559 ( .A(n_42), .Y(n_559) );
INVx1_ASAP7_75t_L g644 ( .A(n_43), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_44), .A2(n_119), .B1(n_1162), .B2(n_1169), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g1069 ( .A1(n_45), .A2(n_137), .B1(n_455), .B2(n_456), .Y(n_1069) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_45), .A2(n_62), .B1(n_399), .B2(n_420), .Y(n_1081) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_46), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_47), .A2(n_215), .B1(n_1162), .B2(n_1172), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_48), .A2(n_188), .B1(n_399), .B2(n_420), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_48), .A2(n_49), .B1(n_455), .B2(n_456), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_49), .A2(n_278), .B1(n_398), .B2(n_419), .Y(n_1024) );
AOI22xp5_ASAP7_75t_L g1207 ( .A1(n_50), .A2(n_108), .B1(n_1162), .B2(n_1169), .Y(n_1207) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_51), .A2(n_162), .B1(n_650), .B2(n_651), .Y(n_649) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_51), .Y(n_661) );
INVx1_ASAP7_75t_L g973 ( .A(n_52), .Y(n_973) );
INVx1_ASAP7_75t_L g1409 ( .A(n_53), .Y(n_1409) );
INVx1_ASAP7_75t_L g321 ( .A(n_54), .Y(n_321) );
INVx1_ASAP7_75t_L g329 ( .A(n_54), .Y(n_329) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_55), .A2(n_90), .B1(n_1463), .B2(n_1465), .Y(n_1462) );
AOI22xp33_ASAP7_75t_SL g1475 ( .A1(n_55), .A2(n_99), .B1(n_470), .B2(n_693), .Y(n_1475) );
INVx1_ASAP7_75t_L g1448 ( .A(n_56), .Y(n_1448) );
OAI221xp5_ASAP7_75t_L g1455 ( .A1(n_56), .A2(n_113), .B1(n_353), .B2(n_651), .C(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g886 ( .A(n_57), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g825 ( .A(n_58), .Y(n_825) );
XOR2x2_ASAP7_75t_L g640 ( .A(n_59), .B(n_641), .Y(n_640) );
XOR2xp5_ASAP7_75t_L g921 ( .A(n_60), .B(n_922), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_61), .A2(n_82), .B1(n_679), .B2(n_681), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_61), .A2(n_252), .B1(n_699), .B2(n_705), .Y(n_704) );
OAI22xp33_ASAP7_75t_L g1074 ( .A1(n_62), .A2(n_213), .B1(n_428), .B2(n_430), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_63), .A2(n_209), .B1(n_1122), .B2(n_1129), .Y(n_1128) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_63), .A2(n_214), .B1(n_1138), .B2(n_1142), .Y(n_1143) );
INVx1_ASAP7_75t_L g288 ( .A(n_64), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g511 ( .A1(n_65), .A2(n_230), .B1(n_512), .B2(n_514), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g533 ( .A1(n_65), .A2(n_230), .B1(n_534), .B2(n_536), .Y(n_533) );
INVx2_ASAP7_75t_L g349 ( .A(n_66), .Y(n_349) );
INVx1_ASAP7_75t_L g607 ( .A(n_67), .Y(n_607) );
INVx1_ASAP7_75t_L g927 ( .A(n_68), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_69), .A2(n_253), .B1(n_920), .B2(n_1010), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_69), .A2(n_190), .B1(n_688), .B2(n_1056), .Y(n_1057) );
INVxp67_ASAP7_75t_SL g647 ( .A(n_70), .Y(n_647) );
OAI22xp33_ASAP7_75t_L g662 ( .A1(n_70), .A2(n_162), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_71), .A2(n_95), .B1(n_1169), .B2(n_1177), .Y(n_1190) );
INVx1_ASAP7_75t_L g1031 ( .A(n_72), .Y(n_1031) );
INVx1_ASAP7_75t_L g1073 ( .A(n_73), .Y(n_1073) );
INVx1_ASAP7_75t_L g1027 ( .A(n_74), .Y(n_1027) );
OAI22xp33_ASAP7_75t_L g418 ( .A1(n_75), .A2(n_269), .B1(n_419), .B2(n_420), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_75), .A2(n_269), .B1(n_455), .B2(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g746 ( .A(n_76), .Y(n_746) );
INVx1_ASAP7_75t_L g485 ( .A(n_77), .Y(n_485) );
OAI22xp33_ASAP7_75t_SL g397 ( .A1(n_78), .A2(n_275), .B1(n_398), .B2(n_399), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g427 ( .A1(n_78), .A2(n_275), .B1(n_428), .B2(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g1088 ( .A(n_79), .Y(n_1088) );
OAI222xp33_ASAP7_75t_L g1115 ( .A1(n_80), .A2(n_117), .B1(n_246), .B2(n_592), .C1(n_811), .C2(n_1116), .Y(n_1115) );
OAI222xp33_ASAP7_75t_L g1150 ( .A1(n_80), .A2(n_117), .B1(n_246), .B2(n_615), .C1(n_663), .C2(n_664), .Y(n_1150) );
INVx1_ASAP7_75t_L g1371 ( .A(n_81), .Y(n_1371) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_82), .A2(n_96), .B1(n_489), .B2(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g991 ( .A(n_83), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_84), .A2(n_279), .B1(n_1125), .B2(n_1127), .Y(n_1124) );
AOI22xp33_ASAP7_75t_SL g1144 ( .A1(n_84), .A2(n_147), .B1(n_1061), .B2(n_1145), .Y(n_1144) );
XOR2xp5_ASAP7_75t_L g862 ( .A(n_85), .B(n_863), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g1196 ( .A1(n_85), .A2(n_140), .B1(n_1162), .B2(n_1169), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_86), .A2(n_147), .B1(n_1013), .B2(n_1131), .Y(n_1130) );
AOI22xp33_ASAP7_75t_SL g1137 ( .A1(n_86), .A2(n_279), .B1(n_1138), .B2(n_1142), .Y(n_1137) );
INVx1_ASAP7_75t_L g331 ( .A(n_87), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g1011 ( .A1(n_88), .A2(n_277), .B1(n_1012), .B2(n_1013), .C(n_1015), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_88), .A2(n_145), .B1(n_1059), .B2(n_1061), .Y(n_1058) );
INVx1_ASAP7_75t_L g509 ( .A(n_89), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_90), .A2(n_203), .B1(n_693), .B2(n_1472), .Y(n_1471) );
INVx1_ASAP7_75t_L g972 ( .A(n_91), .Y(n_972) );
INVx1_ASAP7_75t_L g1375 ( .A(n_92), .Y(n_1375) );
INVx1_ASAP7_75t_L g316 ( .A(n_93), .Y(n_316) );
INVx1_ASAP7_75t_L g802 ( .A(n_94), .Y(n_802) );
OAI211xp5_ASAP7_75t_SL g810 ( .A1(n_94), .A2(n_526), .B(n_811), .C(n_812), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_96), .A2(n_252), .B1(n_677), .B2(n_688), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_97), .A2(n_100), .B1(n_536), .B2(n_628), .Y(n_1405) );
OAI22xp33_ASAP7_75t_L g1415 ( .A1(n_97), .A2(n_120), .B1(n_297), .B2(n_499), .Y(n_1415) );
XOR2x2_ASAP7_75t_L g966 ( .A(n_98), .B(n_967), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g1467 ( .A1(n_99), .A2(n_203), .B1(n_1468), .B2(n_1469), .Y(n_1467) );
OAI22xp5_ASAP7_75t_L g1416 ( .A1(n_100), .A2(n_184), .B1(n_1417), .B2(n_1419), .Y(n_1416) );
AOI22xp5_ASAP7_75t_L g1187 ( .A1(n_101), .A2(n_138), .B1(n_1162), .B2(n_1169), .Y(n_1187) );
OAI221xp5_ASAP7_75t_L g946 ( .A1(n_102), .A2(n_273), .B1(n_399), .B2(n_419), .C(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g960 ( .A(n_102), .Y(n_960) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_103), .A2(n_180), .B1(n_455), .B2(n_456), .Y(n_974) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_103), .A2(n_180), .B1(n_419), .B2(n_420), .Y(n_984) );
AOI22xp5_ASAP7_75t_SL g1186 ( .A1(n_104), .A2(n_265), .B1(n_1172), .B2(n_1177), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1451 ( .A1(n_105), .A2(n_221), .B1(n_455), .B2(n_456), .Y(n_1451) );
OAI22xp5_ASAP7_75t_L g1457 ( .A1(n_105), .A2(n_221), .B1(n_419), .B2(n_420), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_106), .Y(n_290) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_106), .B(n_288), .Y(n_1163) );
OAI211xp5_ASAP7_75t_L g865 ( .A1(n_107), .A2(n_866), .B(n_867), .C(n_877), .Y(n_865) );
INVx1_ASAP7_75t_L g906 ( .A(n_107), .Y(n_906) );
INVx1_ASAP7_75t_L g745 ( .A(n_109), .Y(n_745) );
INVx1_ASAP7_75t_L g929 ( .A(n_110), .Y(n_929) );
INVx1_ASAP7_75t_L g577 ( .A(n_111), .Y(n_577) );
INVx1_ASAP7_75t_L g1388 ( .A(n_112), .Y(n_1388) );
INVx1_ASAP7_75t_L g1450 ( .A(n_113), .Y(n_1450) );
AOI22xp33_ASAP7_75t_SL g1181 ( .A1(n_114), .A2(n_123), .B1(n_1166), .B2(n_1172), .Y(n_1181) );
INVx1_ASAP7_75t_L g1165 ( .A(n_115), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_115), .B(n_1171), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_116), .A2(n_272), .B1(n_1162), .B2(n_1166), .Y(n_1161) );
INVx1_ASAP7_75t_L g930 ( .A(n_118), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_120), .A2(n_184), .B1(n_1412), .B2(n_1413), .Y(n_1411) );
INVx1_ASAP7_75t_L g653 ( .A(n_121), .Y(n_653) );
INVx1_ASAP7_75t_L g545 ( .A(n_122), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_124), .A2(n_236), .B1(n_952), .B2(n_1114), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1149 ( .A1(n_124), .A2(n_236), .B1(n_580), .B2(n_805), .Y(n_1149) );
INVx2_ASAP7_75t_L g348 ( .A(n_125), .Y(n_348) );
INVx1_ASAP7_75t_L g358 ( .A(n_125), .Y(n_358) );
INVx1_ASAP7_75t_L g740 ( .A(n_126), .Y(n_740) );
INVx1_ASAP7_75t_L g1092 ( .A(n_127), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_128), .A2(n_263), .B1(n_679), .B2(n_681), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_128), .A2(n_197), .B1(n_484), .B2(n_693), .Y(n_701) );
INVx1_ASAP7_75t_L g362 ( .A(n_129), .Y(n_362) );
INVx1_ASAP7_75t_L g989 ( .A(n_130), .Y(n_989) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_131), .A2(n_244), .B1(n_1162), .B2(n_1169), .Y(n_1178) );
XNOR2xp5_ASAP7_75t_L g567 ( .A(n_132), .B(n_568), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_133), .A2(n_248), .B1(n_419), .B2(n_420), .Y(n_809) );
OAI22xp33_ASAP7_75t_SL g853 ( .A1(n_134), .A2(n_139), .B1(n_430), .B2(n_455), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_134), .A2(n_143), .B1(n_815), .B2(n_816), .Y(n_860) );
INVx1_ASAP7_75t_L g1110 ( .A(n_135), .Y(n_1110) );
XOR2xp5_ASAP7_75t_L g1436 ( .A(n_136), .B(n_1437), .Y(n_1436) );
OAI22xp5_ASAP7_75t_SL g1076 ( .A1(n_137), .A2(n_213), .B1(n_398), .B2(n_419), .Y(n_1076) );
INVx1_ASAP7_75t_L g1095 ( .A(n_141), .Y(n_1095) );
INVx1_ASAP7_75t_L g997 ( .A(n_142), .Y(n_997) );
INVx1_ASAP7_75t_L g851 ( .A(n_143), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_144), .A2(n_243), .B1(n_398), .B2(n_721), .Y(n_720) );
OAI22xp33_ASAP7_75t_L g731 ( .A1(n_144), .A2(n_243), .B1(n_428), .B2(n_499), .Y(n_731) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_145), .A2(n_228), .B1(n_1012), .B2(n_1013), .C(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g352 ( .A(n_146), .Y(n_352) );
XOR2xp5_ASAP7_75t_L g1106 ( .A(n_148), .B(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g472 ( .A(n_149), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g1194 ( .A1(n_150), .A2(n_256), .B1(n_1172), .B2(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1381 ( .A(n_152), .Y(n_1381) );
INVx1_ASAP7_75t_L g756 ( .A(n_153), .Y(n_756) );
INVx1_ASAP7_75t_L g876 ( .A(n_154), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_154), .A2(n_233), .B1(n_419), .B2(n_420), .Y(n_903) );
INVx1_ASAP7_75t_L g1093 ( .A(n_155), .Y(n_1093) );
AOI31xp33_ASAP7_75t_L g1007 ( .A1(n_156), .A2(n_1008), .A3(n_1023), .B(n_1034), .Y(n_1007) );
NAND2xp33_ASAP7_75t_SL g1051 ( .A(n_156), .B(n_1052), .Y(n_1051) );
INVxp67_ASAP7_75t_SL g1064 ( .A(n_156), .Y(n_1064) );
INVx1_ASAP7_75t_L g1442 ( .A(n_157), .Y(n_1442) );
INVx1_ASAP7_75t_L g417 ( .A(n_158), .Y(n_417) );
OAI211xp5_ASAP7_75t_L g436 ( .A1(n_158), .A2(n_437), .B(n_438), .C(n_444), .Y(n_436) );
INVx1_ASAP7_75t_L g598 ( .A(n_159), .Y(n_598) );
INVx1_ASAP7_75t_L g868 ( .A(n_160), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g888 ( .A(n_161), .Y(n_888) );
BUFx3_ASAP7_75t_L g323 ( .A(n_163), .Y(n_323) );
OAI211xp5_ASAP7_75t_SL g848 ( .A1(n_164), .A2(n_438), .B(n_558), .C(n_849), .Y(n_848) );
OAI211xp5_ASAP7_75t_SL g857 ( .A1(n_164), .A2(n_526), .B(n_858), .C(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g324 ( .A(n_165), .Y(n_324) );
INVx1_ASAP7_75t_L g335 ( .A(n_166), .Y(n_335) );
INVx1_ASAP7_75t_L g1086 ( .A(n_167), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_168), .A2(n_257), .B1(n_297), .B2(n_499), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_168), .A2(n_257), .B1(n_519), .B2(n_521), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_169), .Y(n_414) );
XNOR2x1_ASAP7_75t_L g311 ( .A(n_170), .B(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_171), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_172), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_173), .Y(n_882) );
INVx1_ASAP7_75t_L g486 ( .A(n_174), .Y(n_486) );
INVx1_ASAP7_75t_L g602 ( .A(n_175), .Y(n_602) );
INVx1_ASAP7_75t_L g949 ( .A(n_176), .Y(n_949) );
XOR2x2_ASAP7_75t_L g1066 ( .A(n_177), .B(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_178), .A2(n_214), .B1(n_1028), .B2(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_178), .A2(n_209), .B1(n_679), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g510 ( .A(n_179), .Y(n_510) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_179), .A2(n_524), .B(n_526), .C(n_527), .Y(n_523) );
INVx1_ASAP7_75t_L g751 ( .A(n_181), .Y(n_751) );
INVx1_ASAP7_75t_L g1021 ( .A(n_182), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g1053 ( .A1(n_182), .A2(n_253), .B1(n_681), .B2(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g757 ( .A(n_185), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g1406 ( .A1(n_186), .A2(n_405), .B(n_1407), .C(n_1408), .Y(n_1406) );
INVx1_ASAP7_75t_L g1423 ( .A(n_186), .Y(n_1423) );
CKINVDCx5p33_ASAP7_75t_R g783 ( .A(n_187), .Y(n_783) );
INVxp67_ASAP7_75t_SL g1038 ( .A(n_188), .Y(n_1038) );
INVx1_ASAP7_75t_L g937 ( .A(n_189), .Y(n_937) );
INVx1_ASAP7_75t_L g1019 ( .A(n_190), .Y(n_1019) );
INVx1_ASAP7_75t_L g587 ( .A(n_192), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_193), .A2(n_207), .B1(n_419), .B2(n_635), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_193), .A2(n_207), .B1(n_513), .B2(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g881 ( .A(n_194), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_194), .B(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g645 ( .A(n_195), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_197), .A2(n_205), .B1(n_674), .B2(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g1096 ( .A(n_198), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_199), .B(n_412), .Y(n_948) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_199), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g1256 ( .A1(n_200), .A2(n_201), .B1(n_1166), .B2(n_1172), .Y(n_1256) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_202), .Y(n_791) );
OAI211xp5_ASAP7_75t_L g800 ( .A1(n_204), .A2(n_438), .B(n_558), .C(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g817 ( .A(n_204), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_205), .A2(n_263), .B1(n_484), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g1378 ( .A(n_206), .Y(n_1378) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_208), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_211), .Y(n_780) );
INVx1_ASAP7_75t_L g1072 ( .A(n_212), .Y(n_1072) );
INVx1_ASAP7_75t_L g1384 ( .A(n_216), .Y(n_1384) );
INVx1_ASAP7_75t_L g754 ( .A(n_217), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g1476 ( .A1(n_218), .A2(n_267), .B1(n_489), .B2(n_699), .C(n_1015), .Y(n_1476) );
INVx1_ASAP7_75t_L g933 ( .A(n_219), .Y(n_933) );
OAI211xp5_ASAP7_75t_L g500 ( .A1(n_222), .A2(n_501), .B(n_505), .C(n_508), .Y(n_500) );
INVx1_ASAP7_75t_L g532 ( .A(n_222), .Y(n_532) );
INVx1_ASAP7_75t_L g994 ( .A(n_223), .Y(n_994) );
INVx1_ASAP7_75t_L g351 ( .A(n_224), .Y(n_351) );
INVx1_ASAP7_75t_L g1090 ( .A(n_225), .Y(n_1090) );
INVxp67_ASAP7_75t_SL g959 ( .A(n_226), .Y(n_959) );
INVx1_ASAP7_75t_L g578 ( .A(n_227), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g630 ( .A1(n_227), .A2(n_526), .B(n_631), .C(n_632), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_228), .A2(n_277), .B1(n_688), .B2(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1443 ( .A(n_229), .Y(n_1443) );
XOR2xp5_ASAP7_75t_L g819 ( .A(n_231), .B(n_820), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_232), .Y(n_835) );
INVx1_ASAP7_75t_L g878 ( .A(n_233), .Y(n_878) );
INVx1_ASAP7_75t_L g992 ( .A(n_234), .Y(n_992) );
BUFx3_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
INVx1_ASAP7_75t_L g433 ( .A(n_235), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_237), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_239), .Y(n_827) );
INVx1_ASAP7_75t_L g926 ( .A(n_240), .Y(n_926) );
INVx1_ASAP7_75t_L g1410 ( .A(n_241), .Y(n_1410) );
OAI211xp5_ASAP7_75t_L g1421 ( .A1(n_241), .A2(n_572), .B(n_573), .C(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_242), .A2(n_267), .B1(n_1061), .B2(n_1145), .Y(n_1461) );
INVx1_ASAP7_75t_L g988 ( .A(n_245), .Y(n_988) );
INVx1_ASAP7_75t_L g366 ( .A(n_247), .Y(n_366) );
INVx1_ASAP7_75t_L g346 ( .A(n_249), .Y(n_346) );
INVx2_ASAP7_75t_L g356 ( .A(n_249), .Y(n_356) );
INVx1_ASAP7_75t_L g496 ( .A(n_249), .Y(n_496) );
INVx1_ASAP7_75t_L g717 ( .A(n_250), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g969 ( .A1(n_251), .A2(n_438), .B(n_970), .C(n_971), .Y(n_969) );
INVx1_ASAP7_75t_L g981 ( .A(n_251), .Y(n_981) );
XNOR2x1_ASAP7_75t_L g464 ( .A(n_254), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g1168 ( .A1(n_255), .A2(n_259), .B1(n_1169), .B2(n_1172), .Y(n_1168) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_258), .Y(n_787) );
INVx1_ASAP7_75t_L g594 ( .A(n_260), .Y(n_594) );
INVx1_ASAP7_75t_L g936 ( .A(n_261), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g1447 ( .A(n_262), .Y(n_1447) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_264), .Y(n_557) );
INVx1_ASAP7_75t_L g654 ( .A(n_266), .Y(n_654) );
INVx1_ASAP7_75t_L g474 ( .A(n_268), .Y(n_474) );
AOI21xp33_ASAP7_75t_L g890 ( .A1(n_270), .A2(n_688), .B(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g909 ( .A(n_270), .Y(n_909) );
INVx1_ASAP7_75t_L g1111 ( .A(n_271), .Y(n_1111) );
XOR2x2_ASAP7_75t_L g1366 ( .A(n_272), .B(n_1367), .Y(n_1366) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_272), .A2(n_1430), .B1(n_1435), .B2(n_1477), .Y(n_1429) );
OAI211xp5_ASAP7_75t_L g571 ( .A1(n_274), .A2(n_572), .B(n_573), .C(n_574), .Y(n_571) );
INVx1_ASAP7_75t_L g633 ( .A(n_274), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g874 ( .A(n_276), .Y(n_874) );
INVx1_ASAP7_75t_L g1036 ( .A(n_278), .Y(n_1036) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_280), .A2(n_404), .B(n_405), .C(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g453 ( .A(n_280), .Y(n_453) );
INVx1_ASAP7_75t_L g596 ( .A(n_281), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_306), .B(n_1154), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_291), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g1428 ( .A(n_285), .B(n_294), .Y(n_1428) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1434 ( .A(n_287), .B(n_290), .Y(n_1434) );
INVx1_ASAP7_75t_L g1480 ( .A(n_287), .Y(n_1480) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_290), .B(n_1480), .Y(n_1482) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g458 ( .A(n_294), .B(n_459), .Y(n_458) );
AOI21xp5_ASAP7_75t_SL g864 ( .A1(n_294), .A2(n_865), .B(n_879), .Y(n_864) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g393 ( .A(n_295), .B(n_305), .Y(n_393) );
AND2x4_ASAP7_75t_L g892 ( .A(n_295), .B(n_304), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_296), .A2(n_431), .B1(n_1110), .B2(n_1111), .Y(n_1147) );
AND2x4_ASAP7_75t_SL g1427 ( .A(n_296), .B(n_1428), .Y(n_1427) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
OR2x2_ASAP7_75t_L g455 ( .A(n_298), .B(n_432), .Y(n_455) );
OR2x6_ASAP7_75t_L g513 ( .A(n_298), .B(n_432), .Y(n_513) );
BUFx4f_ASAP7_75t_L g544 ( .A(n_298), .Y(n_544) );
INVx1_ASAP7_75t_L g798 ( .A(n_298), .Y(n_798) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx4f_ASAP7_75t_L g373 ( .A(n_299), .Y(n_373) );
INVx3_ASAP7_75t_L g429 ( .A(n_299), .Y(n_429) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g378 ( .A(n_301), .Y(n_378) );
INVx2_ASAP7_75t_L g382 ( .A(n_301), .Y(n_382) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_301), .B(n_302), .Y(n_385) );
AND2x2_ASAP7_75t_L g434 ( .A(n_301), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g443 ( .A(n_301), .B(n_302), .Y(n_443) );
INVx1_ASAP7_75t_L g452 ( .A(n_301), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_302), .B(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g381 ( .A(n_302), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g435 ( .A(n_302), .Y(n_435) );
BUFx2_ASAP7_75t_L g447 ( .A(n_302), .Y(n_447) );
INVx1_ASAP7_75t_L g669 ( .A(n_302), .Y(n_669) );
AND2x2_ASAP7_75t_L g682 ( .A(n_302), .B(n_378), .Y(n_682) );
OR2x6_ASAP7_75t_L g428 ( .A(n_303), .B(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_303), .A2(n_874), .B1(n_875), .B2(n_876), .Y(n_873) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g440 ( .A(n_304), .Y(n_440) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g446 ( .A(n_305), .Y(n_446) );
AND2x4_ASAP7_75t_L g450 ( .A(n_305), .B(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B1(n_769), .B2(n_770), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
XOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_638), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_461), .B1(n_462), .B2(n_637), .Y(n_309) );
INVx1_ASAP7_75t_L g637 ( .A(n_310), .Y(n_637) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND3x1_ASAP7_75t_L g312 ( .A(n_313), .B(n_396), .C(n_426), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_367), .Y(n_313) );
OAI33xp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_330), .A3(n_342), .B1(n_350), .B2(n_354), .B3(n_360), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_324), .B2(n_325), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_316), .A2(n_362), .B1(n_380), .B2(n_383), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_317), .A2(n_752), .B1(n_787), .B2(n_788), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_317), .A2(n_829), .B1(n_1088), .B2(n_1095), .Y(n_1100) );
INVx2_ASAP7_75t_L g1377 ( .A(n_317), .Y(n_1377) );
INVx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_SL g361 ( .A(n_318), .Y(n_361) );
INVx5_ASAP7_75t_L g601 ( .A(n_318), .Y(n_601) );
INVx2_ASAP7_75t_SL g1473 ( .A(n_318), .Y(n_1473) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_319), .Y(n_402) );
INVx2_ASAP7_75t_L g471 ( .A(n_319), .Y(n_471) );
BUFx8_ASAP7_75t_L g750 ( .A(n_319), .Y(n_750) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g334 ( .A(n_321), .Y(n_334) );
AND2x4_ASAP7_75t_L g478 ( .A(n_322), .B(n_479), .Y(n_478) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_323), .B(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g333 ( .A(n_323), .B(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_323), .Y(n_341) );
AND2x4_ASAP7_75t_L g407 ( .A(n_323), .B(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_324), .A2(n_366), .B1(n_372), .B2(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_325), .A2(n_361), .B1(n_831), .B2(n_832), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_325), .A2(n_595), .B1(n_1090), .B2(n_1096), .Y(n_1101) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g747 ( .A(n_326), .Y(n_747) );
INVx3_ASAP7_75t_L g829 ( .A(n_326), .Y(n_829) );
CKINVDCx8_ASAP7_75t_R g918 ( .A(n_326), .Y(n_918) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g753 ( .A(n_327), .Y(n_753) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g365 ( .A(n_328), .Y(n_365) );
INVx1_ASAP7_75t_L g340 ( .A(n_329), .Y(n_340) );
INVx2_ASAP7_75t_L g408 ( .A(n_329), .Y(n_408) );
OAI22xp5_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_332), .B1(n_335), .B2(n_336), .Y(n_330) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_331), .A2(n_351), .B1(n_372), .B2(n_374), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_332), .A2(n_351), .B1(n_352), .B2(n_353), .Y(n_350) );
OAI22xp33_ASAP7_75t_L g778 ( .A1(n_332), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
OAI22xp33_ASAP7_75t_L g789 ( .A1(n_332), .A2(n_353), .B1(n_790), .B2(n_791), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_332), .A2(n_336), .B1(n_824), .B2(n_825), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_332), .A2(n_353), .B1(n_834), .B2(n_835), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_332), .A2(n_901), .B1(n_926), .B2(n_927), .Y(n_925) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_332), .A2(n_781), .B1(n_936), .B2(n_937), .Y(n_935) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_332), .A2(n_781), .B1(n_988), .B2(n_989), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_332), .A2(n_353), .B1(n_997), .B2(n_998), .Y(n_996) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_332), .A2(n_1086), .B1(n_1093), .B2(n_1103), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_332), .Y(n_1372) );
HB1xp67_ASAP7_75t_L g1386 ( .A(n_332), .Y(n_1386) );
BUFx4f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x4_ASAP7_75t_L g398 ( .A(n_333), .B(n_359), .Y(n_398) );
OR2x4_ASAP7_75t_L g419 ( .A(n_333), .B(n_401), .Y(n_419) );
BUFx3_ASAP7_75t_L g590 ( .A(n_333), .Y(n_590) );
BUFx3_ASAP7_75t_L g605 ( .A(n_333), .Y(n_605) );
INVx2_ASAP7_75t_L g739 ( .A(n_333), .Y(n_739) );
INVx1_ASAP7_75t_L g479 ( .A(n_334), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_335), .A2(n_352), .B1(n_387), .B2(n_389), .Y(n_386) );
INVx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g1407 ( .A(n_337), .Y(n_1407) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx4_ASAP7_75t_L g525 ( .A(n_338), .Y(n_525) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_338), .Y(n_781) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g353 ( .A(n_339), .Y(n_353) );
BUFx2_ASAP7_75t_L g743 ( .A(n_339), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
BUFx2_ASAP7_75t_L g416 ( .A(n_340), .Y(n_416) );
BUFx2_ASAP7_75t_L g413 ( .A(n_341), .Y(n_413) );
AND2x4_ASAP7_75t_L g694 ( .A(n_341), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g816 ( .A(n_341), .Y(n_816) );
BUFx3_ASAP7_75t_L g481 ( .A(n_342), .Y(n_481) );
OAI33xp33_ASAP7_75t_L g585 ( .A1(n_342), .A2(n_586), .A3(n_593), .B1(n_597), .B2(n_603), .B3(n_604), .Y(n_585) );
OAI33xp33_ASAP7_75t_L g777 ( .A1(n_342), .A2(n_354), .A3(n_778), .B1(n_782), .B2(n_786), .B3(n_789), .Y(n_777) );
OAI33xp33_ASAP7_75t_L g822 ( .A1(n_342), .A2(n_354), .A3(n_823), .B1(n_826), .B2(n_830), .B3(n_833), .Y(n_822) );
OAI33xp33_ASAP7_75t_L g986 ( .A1(n_342), .A2(n_354), .A3(n_987), .B1(n_990), .B2(n_993), .B3(n_996), .Y(n_986) );
OAI33xp33_ASAP7_75t_L g1097 ( .A1(n_342), .A2(n_354), .A3(n_1098), .B1(n_1100), .B2(n_1101), .B3(n_1102), .Y(n_1097) );
BUFx4f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx2_ASAP7_75t_L g734 ( .A(n_343), .Y(n_734) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_347), .Y(n_343) );
AND2x2_ASAP7_75t_SL g392 ( .A(n_344), .B(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_344), .Y(n_425) );
INVx1_ASAP7_75t_L g566 ( .A(n_344), .Y(n_566) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g460 ( .A(n_345), .Y(n_460) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_349), .Y(n_347) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_348), .Y(n_423) );
AND3x4_ASAP7_75t_L g696 ( .A(n_348), .B(n_412), .C(n_697), .Y(n_696) );
INVx3_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
BUFx3_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
INVx2_ASAP7_75t_L g715 ( .A(n_353), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_353), .A2(n_738), .B1(n_756), .B2(n_757), .Y(n_755) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_353), .A2(n_1085), .B1(n_1092), .B2(n_1099), .Y(n_1098) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
AND2x4_ASAP7_75t_L g369 ( .A(n_355), .B(n_370), .Y(n_369) );
OR2x6_ASAP7_75t_L g758 ( .A(n_355), .B(n_357), .Y(n_758) );
INVx1_ASAP7_75t_L g896 ( .A(n_355), .Y(n_896) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g697 ( .A(n_356), .Y(n_697) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND3x1_ASAP7_75t_L g494 ( .A(n_358), .B(n_359), .C(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g401 ( .A(n_359), .Y(n_401) );
AND2x4_ASAP7_75t_L g406 ( .A(n_359), .B(n_407), .Y(n_406) );
OR2x6_ASAP7_75t_L g420 ( .A(n_359), .B(n_365), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_363), .B2(n_366), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_363), .A2(n_783), .B1(n_784), .B2(n_785), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g990 ( .A1(n_363), .A2(n_932), .B1(n_991), .B2(n_992), .Y(n_990) );
OAI22xp33_ASAP7_75t_SL g1374 ( .A1(n_363), .A2(n_1375), .B1(n_1376), .B2(n_1378), .Y(n_1374) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g473 ( .A(n_365), .Y(n_473) );
OAI33xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .A3(n_379), .B1(n_386), .B2(n_391), .B3(n_394), .Y(n_367) );
OAI33xp33_ASAP7_75t_L g792 ( .A1(n_368), .A2(n_391), .A3(n_793), .B1(n_794), .B2(n_795), .B3(n_796), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g938 ( .A1(n_368), .A2(n_391), .A3(n_939), .B1(n_940), .B2(n_941), .B3(n_943), .Y(n_938) );
OAI33xp33_ASAP7_75t_L g999 ( .A1(n_368), .A2(n_391), .A3(n_1000), .B1(n_1001), .B2(n_1002), .B3(n_1003), .Y(n_999) );
OAI33xp33_ASAP7_75t_L g1389 ( .A1(n_368), .A2(n_625), .A3(n_1390), .B1(n_1394), .B2(n_1396), .B3(n_1399), .Y(n_1389) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g541 ( .A(n_369), .Y(n_541) );
INVx4_ASAP7_75t_L g685 ( .A(n_369), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_372), .A2(n_395), .B1(n_779), .B2(n_790), .Y(n_793) );
OAI22xp33_ASAP7_75t_L g1000 ( .A1(n_372), .A2(n_613), .B1(n_988), .B2(n_997), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_372), .A2(n_839), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_372), .A2(n_767), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx3_ASAP7_75t_L g612 ( .A(n_373), .Y(n_612) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_373), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_374), .Y(n_624) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx4_ASAP7_75t_L g395 ( .A(n_375), .Y(n_395) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_375), .Y(n_547) );
INVx1_ASAP7_75t_L g613 ( .A(n_375), .Y(n_613) );
INVx2_ASAP7_75t_SL g767 ( .A(n_375), .Y(n_767) );
INVx2_ASAP7_75t_L g840 ( .A(n_375), .Y(n_840) );
INVx8_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g456 ( .A(n_376), .B(n_440), .Y(n_456) );
OR2x2_ASAP7_75t_L g516 ( .A(n_376), .B(n_446), .Y(n_516) );
BUFx2_ASAP7_75t_L g763 ( .A(n_376), .Y(n_763) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_380), .A2(n_503), .B1(n_745), .B2(n_751), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_380), .A2(n_503), .B1(n_740), .B2(n_757), .Y(n_765) );
BUFx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g388 ( .A(n_381), .Y(n_388) );
BUFx2_ASAP7_75t_L g551 ( .A(n_381), .Y(n_551) );
INVx2_ASAP7_75t_L g556 ( .A(n_381), .Y(n_556) );
BUFx3_ASAP7_75t_L g843 ( .A(n_381), .Y(n_843) );
AND2x2_ASAP7_75t_L g668 ( .A(n_382), .B(n_669), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_383), .A2(n_387), .B1(n_827), .B2(n_831), .Y(n_841) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_383), .A2(n_1089), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1394 ( .A1(n_383), .A2(n_1375), .B1(n_1381), .B2(n_1395), .Y(n_1394) );
BUFx4f_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx4_ASAP7_75t_L g390 ( .A(n_384), .Y(n_390) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
BUFx4f_ASAP7_75t_L g558 ( .A(n_384), .Y(n_558) );
BUFx4f_ASAP7_75t_L g889 ( .A(n_384), .Y(n_889) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx3_ASAP7_75t_L g504 ( .A(n_385), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_387), .A2(n_389), .B1(n_783), .B2(n_787), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g795 ( .A1(n_387), .A2(n_389), .B1(n_780), .B2(n_791), .Y(n_795) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_387), .A2(n_389), .B1(n_991), .B2(n_994), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_387), .A2(n_504), .B1(n_989), .B2(n_998), .Y(n_1002) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g942 ( .A(n_388), .Y(n_942) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g844 ( .A(n_390), .Y(n_844) );
INVx1_ASAP7_75t_L g884 ( .A(n_390), .Y(n_884) );
INVx1_ASAP7_75t_L g1403 ( .A(n_390), .Y(n_1403) );
OAI33xp33_ASAP7_75t_L g836 ( .A1(n_391), .A2(n_541), .A3(n_837), .B1(n_841), .B2(n_842), .B3(n_845), .Y(n_836) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g768 ( .A(n_392), .Y(n_768) );
AOI33xp33_ASAP7_75t_L g1052 ( .A1(n_392), .A2(n_684), .A3(n_1053), .B1(n_1055), .B2(n_1057), .B3(n_1058), .Y(n_1052) );
AOI33xp33_ASAP7_75t_L g1459 ( .A1(n_392), .A2(n_1460), .A3(n_1461), .B1(n_1462), .B2(n_1466), .B3(n_1467), .Y(n_1459) );
AND2x4_ASAP7_75t_L g564 ( .A(n_393), .B(n_565), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_393), .A2(n_554), .B1(n_884), .B2(n_885), .C(n_886), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g796 ( .A1(n_395), .A2(n_785), .B1(n_788), .B2(n_797), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_395), .A2(n_828), .B1(n_832), .B2(n_838), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_395), .A2(n_838), .B1(n_926), .B2(n_936), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_395), .A2(n_797), .B1(n_992), .B2(n_995), .Y(n_1003) );
OAI31xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_403), .A3(n_418), .B(n_421), .Y(n_396) );
INVx2_ASAP7_75t_SL g520 ( .A(n_398), .Y(n_520) );
INVx2_ASAP7_75t_SL g629 ( .A(n_398), .Y(n_629) );
INVx1_ASAP7_75t_L g905 ( .A(n_398), .Y(n_905) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_400), .A2(n_874), .B1(n_905), .B2(n_906), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g1453 ( .A1(n_400), .A2(n_520), .B1(n_1442), .B2(n_1443), .Y(n_1453) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AND2x4_ASAP7_75t_L g522 ( .A(n_401), .B(n_402), .Y(n_522) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_402), .Y(n_484) );
INVx2_ASAP7_75t_L g595 ( .A(n_402), .Y(n_595) );
BUFx6f_ASAP7_75t_L g1012 ( .A(n_402), .Y(n_1012) );
OAI22xp33_ASAP7_75t_L g604 ( .A1(n_404), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g1370 ( .A1(n_404), .A2(n_1371), .B1(n_1372), .B2(n_1373), .Y(n_1370) );
NAND3xp33_ASAP7_75t_L g979 ( .A(n_405), .B(n_980), .C(n_982), .Y(n_979) );
NAND3xp33_ASAP7_75t_SL g1025 ( .A(n_405), .B(n_1026), .C(n_1030), .Y(n_1025) );
NAND3xp33_ASAP7_75t_SL g1077 ( .A(n_405), .B(n_1078), .C(n_1079), .Y(n_1077) );
CKINVDCx8_ASAP7_75t_R g405 ( .A(n_406), .Y(n_405) );
CKINVDCx8_ASAP7_75t_R g526 ( .A(n_406), .Y(n_526) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_406), .A2(n_647), .B(n_648), .C(n_649), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g899 ( .A(n_406), .B(n_900), .C(n_903), .Y(n_899) );
NOR3xp33_ASAP7_75t_L g1112 ( .A(n_406), .B(n_1113), .C(n_1115), .Y(n_1112) );
NOR3xp33_ASAP7_75t_L g1454 ( .A(n_406), .B(n_1455), .C(n_1457), .Y(n_1454) );
BUFx2_ASAP7_75t_L g480 ( .A(n_407), .Y(n_480) );
BUFx2_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
BUFx2_ASAP7_75t_L g648 ( .A(n_407), .Y(n_648) );
BUFx3_ASAP7_75t_L g699 ( .A(n_407), .Y(n_699) );
BUFx2_ASAP7_75t_L g912 ( .A(n_407), .Y(n_912) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_407), .Y(n_1010) );
INVx2_ASAP7_75t_L g1029 ( .A(n_407), .Y(n_1029) );
INVx1_ASAP7_75t_L g695 ( .A(n_408), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g409 ( .A1(n_410), .A2(n_414), .B1(n_415), .B2(n_417), .Y(n_409) );
INVx1_ASAP7_75t_L g650 ( .A(n_410), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g859 ( .A1(n_410), .A2(n_813), .B1(n_850), .B2(n_860), .Y(n_859) );
AOI222xp33_ASAP7_75t_L g947 ( .A1(n_410), .A2(n_415), .B1(n_480), .B2(n_948), .C1(n_949), .C2(n_950), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_410), .A2(n_415), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_410), .A2(n_415), .B1(n_1072), .B2(n_1080), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1456 ( .A(n_410), .B(n_1447), .Y(n_1456) );
AND2x4_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
AND2x2_ASAP7_75t_L g415 ( .A(n_411), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g529 ( .A(n_411), .B(n_413), .Y(n_529) );
AND2x4_ASAP7_75t_L g531 ( .A(n_411), .B(n_416), .Y(n_531) );
AND2x4_ASAP7_75t_L g718 ( .A(n_411), .B(n_413), .Y(n_718) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g813 ( .A(n_412), .B(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_414), .A2(n_445), .B1(n_448), .B2(n_453), .Y(n_444) );
INVx1_ASAP7_75t_L g651 ( .A(n_415), .Y(n_651) );
AOI32xp33_ASAP7_75t_L g812 ( .A1(n_415), .A2(n_803), .A3(n_813), .B1(n_815), .B2(n_817), .Y(n_812) );
INVxp67_ASAP7_75t_L g858 ( .A(n_415), .Y(n_858) );
INVxp67_ASAP7_75t_L g902 ( .A(n_415), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_415), .A2(n_718), .B1(n_972), .B2(n_981), .Y(n_980) );
INVx2_ASAP7_75t_SL g537 ( .A(n_419), .Y(n_537) );
BUFx2_ASAP7_75t_L g1114 ( .A(n_419), .Y(n_1114) );
INVx1_ASAP7_75t_L g535 ( .A(n_420), .Y(n_535) );
INVx1_ASAP7_75t_L g636 ( .A(n_420), .Y(n_636) );
INVx2_ASAP7_75t_L g953 ( .A(n_420), .Y(n_953) );
BUFx3_ASAP7_75t_L g1413 ( .A(n_420), .Y(n_1413) );
OAI31xp33_ASAP7_75t_SL g808 ( .A1(n_421), .A2(n_809), .A3(n_810), .B(n_818), .Y(n_808) );
OAI31xp33_ASAP7_75t_SL g854 ( .A1(n_421), .A2(n_855), .A3(n_856), .B(n_857), .Y(n_854) );
OAI21xp5_ASAP7_75t_L g945 ( .A1(n_421), .A2(n_946), .B(n_951), .Y(n_945) );
OAI31xp33_ASAP7_75t_L g976 ( .A1(n_421), .A2(n_977), .A3(n_979), .B(n_984), .Y(n_976) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
AND2x2_ASAP7_75t_SL g538 ( .A(n_422), .B(n_424), .Y(n_538) );
AND2x2_ASAP7_75t_L g722 ( .A(n_422), .B(n_424), .Y(n_722) );
AND2x4_ASAP7_75t_L g1118 ( .A(n_422), .B(n_424), .Y(n_1118) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI31xp33_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_436), .A3(n_454), .B(n_457), .Y(n_426) );
INVx1_ASAP7_75t_L g657 ( .A(n_428), .Y(n_657) );
INVx1_ASAP7_75t_L g1037 ( .A(n_428), .Y(n_1037) );
BUFx3_ASAP7_75t_L g561 ( .A(n_429), .Y(n_561) );
INVx2_ASAP7_75t_SL g762 ( .A(n_429), .Y(n_762) );
BUFx3_ASAP7_75t_L g838 ( .A(n_429), .Y(n_838) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_429), .Y(n_944) );
INVx4_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_431), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_431), .A2(n_644), .B1(n_645), .B2(n_657), .Y(n_656) );
INVx3_ASAP7_75t_SL g866 ( .A(n_431), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_431), .A2(n_1036), .B1(n_1037), .B2(n_1038), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_431), .A2(n_1037), .B1(n_1442), .B2(n_1443), .Y(n_1441) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g676 ( .A(n_434), .Y(n_676) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_434), .Y(n_689) );
INVx2_ASAP7_75t_L g1141 ( .A(n_434), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_437), .A2(n_927), .B1(n_937), .B2(n_942), .Y(n_941) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_437), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_437), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1087) );
NAND3xp33_ASAP7_75t_SL g955 ( .A(n_438), .B(n_956), .C(n_958), .Y(n_955) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_439), .A2(n_659), .B(n_661), .C(n_662), .Y(n_658) );
INVx2_ASAP7_75t_L g1046 ( .A(n_439), .Y(n_1046) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AND2x2_ASAP7_75t_L g506 ( .A(n_440), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g872 ( .A(n_440), .B(n_447), .Y(n_872) );
INVx1_ASAP7_75t_L g1045 ( .A(n_441), .Y(n_1045) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g660 ( .A(n_442), .Y(n_660) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_443), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_445), .A2(n_450), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_445), .A2(n_717), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_445), .A2(n_448), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI222xp33_ASAP7_75t_L g956 ( .A1(n_445), .A2(n_852), .B1(n_869), .B2(n_949), .C1(n_950), .C2(n_957), .Y(n_956) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
AND2x4_ASAP7_75t_L g576 ( .A(n_446), .B(n_447), .Y(n_576) );
AND2x2_ASAP7_75t_L g666 ( .A(n_446), .B(n_667), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g867 ( .A1(n_446), .A2(n_868), .B(n_869), .C(n_870), .Y(n_867) );
INVx1_ASAP7_75t_L g875 ( .A(n_446), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_448), .A2(n_575), .B1(n_577), .B2(n_578), .Y(n_574) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g664 ( .A(n_450), .Y(n_664) );
BUFx3_ASAP7_75t_L g852 ( .A(n_450), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_450), .A2(n_872), .B1(n_1027), .B2(n_1031), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1446 ( .A1(n_450), .A2(n_872), .B1(n_1447), .B2(n_1448), .Y(n_1446) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g961 ( .A(n_456), .Y(n_961) );
OAI31xp33_ASAP7_75t_SL g497 ( .A1(n_457), .A2(n_498), .A3(n_500), .B(n_511), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g799 ( .A1(n_457), .A2(n_800), .A3(n_804), .B(n_807), .Y(n_799) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx3_ASAP7_75t_L g583 ( .A(n_458), .Y(n_583) );
BUFx2_ASAP7_75t_SL g670 ( .A(n_458), .Y(n_670) );
OAI31xp33_ASAP7_75t_L g846 ( .A1(n_458), .A2(n_847), .A3(n_848), .B(n_853), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g954 ( .A1(n_458), .A2(n_955), .B(n_962), .Y(n_954) );
INVx1_ASAP7_75t_L g1047 ( .A(n_458), .Y(n_1047) );
OAI31xp33_ASAP7_75t_L g1068 ( .A1(n_458), .A2(n_1069), .A3(n_1070), .B(n_1074), .Y(n_1068) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
XNOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_567), .Y(n_463) );
NAND4xp75_ASAP7_75t_L g465 ( .A(n_466), .B(n_497), .C(n_517), .D(n_539), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_481), .B1(n_482), .B2(n_492), .Y(n_467) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_472), .B1(n_473), .B2(n_474), .C(n_475), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_469), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g917 ( .A(n_471), .Y(n_917) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_471), .Y(n_1126) );
INVx1_ASAP7_75t_L g1131 ( .A(n_471), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_472), .A2(n_485), .B1(n_549), .B2(n_552), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_473), .A2(n_483), .B1(n_485), .B2(n_486), .C(n_487), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_473), .A2(n_594), .B1(n_595), .B2(n_596), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_473), .A2(n_598), .B1(n_599), .B2(n_602), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_474), .A2(n_486), .B1(n_561), .B2(n_562), .Y(n_560) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g706 ( .A(n_477), .Y(n_706) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx8_ASAP7_75t_L g490 ( .A(n_478), .Y(n_490) );
BUFx3_ASAP7_75t_L g911 ( .A(n_478), .Y(n_911) );
OAI33xp33_ASAP7_75t_L g1369 ( .A1(n_481), .A2(n_492), .A3(n_1370), .B1(n_1374), .B2(n_1379), .B3(n_1385), .Y(n_1369) );
OAI211xp5_ASAP7_75t_L g908 ( .A1(n_483), .A2(n_909), .B(n_910), .C(n_913), .Y(n_908) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx8_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g920 ( .A(n_490), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_491), .B(n_1073), .Y(n_1078) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g603 ( .A(n_493), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_493), .Y(n_915) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g703 ( .A(n_494), .Y(n_703) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g572 ( .A(n_503), .Y(n_572) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_SL g552 ( .A(n_504), .Y(n_552) );
INVx2_ASAP7_75t_SL g616 ( .A(n_504), .Y(n_616) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g573 ( .A(n_506), .Y(n_573) );
INVx3_ASAP7_75t_L g725 ( .A(n_506), .Y(n_725) );
NOR3xp33_ASAP7_75t_L g1148 ( .A(n_506), .B(n_1149), .C(n_1150), .Y(n_1148) );
BUFx3_ASAP7_75t_L g677 ( .A(n_507), .Y(n_677) );
BUFx3_ASAP7_75t_L g869 ( .A(n_507), .Y(n_869) );
BUFx3_ASAP7_75t_L g1056 ( .A(n_507), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_509), .A2(n_528), .B1(n_530), .B2(n_532), .Y(n_527) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_513), .Y(n_580) );
INVx1_ASAP7_75t_L g1418 ( .A(n_513), .Y(n_1418) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_515), .A2(n_653), .B1(n_654), .B2(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_515), .Y(n_730) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
INVx1_ASAP7_75t_L g806 ( .A(n_516), .Y(n_806) );
OAI31xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_523), .A3(n_533), .B(n_538), .Y(n_517) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_520), .A2(n_522), .B1(n_644), .B2(n_645), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_520), .A2(n_522), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g721 ( .A(n_522), .Y(n_721) );
INVx1_ASAP7_75t_L g978 ( .A(n_522), .Y(n_978) );
INVx1_ASAP7_75t_L g1412 ( .A(n_522), .Y(n_1412) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g592 ( .A(n_525), .Y(n_592) );
INVx2_ASAP7_75t_L g631 ( .A(n_525), .Y(n_631) );
INVx2_ASAP7_75t_L g901 ( .A(n_525), .Y(n_901) );
INVx1_ASAP7_75t_L g1103 ( .A(n_525), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_528), .A2(n_530), .B1(n_577), .B2(n_633), .Y(n_632) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_531), .A2(n_717), .B1(n_718), .B2(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g1116 ( .A(n_531), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_531), .A2(n_718), .B1(n_1409), .B2(n_1410), .Y(n_1408) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_535), .A2(n_537), .B1(n_653), .B2(n_654), .Y(n_652) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g626 ( .A1(n_538), .A2(n_627), .A3(n_630), .B(n_634), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_538), .A2(n_642), .B1(n_655), .B2(n_670), .C(n_671), .Y(n_641) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_538), .A2(n_898), .B(n_907), .Y(n_897) );
OAI31xp33_ASAP7_75t_SL g1404 ( .A1(n_538), .A2(n_1405), .A3(n_1406), .B(n_1411), .Y(n_1404) );
OA33x2_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .A3(n_548), .B1(n_553), .B2(n_560), .B3(n_563), .Y(n_539) );
INVx1_ASAP7_75t_L g1134 ( .A(n_540), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI33xp33_ASAP7_75t_L g608 ( .A1(n_541), .A2(n_609), .A3(n_614), .B1(n_617), .B2(n_621), .B3(n_625), .Y(n_608) );
OAI33xp33_ASAP7_75t_L g1083 ( .A1(n_541), .A2(n_768), .A3(n_1084), .B1(n_1087), .B2(n_1091), .B3(n_1094), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_544), .A2(n_546), .B1(n_881), .B2(n_882), .Y(n_880) );
INVx5_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx6_ASAP7_75t_L g562 ( .A(n_547), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_549), .A2(n_594), .B1(n_598), .B2(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g1395 ( .A(n_550), .Y(n_1395) );
INVx4_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_557), .B1(n_558), .B2(n_559), .Y(n_553) );
INVx4_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g620 ( .A(n_556), .Y(n_620) );
INVx2_ASAP7_75t_L g1089 ( .A(n_556), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_558), .A2(n_843), .B1(n_929), .B2(n_933), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g625 ( .A(n_564), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g686 ( .A(n_564), .B(n_687), .C(n_690), .Y(n_686) );
AOI33xp33_ASAP7_75t_L g1133 ( .A1(n_564), .A2(n_1134), .A3(n_1135), .B1(n_1137), .B2(n_1143), .B3(n_1144), .Y(n_1133) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND3x1_ASAP7_75t_L g568 ( .A(n_569), .B(n_584), .C(n_626), .Y(n_568) );
OAI31xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .A3(n_579), .B(n_583), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g1422 ( .A1(n_575), .A2(n_852), .B1(n_1409), .B2(n_1423), .Y(n_1422) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g663 ( .A(n_576), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_576), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_576), .A2(n_852), .B1(n_972), .B2(n_973), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_576), .A2(n_852), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g1420 ( .A(n_582), .Y(n_1420) );
NOR2xp33_ASAP7_75t_SL g584 ( .A(n_585), .B(n_608), .Y(n_584) );
OAI22xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_591), .B2(n_592), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g609 ( .A1(n_587), .A2(n_606), .B1(n_610), .B2(n_613), .Y(n_609) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_591), .A2(n_607), .B1(n_615), .B2(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_595), .A2(n_827), .B1(n_828), .B2(n_829), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_596), .A2(n_602), .B1(n_622), .B2(n_624), .Y(n_621) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx8_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx5_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_SL g1391 ( .A(n_623), .Y(n_1391) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_707), .B2(n_708), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .C(n_652), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_658), .C(n_665), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g1449 ( .A(n_659), .B(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1142 ( .A(n_660), .Y(n_1142) );
INVx2_ASAP7_75t_L g1465 ( .A(n_660), .Y(n_1465) );
INVx2_ASAP7_75t_L g728 ( .A(n_664), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g958 ( .A1(n_666), .A2(n_959), .B1(n_960), .B2(n_961), .Y(n_958) );
INVx3_ASAP7_75t_L g1060 ( .A(n_667), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx3_ASAP7_75t_L g680 ( .A(n_668), .Y(n_680) );
OAI31xp33_ASAP7_75t_L g723 ( .A1(n_670), .A2(n_724), .A3(n_729), .B(n_731), .Y(n_723) );
OAI31xp33_ASAP7_75t_SL g968 ( .A1(n_670), .A2(n_969), .A3(n_974), .B(n_975), .Y(n_968) );
OAI31xp33_ASAP7_75t_L g1414 ( .A1(n_670), .A2(n_1415), .A3(n_1416), .B(n_1421), .Y(n_1414) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_686), .C(n_691), .D(n_700), .Y(n_671) );
NAND3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_678), .C(n_683), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g894 ( .A(n_680), .Y(n_894) );
INVx2_ASAP7_75t_L g1054 ( .A(n_680), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1145 ( .A(n_680), .Y(n_1145) );
INVx1_ASAP7_75t_L g1468 ( .A(n_680), .Y(n_1468) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_681), .Y(n_1136) );
BUFx3_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g1062 ( .A(n_682), .Y(n_1062) );
BUFx6f_ASAP7_75t_L g1469 ( .A(n_682), .Y(n_1469) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
OAI33xp33_ASAP7_75t_L g759 ( .A1(n_685), .A2(n_760), .A3(n_764), .B1(n_765), .B2(n_766), .B3(n_768), .Y(n_759) );
INVx2_ASAP7_75t_SL g1460 ( .A(n_685), .Y(n_1460) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g1464 ( .A(n_689), .Y(n_1464) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_692), .B(n_696), .C(n_698), .Y(n_691) );
BUFx12f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g914 ( .A(n_694), .Y(n_914) );
INVx5_ASAP7_75t_L g1014 ( .A(n_694), .Y(n_1014) );
INVx1_ASAP7_75t_L g814 ( .A(n_695), .Y(n_814) );
INVx1_ASAP7_75t_L g1015 ( .A(n_696), .Y(n_1015) );
BUFx3_ASAP7_75t_L g1120 ( .A(n_696), .Y(n_1120) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_699), .Y(n_983) );
INVx1_ASAP7_75t_L g1018 ( .A(n_699), .Y(n_1018) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .C(n_704), .Y(n_700) );
BUFx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_723), .C(n_732), .Y(n_710) );
OAI31xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .A3(n_720), .B(n_722), .Y(n_711) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g811 ( .A(n_718), .Y(n_811) );
OAI31xp33_ASAP7_75t_SL g1023 ( .A1(n_722), .A2(n_1024), .A3(n_1025), .B(n_1033), .Y(n_1023) );
OAI31xp33_ASAP7_75t_SL g1075 ( .A1(n_722), .A2(n_1076), .A3(n_1077), .B(n_1081), .Y(n_1075) );
INVx1_ASAP7_75t_L g1458 ( .A(n_722), .Y(n_1458) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_759), .Y(n_732) );
OAI33xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .A3(n_744), .B1(n_748), .B2(n_755), .B3(n_758), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_734), .A2(n_908), .B1(n_915), .B2(n_916), .Y(n_907) );
OAI33xp33_ASAP7_75t_L g924 ( .A1(n_734), .A2(n_758), .A3(n_925), .B1(n_928), .B2(n_931), .B3(n_935), .Y(n_924) );
OAI22xp33_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_740), .B2(n_741), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_736), .A2(n_756), .B1(n_761), .B2(n_763), .Y(n_760) );
BUFx4f_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx2_ASAP7_75t_SL g1099 ( .A(n_739), .Y(n_1099) );
INVxp67_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_746), .A2(n_754), .B1(n_761), .B2(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_747), .A2(n_932), .B1(n_933), .B2(n_934), .Y(n_931) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_751), .B1(n_752), .B2(n_754), .Y(n_748) );
INVx2_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_SL g784 ( .A(n_750), .Y(n_784) );
INVx3_ASAP7_75t_L g932 ( .A(n_750), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g928 ( .A1(n_752), .A2(n_917), .B1(n_929), .B2(n_930), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_752), .A2(n_784), .B1(n_994), .B2(n_995), .Y(n_993) );
BUFx3_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g1022 ( .A(n_758), .Y(n_1022) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g1393 ( .A(n_767), .Y(n_1393) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OA22x2_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_963), .B1(n_964), .B2(n_1153), .Y(n_770) );
INVx1_ASAP7_75t_L g1153 ( .A(n_771), .Y(n_1153) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
XNOR2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_861), .Y(n_772) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_819), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_799), .C(n_808), .Y(n_775) );
NOR2xp33_ASAP7_75t_SL g776 ( .A(n_777), .B(n_792), .Y(n_776) );
INVx1_ASAP7_75t_L g1383 ( .A(n_781), .Y(n_1383) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1402 ( .A(n_798), .Y(n_1402) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g877 ( .A(n_806), .B(n_878), .Y(n_877) );
INVx3_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_846), .C(n_854), .Y(n_820) );
NOR2xp33_ASAP7_75t_SL g821 ( .A(n_822), .B(n_836), .Y(n_821) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_824), .A2(n_834), .B1(n_838), .B2(n_839), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g842 ( .A1(n_825), .A2(n_835), .B1(n_843), .B2(n_844), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_829), .A2(n_1386), .B1(n_1387), .B2(n_1388), .Y(n_1385) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_839), .A2(n_930), .B1(n_934), .B2(n_944), .Y(n_943) );
BUFx6f_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g1398 ( .A(n_843), .Y(n_1398) );
XOR2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_921), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_895), .B(n_897), .Y(n_863) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_883), .B(n_887), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g916 ( .A1(n_882), .A2(n_888), .B1(n_917), .B2(n_918), .C(n_919), .Y(n_916) );
OAI211xp5_ASAP7_75t_SL g887 ( .A1(n_888), .A2(n_889), .B(n_890), .C(n_893), .Y(n_887) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
BUFx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_SL g898 ( .A(n_899), .B(n_904), .Y(n_898) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_911), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_912), .Y(n_1129) );
INVx1_ASAP7_75t_L g1132 ( .A(n_915), .Y(n_1132) );
NAND3xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_945), .C(n_954), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g923 ( .A(n_924), .B(n_938), .Y(n_923) );
INVx2_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
XNOR2xp5_ASAP7_75t_L g964 ( .A(n_965), .B(n_1004), .Y(n_964) );
INVx2_ASAP7_75t_SL g965 ( .A(n_966), .Y(n_965) );
NAND3xp33_ASAP7_75t_L g967 ( .A(n_968), .B(n_976), .C(n_985), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_973), .B(n_983), .Y(n_982) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_999), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1104), .B1(n_1151), .B2(n_1152), .Y(n_1004) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1005), .Y(n_1152) );
XNOR2x1_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1066), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1048), .Y(n_1006) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1008), .Y(n_1050) );
AOI21xp5_ASAP7_75t_L g1008 ( .A1(n_1009), .A2(n_1011), .B(n_1016), .Y(n_1008) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1014), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_1018), .A2(n_1019), .B1(n_1020), .B2(n_1021), .C(n_1022), .Y(n_1017) );
INVx2_ASAP7_75t_L g1123 ( .A(n_1020), .Y(n_1123) );
AOI32xp33_ASAP7_75t_L g1470 ( .A1(n_1022), .A2(n_1471), .A3(n_1474), .B1(n_1475), .B2(n_1476), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1023), .B(n_1034), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_1027), .B(n_1028), .Y(n_1026) );
INVx2_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_1032), .B(n_1044), .Y(n_1043) );
AO21x1_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1039), .B(n_1047), .Y(n_1034) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1041), .Y(n_1039) );
NAND3xp33_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .C(n_1046), .Y(n_1041) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
NAND3xp33_ASAP7_75t_L g1445 ( .A(n_1046), .B(n_1446), .C(n_1449), .Y(n_1445) );
AO21x1_ASAP7_75t_L g1146 ( .A1(n_1047), .A2(n_1147), .B(n_1148), .Y(n_1146) );
AO21x1_ASAP7_75t_L g1440 ( .A1(n_1047), .A2(n_1441), .B(n_1444), .Y(n_1440) );
OAI31xp33_ASAP7_75t_L g1048 ( .A1(n_1049), .A2(n_1050), .A3(n_1051), .B(n_1063), .Y(n_1048) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1052), .Y(n_1065) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1064), .B(n_1065), .Y(n_1063) );
NAND3xp33_ASAP7_75t_SL g1067 ( .A(n_1068), .B(n_1075), .C(n_1082), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1097), .Y(n_1082) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1106), .Y(n_1151) );
NAND4xp25_ASAP7_75t_SL g1107 ( .A(n_1108), .B(n_1119), .C(n_1133), .D(n_1146), .Y(n_1107) );
AO21x1_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1112), .B(n_1117), .Y(n_1108) );
CKINVDCx14_ASAP7_75t_R g1117 ( .A(n_1118), .Y(n_1117) );
AOI33xp33_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1121), .A3(n_1124), .B1(n_1128), .B2(n_1130), .B3(n_1132), .Y(n_1119) );
BUFx2_ASAP7_75t_SL g1122 ( .A(n_1123), .Y(n_1122) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1131), .Y(n_1380) );
INVx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx2_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_1155), .A2(n_1364), .B1(n_1366), .B2(n_1424), .C(n_1429), .Y(n_1154) );
NOR3xp33_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1302), .C(n_1344), .Y(n_1155) );
A2O1A1Ixp33_ASAP7_75t_L g1156 ( .A1(n_1157), .A2(n_1236), .B(n_1254), .C(n_1258), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1183), .B1(n_1191), .B2(n_1202), .C(n_1209), .Y(n_1157) );
AOI221xp5_ASAP7_75t_SL g1303 ( .A1(n_1158), .A2(n_1242), .B1(n_1304), .B2(n_1306), .C(n_1308), .Y(n_1303) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1174), .Y(n_1159) );
INVx3_ASAP7_75t_L g1235 ( .A(n_1160), .Y(n_1235) );
NOR2xp33_ASAP7_75t_L g1244 ( .A(n_1160), .B(n_1225), .Y(n_1244) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1160), .B(n_1175), .Y(n_1246) );
INVx3_ASAP7_75t_L g1260 ( .A(n_1160), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1160), .B(n_1268), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1160), .B(n_1216), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1160), .B(n_1175), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1160), .B(n_1223), .Y(n_1363) );
AND2x4_ASAP7_75t_SL g1160 ( .A(n_1161), .B(n_1168), .Y(n_1160) );
AND2x6_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1164), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1163), .B(n_1167), .Y(n_1166) );
AND2x4_ASAP7_75t_L g1169 ( .A(n_1163), .B(n_1170), .Y(n_1169) );
AND2x6_ASAP7_75t_L g1172 ( .A(n_1163), .B(n_1173), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1163), .B(n_1167), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1163), .B(n_1167), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1165), .B(n_1171), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1365 ( .A(n_1166), .Y(n_1365) );
OAI21xp5_ASAP7_75t_L g1479 ( .A1(n_1167), .A2(n_1480), .B(n_1481), .Y(n_1479) );
INVx2_ASAP7_75t_SL g1295 ( .A(n_1174), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1179), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_1175), .B(n_1204), .Y(n_1203) );
NAND2xp5_ASAP7_75t_SL g1210 ( .A(n_1175), .B(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1175), .B(n_1180), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1175), .B(n_1235), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1175), .B(n_1180), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1343 ( .A(n_1175), .B(n_1255), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1178), .Y(n_1175) );
AND2x4_ASAP7_75t_L g1264 ( .A(n_1176), .B(n_1178), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1179), .B(n_1264), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1179), .B(n_1231), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_1179), .B(n_1206), .Y(n_1336) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1180), .Y(n_1216) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1180), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1182), .Y(n_1180) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1183), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1252 ( .A(n_1183), .B(n_1253), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1183), .B(n_1219), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1183), .B(n_1271), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1188), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1184), .B(n_1201), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1243 ( .A(n_1184), .B(n_1188), .Y(n_1243) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1184), .Y(n_1285) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1185), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1240 ( .A(n_1185), .B(n_1188), .Y(n_1240) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1187), .Y(n_1185) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1188), .Y(n_1201) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1188), .Y(n_1233) );
NOR2xp33_ASAP7_75t_L g1347 ( .A(n_1188), .B(n_1214), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1198), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_1192), .A2(n_1266), .B1(n_1328), .B2(n_1362), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1197), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1193), .B(n_1200), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1193), .B(n_1252), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1196), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1194), .B(n_1196), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1221 ( .A(n_1197), .B(n_1222), .Y(n_1221) );
A2O1A1Ixp33_ASAP7_75t_L g1287 ( .A1(n_1198), .A2(n_1288), .B(n_1290), .C(n_1294), .Y(n_1287) );
OAI221xp5_ASAP7_75t_L g1327 ( .A1(n_1198), .A2(n_1328), .B1(n_1329), .B2(n_1330), .C(n_1331), .Y(n_1327) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1199), .B(n_1231), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1218 ( .A(n_1200), .B(n_1219), .Y(n_1218) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1200), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1200), .B(n_1222), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1201), .B(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1204), .B(n_1232), .Y(n_1267) );
AOI32xp33_ASAP7_75t_L g1276 ( .A1(n_1204), .A2(n_1277), .A3(n_1281), .B1(n_1282), .B2(n_1286), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1204), .B(n_1319), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1204), .B(n_1240), .Y(n_1329) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1205), .B(n_1239), .Y(n_1238) );
NAND2xp5_ASAP7_75t_SL g1262 ( .A(n_1205), .B(n_1263), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1205), .B(n_1292), .Y(n_1291) );
NAND2xp5_ASAP7_75t_SL g1353 ( .A(n_1205), .B(n_1242), .Y(n_1353) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1206), .B(n_1216), .Y(n_1215) );
NOR2xp33_ASAP7_75t_L g1219 ( .A(n_1206), .B(n_1214), .Y(n_1219) );
INVx3_ASAP7_75t_L g1231 ( .A(n_1206), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1206), .B(n_1214), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1206), .B(n_1235), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1208), .Y(n_1206) );
NAND3xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1217), .C(n_1224), .Y(n_1209) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1215), .Y(n_1211) );
CKINVDCx14_ASAP7_75t_R g1212 ( .A(n_1213), .Y(n_1212) );
AOI32xp33_ASAP7_75t_L g1294 ( .A1(n_1213), .A2(n_1295), .A3(n_1296), .B1(n_1297), .B2(n_1301), .Y(n_1294) );
CKINVDCx5p33_ASAP7_75t_R g1222 ( .A(n_1214), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_1214), .B(n_1229), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1214), .B(n_1233), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1214), .B(n_1240), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1214), .B(n_1285), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1214), .B(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1216), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1216), .B(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1216), .Y(n_1299) );
OAI322xp33_ASAP7_75t_L g1308 ( .A1(n_1216), .A2(n_1265), .A3(n_1268), .B1(n_1309), .B2(n_1310), .C1(n_1313), .C2(n_1314), .Y(n_1308) );
O2A1O1Ixp33_ASAP7_75t_L g1337 ( .A1(n_1216), .A2(n_1338), .B(n_1339), .C(n_1342), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1348 ( .A1(n_1216), .A2(n_1220), .B1(n_1349), .B2(n_1351), .Y(n_1348) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1216), .B(n_1350), .Y(n_1349) );
OAI21xp5_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1220), .B(n_1223), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1219), .B(n_1242), .Y(n_1301) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1222), .B(n_1242), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1222), .B(n_1278), .Y(n_1277) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1222), .B(n_1285), .Y(n_1289) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1222), .B(n_1353), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1222), .B(n_1240), .Y(n_1360) );
AOI222xp33_ASAP7_75t_L g1345 ( .A1(n_1223), .A2(n_1239), .B1(n_1263), .B2(n_1271), .C1(n_1295), .C2(n_1346), .Y(n_1345) );
A2O1A1Ixp33_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1227), .B(n_1230), .C(n_1234), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1225), .B(n_1234), .Y(n_1286) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1226), .B(n_1239), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1226), .B(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1229), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1232), .Y(n_1230) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1231), .Y(n_1253) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1233), .Y(n_1307) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1234), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1235), .B(n_1292), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1235), .B(n_1293), .Y(n_1328) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1235), .B(n_1279), .C(n_1336), .Y(n_1335) );
NOR2xp33_ASAP7_75t_L g1356 ( .A(n_1235), .B(n_1357), .Y(n_1356) );
O2A1O1Ixp33_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1241), .B(n_1244), .C(n_1245), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1240), .B(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1240), .Y(n_1280) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1241), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1242), .B(n_1271), .Y(n_1350) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
OAI21xp5_ASAP7_75t_L g1245 ( .A1(n_1246), .A2(n_1247), .B(n_1248), .Y(n_1245) );
A2O1A1Ixp33_ASAP7_75t_L g1297 ( .A1(n_1246), .A2(n_1298), .B(n_1299), .C(n_1300), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1250), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1249), .B(n_1253), .Y(n_1334) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1283 ( .A(n_1253), .B(n_1284), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1253), .B(n_1347), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1254), .B(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1254), .Y(n_1298) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_1254), .A2(n_1324), .B1(n_1325), .B2(n_1327), .C(n_1337), .Y(n_1323) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_1255), .A2(n_1298), .B1(n_1303), .B2(n_1315), .C(n_1323), .Y(n_1302) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1255), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1256), .B(n_1257), .Y(n_1255) );
AOI211xp5_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1261), .B(n_1272), .C(n_1287), .Y(n_1258) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1260), .Y(n_1313) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_1262), .A2(n_1265), .B1(n_1266), .B2(n_1268), .C(n_1269), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1263), .B(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1263), .Y(n_1317) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1264), .Y(n_1268) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1264), .B(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
OAI21xp33_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1274), .B(n_1276), .Y(n_1272) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1275), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1280), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_1279), .B(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1281), .Y(n_1330) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1296), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1298), .B(n_1313), .Y(n_1354) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1299), .B(n_1321), .Y(n_1320) );
INVxp67_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
AOI31xp33_ASAP7_75t_SL g1331 ( .A1(n_1307), .A2(n_1332), .A3(n_1334), .B(n_1335), .Y(n_1331) );
INVxp67_ASAP7_75t_SL g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1312), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1320), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1317), .B(n_1318), .Y(n_1316) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
AOI211xp5_ASAP7_75t_L g1355 ( .A1(n_1322), .A2(n_1343), .B(n_1356), .C(n_1361), .Y(n_1355) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
A2O1A1Ixp33_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1348), .B(n_1354), .C(n_1355), .Y(n_1344) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVxp67_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1359), .B(n_1360), .Y(n_1358) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
INVx4_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
NAND3xp33_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1404), .C(n_1414), .Y(n_1367) );
NOR2xp33_ASAP7_75t_SL g1368 ( .A(n_1369), .B(n_1389), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_1371), .A2(n_1387), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_1373), .A2(n_1388), .B1(n_1392), .B2(n_1397), .Y(n_1396) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
OAI22xp33_ASAP7_75t_L g1399 ( .A1(n_1378), .A2(n_1384), .B1(n_1400), .B2(n_1403), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1381), .B1(n_1382), .B2(n_1384), .Y(n_1379) );
INVx2_ASAP7_75t_SL g1382 ( .A(n_1383), .Y(n_1382) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx3_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
CKINVDCx20_ASAP7_75t_R g1424 ( .A(n_1425), .Y(n_1424) );
CKINVDCx20_ASAP7_75t_R g1425 ( .A(n_1426), .Y(n_1425) );
INVx3_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
HB1xp67_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
BUFx3_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVxp33_ASAP7_75t_SL g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
NAND4xp75_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1452), .C(n_1459), .D(n_1470), .Y(n_1439) );
NOR2xp33_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1451), .Y(n_1444) );
AO21x1_ASAP7_75t_L g1452 ( .A1(n_1453), .A2(n_1454), .B(n_1458), .Y(n_1452) );
INVx2_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx2_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
endmodule