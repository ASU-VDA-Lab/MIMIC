module real_jpeg_4646_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_1),
.A2(n_39),
.B1(n_47),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_1),
.A2(n_47),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_1),
.A2(n_47),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_2),
.A2(n_250),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_2),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_2),
.A2(n_100),
.B1(n_287),
.B2(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_2),
.A2(n_287),
.B1(n_387),
.B2(n_390),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_2),
.A2(n_219),
.B1(n_287),
.B2(n_404),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_3),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_4),
.A2(n_179),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_4),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_4),
.A2(n_194),
.B1(n_236),
.B2(n_277),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g393 ( 
.A1(n_4),
.A2(n_236),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_4),
.A2(n_236),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_5),
.A2(n_98),
.B1(n_99),
.B2(n_101),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_5),
.A2(n_98),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_5),
.A2(n_98),
.B1(n_131),
.B2(n_142),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_5),
.A2(n_98),
.B1(n_266),
.B2(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_7),
.A2(n_69),
.B1(n_91),
.B2(n_111),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_7),
.A2(n_69),
.B1(n_130),
.B2(n_136),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_7),
.A2(n_69),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_75),
.B1(n_79),
.B2(n_80),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_8),
.A2(n_79),
.B1(n_128),
.B2(n_131),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_8),
.A2(n_48),
.B1(n_79),
.B2(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_8),
.A2(n_79),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_9),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_9),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_10),
.A2(n_130),
.B1(n_281),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_10),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_10),
.A2(n_112),
.B1(n_284),
.B2(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_10),
.A2(n_48),
.B1(n_284),
.B2(n_379),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_10),
.A2(n_284),
.B1(n_414),
.B2(n_416),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_11),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_11),
.Y(n_144)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_14),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_14),
.Y(n_136)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_14),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_14),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_14),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_14),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_17),
.B(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_17),
.A2(n_142),
.B(n_259),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_17),
.B(n_198),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_17),
.B(n_363),
.C(n_367),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_17),
.A2(n_373),
.B1(n_374),
.B2(n_377),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_17),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_17),
.B(n_96),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_17),
.A2(n_148),
.B1(n_413),
.B2(n_421),
.Y(n_420)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_202),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_200),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_182),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_27),
.B(n_182),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_27),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_27),
.B(n_204),
.Y(n_488)
);

FAx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_103),
.CI(n_146),
.CON(n_27),
.SN(n_27)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_28),
.A2(n_29),
.B(n_72),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_72),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_50),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_30),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_31),
.A2(n_42),
.B(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_31),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_31),
.A2(n_51),
.B1(n_63),
.B2(n_228),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_31),
.B(n_373),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g398 ( 
.A(n_38),
.Y(n_398)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_38),
.Y(n_429)
);

INVx8_ASAP7_75t_L g266 ( 
.A(n_39),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_39),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_42),
.A2(n_51),
.B(n_172),
.Y(n_292)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_43),
.Y(n_170)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_45),
.Y(n_230)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_45),
.Y(n_361)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_45),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_45),
.Y(n_459)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_46),
.Y(n_377)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_46),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g390 ( 
.A(n_46),
.Y(n_390)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_46),
.Y(n_450)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_48),
.Y(n_171)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_82)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_49),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_63),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_51),
.A2(n_168),
.B(n_172),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_51),
.A2(n_471),
.B(n_472),
.Y(n_470)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_52),
.A2(n_169),
.B1(n_173),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_52),
.A2(n_173),
.B1(n_372),
.B2(n_378),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_52),
.A2(n_173),
.B1(n_378),
.B2(n_386),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_52),
.A2(n_173),
.B1(n_386),
.B2(n_456),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_58),
.B2(n_61),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g366 ( 
.A(n_60),
.Y(n_366)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_64),
.B(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_71),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_81),
.B1(n_96),
.B2(n_97),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_74),
.A2(n_82),
.B(n_195),
.Y(n_239)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_77),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_77),
.Y(n_443)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_78),
.Y(n_249)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_97),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_81),
.B(n_110),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_81),
.A2(n_191),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_81),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_81),
.A2(n_96),
.B1(n_331),
.B2(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_90),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_82),
.B(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_82),
.A2(n_297),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_82),
.A2(n_297),
.B1(n_301),
.B2(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_86),
.Y(n_446)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_92),
.Y(n_193)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_94),
.Y(n_255)
);

INVx6_ASAP7_75t_L g440 ( 
.A(n_95),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_110),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g454 ( 
.A1(n_99),
.A2(n_373),
.B(n_441),
.Y(n_454)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_102),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_116),
.B2(n_145),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_114),
.B2(n_115),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_106),
.A2(n_115),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_107),
.B(n_115),
.C(n_116),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_109),
.A2(n_192),
.B(n_301),
.Y(n_316)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g437 ( 
.A1(n_112),
.A2(n_438),
.A3(n_440),
.B1(n_441),
.B2(n_444),
.Y(n_437)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_145),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_127),
.B(n_133),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_135),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_117),
.A2(n_138),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_117),
.A2(n_138),
.B1(n_233),
.B2(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_126),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_127),
.Y(n_197)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_130),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_137),
.A2(n_175),
.B(n_181),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_137),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_137),
.A2(n_198),
.B1(n_280),
.B2(n_285),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_138),
.A2(n_233),
.B(n_237),
.Y(n_232)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_166),
.B(n_174),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_174),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_147),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_147),
.A2(n_167),
.B1(n_207),
.B2(n_342),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_157),
.B(n_161),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_148),
.B(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_148),
.A2(n_263),
.B1(n_269),
.B2(n_271),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_148),
.A2(n_271),
.B(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_148),
.A2(n_222),
.B(n_393),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_148),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_148),
.A2(n_403),
.B1(n_413),
.B2(n_417),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_148),
.A2(n_161),
.B(n_305),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_149),
.Y(n_404)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_151),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_153),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_154),
.B(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_154),
.A2(n_214),
.B(n_264),
.Y(n_326)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_156),
.Y(n_425)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_157),
.Y(n_407)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_206),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_167),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_175),
.B(n_198),
.Y(n_237)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_240),
.B(n_487),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_209),
.C(n_210),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_205),
.B(n_209),
.CI(n_210),
.CON(n_350),
.SN(n_350)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_231),
.C(n_238),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_211),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_225),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_212),
.A2(n_225),
.B1(n_226),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_212),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_215),
.Y(n_306)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_221),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_231),
.A2(n_232),
.B1(n_238),
.B2(n_239),
.Y(n_344)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_351),
.B(n_481),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_336),
.C(n_348),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_320),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_243),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_308),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_244),
.B(n_308),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_291),
.C(n_303),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_245),
.B(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_274),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_246),
.B(n_275),
.C(n_279),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_262),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_247),
.B(n_262),
.Y(n_323)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_250),
.A3(n_252),
.B1(n_254),
.B2(n_258),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx8_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_303),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.C(n_296),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_292),
.B(n_293),
.CI(n_296),
.CON(n_322),
.SN(n_322)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_304),
.B(n_307),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_311),
.C(n_313),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_318),
.C(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_334),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_321),
.B(n_334),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.C(n_324),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_322),
.B(n_479),
.Y(n_478)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_322),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_323),
.B(n_324),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.C(n_329),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_466)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_329),
.B(n_466),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

A2O1A1O1Ixp25_ASAP7_75t_L g481 ( 
.A1(n_336),
.A2(n_348),
.B(n_482),
.C(n_485),
.D(n_486),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_347),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_337),
.B(n_347),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_341),
.C(n_346),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_343),
.B1(n_345),
.B2(n_346),
.Y(n_340)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_341),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_349),
.B(n_350),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_350),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_352),
.A2(n_476),
.B(n_480),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_353),
.A2(n_461),
.B(n_475),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_433),
.B(n_460),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_399),
.B(n_432),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_381),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_356),
.B(n_381),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_371),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_371),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_373),
.B(n_442),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_392),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_384),
.B1(n_385),
.B2(n_391),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_383),
.B(n_391),
.C(n_392),
.Y(n_434)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_385),
.Y(n_391)
);

INVx4_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_409),
.B(n_431),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_408),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_401),
.B(n_408),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_405),
.B1(n_406),
.B2(n_407),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_419),
.B(n_430),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_411),
.B(n_412),
.Y(n_430)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_417),
.Y(n_422)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_423),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_434),
.B(n_435),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_452),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_453),
.C(n_455),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_451),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_451),
.Y(n_469)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

INVx6_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_449),
.Y(n_457)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_455),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_456),
.Y(n_471)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_462),
.B(n_463),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_464),
.A2(n_465),
.B1(n_467),
.B2(n_468),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_470),
.C(n_473),
.Y(n_477)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_473),
.B2(n_474),
.Y(n_468)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_469),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_470),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_478),
.Y(n_480)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);


endmodule