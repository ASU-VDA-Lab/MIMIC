module fake_jpeg_32028_n_114 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_114);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_19),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_30),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

CKINVDCx12_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_37),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_48),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_3),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_50),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_70),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_43),
.B(n_1),
.C(n_2),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_76),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_60),
.A2(n_65),
.B1(n_71),
.B2(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_83),
.B1(n_9),
.B2(n_10),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_38),
.C(n_42),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_80),
.C(n_81),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_0),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_46),
.B(n_20),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_17),
.C(n_34),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_16),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_79),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_88),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_81),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_86),
.A2(n_14),
.B1(n_15),
.B2(n_23),
.Y(n_97)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_8),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_95),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_12),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_29),
.C(n_32),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_102),
.B1(n_84),
.B2(n_96),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_106),
.A2(n_99),
.B1(n_104),
.B2(n_100),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_109),
.C(n_94),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_101),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_109),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

AOI211xp5_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_105),
.B(n_103),
.C(n_85),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_98),
.Y(n_114)
);


endmodule