module real_jpeg_5207_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_0),
.A2(n_96),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_0),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_0),
.A2(n_288),
.B1(n_293),
.B2(n_306),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_0),
.A2(n_125),
.B1(n_306),
.B2(n_389),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_0),
.A2(n_34),
.B1(n_306),
.B2(n_468),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_1),
.A2(n_61),
.B1(n_147),
.B2(n_177),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_1),
.A2(n_61),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_1),
.A2(n_61),
.B1(n_397),
.B2(n_399),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_93),
.B1(n_95),
.B2(n_98),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_2),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_2),
.A2(n_98),
.B1(n_146),
.B2(n_150),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_2),
.A2(n_98),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_3),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_137),
.B1(n_166),
.B2(n_169),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_3),
.A2(n_137),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_4),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_4),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_4),
.Y(n_237)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_4),
.Y(n_319)
);

INVx8_ASAP7_75t_L g334 ( 
.A(n_4),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_4),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_5),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_5),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_5),
.A2(n_209),
.B1(n_241),
.B2(n_276),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_5),
.A2(n_209),
.B1(n_297),
.B2(n_301),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_5),
.A2(n_135),
.B1(n_151),
.B2(n_209),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_6),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_6),
.Y(n_214)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_7),
.Y(n_418)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_8),
.Y(n_515)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_125),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_13),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_13),
.A2(n_127),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_13),
.A2(n_127),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g425 ( 
.A1(n_13),
.A2(n_127),
.B1(n_426),
.B2(n_430),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_14),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_14),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_14),
.A2(n_255),
.B1(n_288),
.B2(n_293),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_14),
.A2(n_93),
.B1(n_255),
.B2(n_346),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_14),
.A2(n_255),
.B1(n_419),
.B2(n_443),
.Y(n_442)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_16),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_16),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_16),
.B(n_283),
.C(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_16),
.B(n_116),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_16),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_16),
.B(n_91),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_16),
.B(n_356),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_17),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_18),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_18),
.A2(n_50),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_18),
.A2(n_50),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_18),
.A2(n_50),
.B1(n_241),
.B2(n_447),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_513),
.B(n_516),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_216),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_215),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_159),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_24),
.B(n_159),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_138),
.B2(n_139),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_62),
.C(n_99),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_27),
.A2(n_140),
.B1(n_141),
.B2(n_158),
.Y(n_139)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_27),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_27),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_28),
.A2(n_53),
.B1(n_55),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_28),
.A2(n_253),
.B(n_258),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_28),
.A2(n_38),
.B1(n_253),
.B2(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_29),
.B(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_29),
.A2(n_438),
.B(n_439),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_35),
.Y(n_468)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_38),
.B(n_273),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_41),
.Y(n_251)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_42),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_42),
.Y(n_444)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_43),
.Y(n_115)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_44),
.Y(n_135)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_44),
.Y(n_414)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g410 ( 
.A1(n_46),
.A2(n_411),
.A3(n_415),
.B1(n_416),
.B2(n_420),
.Y(n_410)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_49),
.B(n_54),
.Y(n_206)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_51),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_53),
.A2(n_207),
.B(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_54),
.B(n_208),
.Y(n_258)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_63),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_62),
.A2(n_63),
.B1(n_99),
.B2(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_90),
.B(n_92),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_64),
.A2(n_269),
.B(n_274),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_64),
.A2(n_90),
.B1(n_305),
.B2(n_345),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_64),
.A2(n_274),
.B(n_345),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_64),
.A2(n_90),
.B1(n_446),
.B2(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_65),
.A2(n_91),
.B1(n_165),
.B2(n_172),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_65),
.A2(n_91),
.B1(n_165),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_65),
.A2(n_91),
.B1(n_200),
.B2(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_65),
.B(n_275),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_80),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B1(n_75),
.B2(n_78),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_69),
.Y(n_281)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_70),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_70),
.Y(n_272)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_71),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_71),
.Y(n_350)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_79),
.Y(n_308)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_80),
.A2(n_305),
.B(n_309),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_82),
.Y(n_283)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_85),
.Y(n_194)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_85),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g284 ( 
.A(n_85),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_85),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_86),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g365 ( 
.A(n_87),
.Y(n_365)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_87),
.Y(n_429)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_90),
.A2(n_309),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_91),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g374 ( 
.A(n_95),
.B(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_123),
.B1(n_131),
.B2(n_132),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_131),
.B1(n_132),
.B2(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_101),
.A2(n_131),
.B1(n_176),
.B2(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_101),
.A2(n_131),
.B1(n_388),
.B2(n_442),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_106),
.B1(n_110),
.B2(n_115),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_104),
.Y(n_373)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_105),
.Y(n_377)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_109),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_116),
.A2(n_124),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g469 ( 
.A1(n_116),
.A2(n_174),
.B1(n_392),
.B2(n_470),
.Y(n_469)
);

AO22x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_122),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_130),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_130),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_131),
.B(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_131),
.A2(n_388),
.B(n_391),
.Y(n_387)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_152),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_181),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g218 ( 
.A(n_160),
.B(n_163),
.CI(n_181),
.CON(n_218),
.SN(n_218)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_163),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_173),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI32xp33_ASAP7_75t_L g370 ( 
.A1(n_169),
.A2(n_250),
.A3(n_355),
.B1(n_371),
.B2(n_374),
.Y(n_370)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_171),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_174),
.A2(n_353),
.B(n_358),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_174),
.B(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_174),
.A2(n_358),
.B(n_486),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_SL g353 ( 
.A1(n_178),
.A2(n_273),
.B(n_354),
.Y(n_353)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B(n_205),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_199),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_205),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_183),
.A2(n_199),
.B1(n_224),
.B2(n_457),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_190),
.B(n_193),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_184),
.A2(n_193),
.B1(n_231),
.B2(n_235),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_184),
.A2(n_287),
.B(n_295),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_184),
.A2(n_273),
.B(n_295),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_184),
.A2(n_235),
.B1(n_423),
.B2(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_185),
.B(n_296),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_185),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_185),
.A2(n_363),
.B1(n_396),
.B2(n_400),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_185),
.A2(n_425),
.B1(n_463),
.B2(n_464),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_192),
.Y(n_464)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_197),
.Y(n_294)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_197),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_198),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_199),
.Y(n_457)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_210),
.B(n_273),
.Y(n_420)
);

OAI21xp33_ASAP7_75t_SL g438 ( 
.A1(n_210),
.A2(n_273),
.B(n_420),
.Y(n_438)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_259),
.B(n_512),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_218),
.B(n_219),
.Y(n_512)
);

BUFx24_ASAP7_75t_SL g521 ( 
.A(n_218),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.C(n_228),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_225),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_228),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_244),
.C(n_252),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_229),
.B(n_455),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_230),
.B(n_238),
.Y(n_480)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_231),
.Y(n_463)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_233),
.Y(n_398)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_233),
.Y(n_431)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_236),
.B(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_239),
.Y(n_461)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_244),
.B(n_252),
.Y(n_455)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_245),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_247),
.Y(n_246)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_258),
.Y(n_439)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI311xp33_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_451),
.A3(n_488),
.B1(n_506),
.C1(n_511),
.Y(n_261)
);

AOI21x1_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_404),
.B(n_450),
.Y(n_262)
);

AO21x1_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_379),
.B(n_403),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_339),
.B(n_378),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_312),
.B(n_338),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_285),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_267),
.B(n_285),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_268),
.A2(n_278),
.B1(n_279),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_268),
.Y(n_336)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx11_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_302),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_303),
.C(n_311),
.Y(n_340)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_292),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_310),
.B2(n_311),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_328),
.B(n_337),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_321),
.B(n_327),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_326),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_324),
.B(n_325),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_325),
.A2(n_362),
.B(n_367),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_335),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_335),
.Y(n_337)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_341),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_360),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_351),
.B2(n_352),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_344),
.B(n_351),
.C(n_360),
.Y(n_380)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx5_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx6_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_359),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_370),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_370),
.Y(n_385)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_380),
.B(n_381),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_386),
.B2(n_402),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_385),
.C(n_402),
.Y(n_405)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_386),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_393),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_387),
.B(n_394),
.C(n_395),
.Y(n_432)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_405),
.B(n_406),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_435),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_432),
.B1(n_433),
.B2(n_434),
.Y(n_407)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_421),
.B2(n_422),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_410),
.B(n_421),
.Y(n_484)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_432),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_432),
.B(n_433),
.C(n_435),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_440),
.B2(n_449),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_436),
.B(n_441),
.C(n_445),
.Y(n_497)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_440),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_445),
.Y(n_440)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_442),
.Y(n_486)
);

INVx6_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_474),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_452),
.A2(n_474),
.B(n_507),
.C(n_510),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_471),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_453),
.B(n_471),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.C(n_458),
.Y(n_453)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_454),
.B(n_456),
.CI(n_458),
.CON(n_487),
.SN(n_487)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_465),
.C(n_469),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_462),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_462),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_465),
.A2(n_466),
.B1(n_469),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_469),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_487),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.C(n_481),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.C(n_485),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_482),
.A2(n_483),
.B1(n_485),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g520 ( 
.A(n_487),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_501),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_498),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_498),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.C(n_497),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_504),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_496),
.B1(n_497),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_497),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_503),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_514),
.Y(n_517)
);

INVx13_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);


endmodule