module fake_jpeg_30891_n_405 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_405);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_405;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_51),
.Y(n_92)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_49),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_0),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_40),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_53),
.B(n_65),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_58),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_68),
.Y(n_110)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx2_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_71),
.B(n_82),
.Y(n_117)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_88),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx11_ASAP7_75t_SL g83 ( 
.A(n_40),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_84),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_86),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_24),
.Y(n_124)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_36),
.B1(n_28),
.B2(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_90),
.A2(n_128),
.B1(n_133),
.B2(n_24),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_43),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_25),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_22),
.B1(n_20),
.B2(n_41),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_54),
.A2(n_41),
.B1(n_16),
.B2(n_17),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_119),
.A2(n_138),
.B1(n_139),
.B2(n_7),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_124),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_60),
.A2(n_28),
.B1(n_34),
.B2(n_26),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_71),
.B(n_24),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_56),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_61),
.A2(n_34),
.B1(n_41),
.B2(n_27),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_27),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_100),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_27),
.B1(n_23),
.B2(n_17),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_75),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_23),
.B1(n_16),
.B2(n_15),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_140),
.A2(n_15),
.B1(n_79),
.B2(n_74),
.Y(n_142)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_109),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_141),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_150),
.B1(n_156),
.B2(n_108),
.Y(n_200)
);

BUFx4f_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_143),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_103),
.B(n_15),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_144),
.B(n_157),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_148),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_56),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_155),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_104),
.A2(n_63),
.B1(n_52),
.B2(n_49),
.Y(n_150)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

OA22x2_ASAP7_75t_SL g153 ( 
.A1(n_112),
.A2(n_83),
.B1(n_48),
.B2(n_46),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

OA22x2_ASAP7_75t_SL g154 ( 
.A1(n_112),
.A2(n_84),
.B1(n_85),
.B2(n_87),
.Y(n_154)
);

AO22x1_ASAP7_75t_SL g205 ( 
.A1(n_154),
.A2(n_161),
.B1(n_166),
.B2(n_178),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_57),
.B1(n_64),
.B2(n_78),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_98),
.B(n_84),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_99),
.B(n_24),
.C(n_2),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_165),
.C(n_167),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_111),
.A2(n_24),
.B1(n_2),
.B2(n_4),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_179),
.B1(n_108),
.B2(n_126),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g165 ( 
.A(n_91),
.B(n_1),
.Y(n_165)
);

AOI22x1_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_139),
.A2(n_132),
.B1(n_125),
.B2(n_101),
.Y(n_167)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_123),
.Y(n_169)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_5),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_177),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_121),
.B(n_5),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_7),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_89),
.A2(n_118),
.B(n_114),
.C(n_127),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_100),
.B(n_7),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_11),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_117),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_183),
.Y(n_213)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_102),
.Y(n_182)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_109),
.B(n_8),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_137),
.Y(n_184)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_101),
.B(n_8),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_185),
.B(n_11),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_89),
.B(n_8),
.C(n_9),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_102),
.C(n_129),
.Y(n_199)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_137),
.B1(n_118),
.B2(n_120),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_210),
.B1(n_221),
.B2(n_157),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_209),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_166),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_142),
.A2(n_156),
.B1(n_155),
.B2(n_149),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_203),
.A2(n_204),
.B1(n_211),
.B2(n_218),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_150),
.A2(n_134),
.B1(n_120),
.B2(n_113),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_215),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_129),
.C(n_115),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_217),
.C(n_165),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_179),
.A2(n_134),
.B1(n_113),
.B2(n_97),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_115),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_212),
.B(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_107),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_180),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_126),
.B1(n_131),
.B2(n_14),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_170),
.A2(n_146),
.B1(n_154),
.B2(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_228),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_154),
.B(n_153),
.Y(n_227)
);

AOI221xp5_ASAP7_75t_L g267 ( 
.A1(n_227),
.A2(n_237),
.B1(n_206),
.B2(n_209),
.C(n_199),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_193),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_222),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_232),
.B(n_246),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_252),
.Y(n_277)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_188),
.A2(n_175),
.B(n_185),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_193),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_239),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_225),
.B1(n_223),
.B2(n_212),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_240),
.A2(n_242),
.B1(n_243),
.B2(n_250),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_224),
.A2(n_181),
.B1(n_141),
.B2(n_153),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_241),
.A2(n_255),
.B(n_191),
.C(n_224),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_146),
.B1(n_164),
.B2(n_172),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_201),
.B(n_174),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_245),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_165),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_216),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_248),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_152),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_166),
.B1(n_161),
.B2(n_158),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_161),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_254),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_210),
.A2(n_163),
.B1(n_143),
.B2(n_160),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_169),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_205),
.A2(n_184),
.B1(n_159),
.B2(n_143),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_189),
.A2(n_186),
.B(n_182),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_202),
.B(n_219),
.Y(n_278)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_214),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_205),
.A2(n_131),
.B1(n_168),
.B2(n_176),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_258),
.A2(n_234),
.B1(n_252),
.B2(n_241),
.Y(n_263)
);

NOR2x1_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_205),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_260),
.A2(n_281),
.B(n_282),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_217),
.C(n_196),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_274),
.C(n_242),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_263),
.A2(n_265),
.B1(n_280),
.B2(n_255),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_189),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_238),
.C(n_256),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_233),
.A2(n_191),
.B1(n_190),
.B2(n_219),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_266),
.A2(n_278),
.B(n_279),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_267),
.B(n_238),
.Y(n_307)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_208),
.B(n_202),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_234),
.A2(n_190),
.B1(n_195),
.B2(n_214),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_233),
.A2(n_208),
.B(n_190),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_251),
.A2(n_195),
.B(n_177),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_249),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_287),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_243),
.A2(n_195),
.B(n_13),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_245),
.B(n_243),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_254),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_258),
.B1(n_247),
.B2(n_240),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_304),
.B1(n_280),
.B2(n_260),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_291),
.A2(n_305),
.B1(n_309),
.B2(n_265),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_298),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_278),
.B(n_270),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_294),
.A2(n_310),
.B(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_303),
.C(n_312),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_235),
.Y(n_298)
);

XOR2x1_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_237),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_300),
.B(n_307),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_259),
.B(n_235),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_308),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_257),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_302),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_274),
.C(n_262),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_284),
.A2(n_258),
.B1(n_286),
.B2(n_263),
.Y(n_304)
);

HAxp5_ASAP7_75t_SL g305 ( 
.A(n_259),
.B(n_244),
.CON(n_305),
.SN(n_305)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_261),
.B(n_250),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_277),
.A2(n_243),
.B1(n_229),
.B2(n_242),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_270),
.A2(n_248),
.B(n_236),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_271),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_283),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_277),
.B(n_265),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_290),
.Y(n_346)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_298),
.Y(n_315)
);

INVx13_ASAP7_75t_L g338 ( 
.A(n_315),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_316),
.A2(n_304),
.B1(n_314),
.B2(n_288),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_317),
.A2(n_309),
.B1(n_299),
.B2(n_306),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_268),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_329),
.C(n_331),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_268),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_333),
.C(n_289),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_324),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_273),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_276),
.C(n_272),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_269),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_334),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_307),
.B(n_272),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_299),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_321),
.Y(n_359)
);

AOI322xp5_ASAP7_75t_L g340 ( 
.A1(n_313),
.A2(n_319),
.A3(n_294),
.B1(n_290),
.B2(n_334),
.C1(n_315),
.C2(n_317),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_340),
.A2(n_351),
.B1(n_292),
.B2(n_300),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_341),
.A2(n_344),
.B1(n_347),
.B2(n_276),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_332),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_350),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_323),
.A2(n_292),
.B1(n_295),
.B2(n_291),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g357 ( 
.A(n_346),
.B(n_318),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_330),
.Y(n_348)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_348),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_301),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_349),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_261),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_326),
.B(n_310),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_269),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_352),
.B(n_320),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_353),
.B(n_354),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_321),
.C(n_339),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_SL g356 ( 
.A1(n_346),
.A2(n_265),
.B(n_318),
.C(n_281),
.Y(n_356)
);

AO21x1_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_357),
.B(n_335),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_365),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_322),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_360),
.B(n_363),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_361),
.A2(n_364),
.B1(n_336),
.B2(n_342),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_341),
.A2(n_265),
.B1(n_300),
.B2(n_325),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_333),
.C(n_325),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_351),
.Y(n_372)
);

OA21x2_ASAP7_75t_SL g367 ( 
.A1(n_362),
.A2(n_349),
.B(n_348),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_367),
.A2(n_345),
.B(n_344),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_369),
.B(n_375),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_355),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_370),
.B(n_371),
.Y(n_381)
);

AOI322xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_338),
.A3(n_350),
.B1(n_343),
.B2(n_345),
.C1(n_342),
.C2(n_336),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_354),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_347),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_361),
.C(n_366),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_374),
.A2(n_375),
.B1(n_356),
.B2(n_377),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_357),
.A2(n_335),
.B(n_340),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_378),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_380),
.B(n_376),
.C(n_365),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_373),
.A2(n_356),
.B1(n_229),
.B2(n_338),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_383),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_369),
.B(n_338),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_386),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_374),
.A2(n_356),
.B(n_311),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_385),
.A2(n_296),
.B(n_368),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_387),
.B(n_391),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_388),
.Y(n_396)
);

FAx1_ASAP7_75t_SL g390 ( 
.A(n_385),
.B(n_377),
.CI(n_376),
.CON(n_390),
.SN(n_390)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_390),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_379),
.A2(n_359),
.B(n_360),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_381),
.B1(n_392),
.B2(n_389),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_395),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_389),
.A2(n_379),
.B1(n_383),
.B2(n_382),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_397),
.B(n_380),
.C(n_390),
.Y(n_399)
);

AOI321xp33_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_12),
.A3(n_13),
.B1(n_396),
.B2(n_397),
.C(n_387),
.Y(n_403)
);

AOI211xp5_ASAP7_75t_L g400 ( 
.A1(n_398),
.A2(n_283),
.B(n_239),
.C(n_228),
.Y(n_400)
);

OAI321xp33_ASAP7_75t_L g402 ( 
.A1(n_400),
.A2(n_396),
.A3(n_232),
.B1(n_246),
.B2(n_13),
.C(n_14),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_403),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_404),
.B(n_401),
.Y(n_405)
);


endmodule