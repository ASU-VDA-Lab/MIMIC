module fake_netlist_1_8170_n_781 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_781);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_781;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_466;
wire n_302;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_59), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_39), .Y(n_95) );
BUFx10_ASAP7_75t_L g96 ( .A(n_39), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_20), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_33), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_22), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_9), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_50), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_79), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_76), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_2), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_67), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_78), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_84), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_53), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_47), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_69), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_80), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_42), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_30), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_49), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_5), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_82), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_66), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_87), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_90), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_83), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_9), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_57), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_60), .Y(n_126) );
BUFx10_ASAP7_75t_L g127 ( .A(n_41), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_6), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_33), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_10), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_15), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_24), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_31), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_10), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_55), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_65), .Y(n_137) );
XNOR2xp5_ASAP7_75t_L g138 ( .A(n_117), .B(n_0), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_123), .Y(n_139) );
INVx5_ASAP7_75t_L g140 ( .A(n_103), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_95), .B(n_93), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_95), .B(n_43), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_114), .B(n_0), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_114), .B(n_1), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_106), .B(n_1), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_127), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_103), .B(n_95), .Y(n_147) );
INVx5_ASAP7_75t_L g148 ( .A(n_103), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_99), .B(n_2), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_106), .B(n_96), .Y(n_150) );
BUFx12f_ASAP7_75t_L g151 ( .A(n_127), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_105), .B(n_3), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_105), .B(n_3), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_96), .B(n_4), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_116), .B(n_4), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_99), .B(n_5), .Y(n_158) );
BUFx3_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_109), .B(n_6), .Y(n_160) );
INVx5_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
OAI22xp33_ASAP7_75t_SL g163 ( .A1(n_143), .A2(n_131), .B1(n_97), .B2(n_135), .Y(n_163) );
OAI22xp33_ASAP7_75t_L g164 ( .A1(n_143), .A2(n_117), .B1(n_129), .B2(n_115), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_147), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_150), .B(n_96), .Y(n_167) );
OAI22xp33_ASAP7_75t_L g168 ( .A1(n_143), .A2(n_129), .B1(n_128), .B2(n_115), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_150), .B(n_96), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_138), .A2(n_109), .B1(n_128), .B2(n_124), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_150), .B(n_96), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_150), .A2(n_130), .B1(n_98), .B2(n_134), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g173 ( .A1(n_144), .A2(n_124), .B1(n_100), .B2(n_133), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_144), .A2(n_104), .B1(n_116), .B2(n_120), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_144), .B(n_123), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_147), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
AO22x2_ASAP7_75t_L g178 ( .A1(n_155), .A2(n_118), .B1(n_120), .B2(n_119), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_152), .B(n_118), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_155), .A2(n_111), .B1(n_137), .B2(n_113), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_152), .B(n_127), .Y(n_182) );
BUFx6f_ASAP7_75t_SL g183 ( .A(n_152), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_152), .B(n_125), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_155), .A2(n_125), .B1(n_132), .B2(n_127), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_155), .A2(n_125), .B1(n_132), .B2(n_11), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_149), .A2(n_136), .B1(n_126), .B2(n_122), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g189 ( .A1(n_145), .A2(n_121), .B1(n_112), .B2(n_110), .Y(n_189) );
BUFx10_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
BUFx2_ASAP7_75t_L g191 ( .A(n_151), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_152), .B(n_94), .Y(n_192) );
OAI22xp33_ASAP7_75t_SL g193 ( .A1(n_149), .A2(n_108), .B1(n_107), .B2(n_102), .Y(n_193) );
AO22x2_ASAP7_75t_L g194 ( .A1(n_145), .A2(n_7), .B1(n_8), .B2(n_11), .Y(n_194) );
OA22x2_ASAP7_75t_L g195 ( .A1(n_147), .A2(n_101), .B1(n_8), .B2(n_12), .Y(n_195) );
OAI22xp33_ASAP7_75t_SL g196 ( .A1(n_158), .A2(n_7), .B1(n_12), .B2(n_13), .Y(n_196) );
AO22x2_ASAP7_75t_L g197 ( .A1(n_145), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_145), .A2(n_14), .B1(n_16), .B2(n_17), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_151), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_152), .A2(n_18), .B1(n_19), .B2(n_20), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_151), .A2(n_19), .B1(n_21), .B2(n_23), .Y(n_201) );
OAI22xp33_ASAP7_75t_L g202 ( .A1(n_158), .A2(n_21), .B1(n_23), .B2(n_24), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
BUFx6f_ASAP7_75t_SL g204 ( .A(n_141), .Y(n_204) );
AOI22xp5_ASAP7_75t_SL g205 ( .A1(n_138), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_151), .A2(n_25), .B1(n_26), .B2(n_27), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_190), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_190), .Y(n_208) );
XOR2xp5_ASAP7_75t_L g209 ( .A(n_170), .B(n_138), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_203), .B(n_151), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_178), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_178), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_191), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_166), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_167), .B(n_146), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_176), .Y(n_217) );
XOR2xp5_ASAP7_75t_L g218 ( .A(n_170), .B(n_138), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_177), .B(n_146), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_169), .B(n_146), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_187), .B(n_146), .Y(n_221) );
AND2x6_ASAP7_75t_L g222 ( .A(n_171), .B(n_146), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_180), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_175), .B(n_146), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_185), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_179), .A2(n_146), .B(n_148), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_162), .B(n_140), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_188), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_186), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_165), .B(n_160), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_186), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_184), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_195), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_195), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_182), .B(n_160), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_173), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_173), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_172), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_192), .B(n_148), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_199), .Y(n_245) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_168), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_189), .B(n_156), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_193), .B(n_156), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_164), .B(n_153), .Y(n_249) );
NAND2x1p5_ASAP7_75t_L g250 ( .A(n_201), .B(n_148), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_206), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_183), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_205), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_181), .B(n_154), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_194), .Y(n_255) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_174), .A2(n_148), .B(n_140), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_163), .B(n_154), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_194), .B(n_153), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_183), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_194), .B(n_159), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_197), .Y(n_261) );
XOR2xp5_ASAP7_75t_L g262 ( .A(n_164), .B(n_28), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_197), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_168), .B(n_174), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
INVxp33_ASAP7_75t_SL g266 ( .A(n_200), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_200), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_200), .Y(n_268) );
OR2x2_ASAP7_75t_L g269 ( .A(n_187), .B(n_139), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_254), .B(n_204), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_232), .B(n_139), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_219), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_232), .B(n_139), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_210), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_210), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_239), .B(n_139), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_239), .B(n_159), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_230), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_239), .B(n_140), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_219), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_215), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_264), .B(n_159), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_217), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_264), .B(n_159), .Y(n_287) );
INVx3_ASAP7_75t_SL g288 ( .A(n_259), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_223), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_258), .B(n_159), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_235), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_240), .B(n_148), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_213), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_216), .B(n_140), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_235), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_254), .B(n_204), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_236), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_258), .B(n_140), .Y(n_299) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_259), .B(n_141), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_236), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_241), .B(n_148), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_216), .B(n_140), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_220), .B(n_140), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_220), .B(n_140), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_211), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_254), .B(n_148), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_212), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_246), .B(n_148), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_259), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_213), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_214), .Y(n_313) );
NOR2xp33_ASAP7_75t_SL g314 ( .A(n_266), .B(n_141), .Y(n_314) );
AND2x2_ASAP7_75t_SL g315 ( .A(n_260), .B(n_141), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_225), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_231), .B(n_148), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_225), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_207), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_222), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_207), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_242), .B(n_140), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_140), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_275), .B(n_237), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_271), .Y(n_325) );
NOR2x1_ASAP7_75t_R g326 ( .A(n_307), .B(n_253), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_275), .B(n_251), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_288), .Y(n_328) );
AND2x6_ASAP7_75t_L g329 ( .A(n_283), .B(n_231), .Y(n_329) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_273), .B(n_226), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g331 ( .A(n_273), .B(n_226), .Y(n_331) );
NAND2x1_ASAP7_75t_SL g332 ( .A(n_288), .B(n_267), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_273), .Y(n_333) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_273), .B(n_227), .Y(n_334) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_283), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
BUFx4f_ASAP7_75t_L g338 ( .A(n_283), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_271), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_273), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_273), .B(n_208), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_275), .B(n_237), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_280), .Y(n_344) );
AND2x2_ASAP7_75t_SL g345 ( .A(n_314), .B(n_233), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_280), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_293), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_280), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_276), .B(n_209), .Y(n_349) );
INVx6_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
NOR2xp33_ASAP7_75t_SL g351 ( .A(n_314), .B(n_266), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_281), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_288), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_288), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_281), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_276), .B(n_238), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_273), .B(n_227), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_335), .B(n_307), .Y(n_358) );
INVx5_ASAP7_75t_L g359 ( .A(n_333), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_335), .B(n_307), .Y(n_360) );
CKINVDCx11_ASAP7_75t_R g361 ( .A(n_328), .Y(n_361) );
BUFx2_ASAP7_75t_SL g362 ( .A(n_353), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_335), .Y(n_363) );
INVx5_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_336), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_333), .Y(n_366) );
BUFx3_ASAP7_75t_L g367 ( .A(n_335), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_349), .B(n_253), .Y(n_368) );
BUFx4f_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_336), .Y(n_370) );
INVx4_ASAP7_75t_L g371 ( .A(n_338), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_336), .Y(n_372) );
BUFx8_ASAP7_75t_L g373 ( .A(n_353), .Y(n_373) );
BUFx2_ASAP7_75t_SL g374 ( .A(n_353), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_338), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_338), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_336), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_341), .Y(n_379) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_338), .Y(n_381) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
INVx6_ASAP7_75t_SL g383 ( .A(n_342), .Y(n_383) );
BUFx3_ASAP7_75t_L g384 ( .A(n_350), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_341), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_336), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_368), .B(n_327), .Y(n_388) );
BUFx8_ASAP7_75t_L g389 ( .A(n_382), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_382), .Y(n_390) );
INVx6_ASAP7_75t_L g391 ( .A(n_382), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_379), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_369), .A2(n_351), .B1(n_349), .B2(n_371), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_379), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_385), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_382), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_385), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_369), .A2(n_209), .B1(n_218), .B2(n_345), .Y(n_399) );
BUFx12f_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
OAI22xp33_ASAP7_75t_SL g401 ( .A1(n_358), .A2(n_261), .B1(n_265), .B2(n_263), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_369), .A2(n_262), .B1(n_248), .B2(n_257), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_385), .Y(n_403) );
CKINVDCx11_ASAP7_75t_R g404 ( .A(n_361), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_373), .Y(n_405) );
BUFx8_ASAP7_75t_L g406 ( .A(n_382), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_369), .A2(n_218), .B1(n_255), .B2(n_345), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_369), .A2(n_314), .B1(n_276), .B2(n_327), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_369), .A2(n_341), .B1(n_267), .B2(n_268), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_371), .A2(n_268), .B1(n_233), .B2(n_234), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_387), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_373), .A2(n_250), .B1(n_315), .B2(n_270), .Y(n_414) );
AOI21xp5_ASAP7_75t_SL g415 ( .A1(n_371), .A2(n_367), .B(n_363), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_373), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_383), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_373), .A2(n_250), .B1(n_315), .B2(n_270), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_373), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_371), .A2(n_350), .B1(n_325), .B2(n_344), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_373), .A2(n_315), .B1(n_270), .B2(n_297), .Y(n_421) );
CKINVDCx11_ASAP7_75t_R g422 ( .A(n_363), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_366), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_383), .A2(n_315), .B1(n_297), .B2(n_249), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_366), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_371), .A2(n_350), .B1(n_325), .B2(n_346), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_371), .A2(n_350), .B1(n_339), .B2(n_346), .Y(n_428) );
BUFx10_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_399), .A2(n_383), .B1(n_315), .B2(n_367), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_402), .A2(n_383), .B1(n_363), .B2(n_367), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_389), .A2(n_383), .B1(n_363), .B2(n_367), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
INVx8_ASAP7_75t_L g434 ( .A(n_405), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_397), .A2(n_360), .B(n_358), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_388), .A2(n_297), .B1(n_375), .B2(n_377), .Y(n_436) );
OAI21xp33_ASAP7_75t_L g437 ( .A1(n_408), .A2(n_196), .B(n_260), .Y(n_437) );
OAI222xp33_ASAP7_75t_L g438 ( .A1(n_397), .A2(n_364), .B1(n_359), .B2(n_360), .C1(n_358), .C2(n_376), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_389), .A2(n_383), .B1(n_377), .B2(n_381), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_389), .A2(n_377), .B1(n_375), .B2(n_381), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_406), .A2(n_394), .B1(n_391), .B2(n_425), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_391), .A2(n_375), .B1(n_359), .B2(n_364), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_406), .A2(n_375), .B1(n_364), .B2(n_359), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_404), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_390), .B(n_359), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_414), .A2(n_360), .B(n_358), .Y(n_447) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_429), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_393), .B(n_238), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_406), .A2(n_359), .B1(n_364), .B2(n_290), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_429), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_359), .B1(n_364), .B2(n_290), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_390), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_352), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_395), .B(n_352), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g458 ( .A1(n_418), .A2(n_360), .B(n_358), .Y(n_458) );
INVx2_ASAP7_75t_SL g459 ( .A(n_416), .Y(n_459) );
INVx5_ASAP7_75t_SL g460 ( .A(n_416), .Y(n_460) );
BUFx4f_ASAP7_75t_SL g461 ( .A(n_400), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_396), .B(n_352), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_429), .Y(n_463) );
AOI22xp33_ASAP7_75t_SL g464 ( .A1(n_419), .A2(n_362), .B1(n_374), .B2(n_364), .Y(n_464) );
INVx6_ASAP7_75t_L g465 ( .A(n_400), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_422), .A2(n_364), .B1(n_359), .B2(n_329), .Y(n_466) );
INVx4_ASAP7_75t_SL g467 ( .A(n_403), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_417), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_401), .B(n_324), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_407), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_421), .A2(n_364), .B1(n_359), .B2(n_360), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_420), .A2(n_359), .B1(n_364), .B2(n_358), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_423), .Y(n_474) );
INVx5_ASAP7_75t_SL g475 ( .A(n_415), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_410), .A2(n_360), .B1(n_376), .B2(n_366), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_409), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_409), .B(n_355), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_424), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_424), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_415), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_427), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_426), .B(n_355), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_426), .Y(n_484) );
OAI21xp5_ASAP7_75t_SL g485 ( .A1(n_428), .A2(n_202), .B(n_326), .Y(n_485) );
OAI222xp33_ASAP7_75t_L g486 ( .A1(n_411), .A2(n_366), .B1(n_376), .B2(n_326), .C1(n_354), .C2(n_328), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_412), .B(n_243), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_398), .B(n_355), .Y(n_488) );
INVx5_ASAP7_75t_SL g489 ( .A(n_389), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_388), .B(n_339), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_397), .Y(n_491) );
OAI21xp5_ASAP7_75t_SL g492 ( .A1(n_435), .A2(n_376), .B(n_366), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_441), .A2(n_374), .B1(n_362), .B2(n_376), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_430), .A2(n_386), .B1(n_384), .B2(n_350), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_482), .A2(n_386), .B1(n_384), .B2(n_362), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_482), .A2(n_386), .B1(n_384), .B2(n_374), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_437), .A2(n_329), .B1(n_376), .B2(n_285), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_487), .A2(n_329), .B1(n_287), .B2(n_285), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_485), .A2(n_247), .B1(n_332), .B2(n_340), .C(n_269), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_489), .A2(n_340), .B1(n_344), .B2(n_348), .Y(n_501) );
OAI222xp33_ASAP7_75t_L g502 ( .A1(n_481), .A2(n_378), .B1(n_370), .B2(n_365), .C1(n_354), .C2(n_340), .Y(n_502) );
OAI21xp5_ASAP7_75t_SL g503 ( .A1(n_438), .A2(n_300), .B(n_287), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_443), .B(n_387), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_431), .A2(n_329), .B1(n_285), .B2(n_287), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_434), .A2(n_340), .B1(n_142), .B2(n_141), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_491), .B(n_247), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_434), .A2(n_142), .B1(n_141), .B2(n_342), .Y(n_508) );
INVxp67_ASAP7_75t_SL g509 ( .A(n_474), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_453), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_434), .A2(n_142), .B1(n_141), .B2(n_342), .Y(n_511) );
OAI222xp33_ASAP7_75t_L g512 ( .A1(n_481), .A2(n_378), .B1(n_370), .B2(n_365), .C1(n_334), .C2(n_357), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_459), .A2(n_142), .B1(n_141), .B2(n_342), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_447), .A2(n_284), .B1(n_286), .B2(n_289), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_470), .A2(n_141), .B1(n_142), .B2(n_300), .Y(n_515) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_458), .A2(n_357), .B1(n_331), .B2(n_330), .Y(n_516) );
OAI222xp33_ASAP7_75t_L g517 ( .A1(n_446), .A2(n_378), .B1(n_370), .B2(n_365), .C1(n_334), .C2(n_357), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g518 ( .A1(n_489), .A2(n_307), .B1(n_372), .B2(n_380), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_472), .A2(n_141), .B1(n_142), .B2(n_299), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_457), .B(n_387), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_444), .A2(n_330), .B1(n_331), .B2(n_334), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g522 ( .A1(n_442), .A2(n_330), .B1(n_331), .B2(n_387), .C1(n_307), .C2(n_269), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_455), .B(n_372), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_466), .A2(n_330), .B1(n_356), .B2(n_343), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_464), .A2(n_356), .B1(n_343), .B2(n_372), .Y(n_525) );
AOI222xp33_ASAP7_75t_L g526 ( .A1(n_461), .A2(n_142), .B1(n_284), .B2(n_313), .C1(n_309), .C2(n_306), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_489), .A2(n_316), .B1(n_318), .B2(n_313), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_450), .A2(n_316), .B1(n_318), .B2(n_306), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_457), .B(n_332), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_467), .B(n_372), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_456), .B(n_372), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_436), .A2(n_323), .B1(n_322), .B2(n_308), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_468), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_475), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_452), .A2(n_316), .B1(n_318), .B2(n_306), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_453), .A2(n_313), .B1(n_309), .B2(n_323), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_465), .A2(n_323), .B1(n_322), .B2(n_308), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_432), .A2(n_320), .B1(n_308), .B2(n_372), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_439), .A2(n_320), .B1(n_372), .B2(n_380), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_440), .A2(n_372), .B1(n_380), .B2(n_321), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_476), .A2(n_309), .B1(n_322), .B2(n_295), .Y(n_541) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_486), .A2(n_490), .B(n_454), .Y(n_542) );
OAI21xp5_ASAP7_75t_SL g543 ( .A1(n_473), .A2(n_256), .B(n_277), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_465), .A2(n_293), .B1(n_295), .B2(n_312), .Y(n_544) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_465), .A2(n_288), .B1(n_372), .B2(n_380), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_475), .A2(n_380), .B1(n_347), .B2(n_337), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_465), .A2(n_295), .B1(n_312), .B2(n_293), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_479), .A2(n_295), .B1(n_312), .B2(n_293), .Y(n_548) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_460), .A2(n_380), .B1(n_278), .B2(n_311), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_484), .A2(n_295), .B1(n_312), .B2(n_293), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_484), .A2(n_295), .B1(n_312), .B2(n_293), .Y(n_551) );
OAI222xp33_ASAP7_75t_L g552 ( .A1(n_469), .A2(n_161), .B1(n_281), .B2(n_221), .C1(n_321), .C2(n_274), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_460), .A2(n_295), .B1(n_312), .B2(n_293), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_460), .A2(n_295), .B1(n_293), .B2(n_312), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_488), .B(n_29), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_471), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_477), .B(n_161), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_448), .A2(n_278), .B1(n_311), .B2(n_336), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_480), .A2(n_295), .B1(n_312), .B2(n_278), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_478), .A2(n_281), .B1(n_291), .B2(n_298), .Y(n_560) );
OAI222xp33_ASAP7_75t_L g561 ( .A1(n_462), .A2(n_161), .B1(n_321), .B2(n_274), .C1(n_272), .C2(n_279), .Y(n_561) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_451), .A2(n_347), .B1(n_337), .B2(n_274), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_483), .A2(n_291), .B1(n_321), .B2(n_274), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_451), .A2(n_317), .B1(n_222), .B2(n_296), .Y(n_564) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_514), .A2(n_463), .B(n_451), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_509), .B(n_467), .Y(n_566) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_542), .A2(n_449), .B(n_483), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_510), .B(n_514), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_503), .A2(n_463), .B1(n_451), .B2(n_454), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_516), .B(n_451), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_496), .B(n_463), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_507), .B(n_463), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_500), .B(n_463), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_492), .B(n_445), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_510), .B(n_467), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_492), .B(n_445), .Y(n_576) );
AOI221xp5_ASAP7_75t_L g577 ( .A1(n_542), .A2(n_161), .B1(n_272), .B2(n_277), .C(n_279), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_518), .B(n_337), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_503), .A2(n_288), .B1(n_337), .B2(n_347), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g580 ( .A(n_534), .B(n_337), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_533), .Y(n_581) );
AND2x2_ASAP7_75t_SL g582 ( .A(n_530), .B(n_534), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_521), .A2(n_347), .B1(n_337), .B2(n_272), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g584 ( .A1(n_512), .A2(n_277), .B(n_279), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_556), .B(n_32), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_529), .B(n_32), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_526), .B(n_161), .C(n_292), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_555), .B(n_34), .Y(n_588) );
OAI221xp5_ASAP7_75t_SL g589 ( .A1(n_499), .A2(n_310), .B1(n_292), .B2(n_302), .C(n_296), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_495), .A2(n_319), .B1(n_296), .B2(n_301), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_504), .B(n_34), .Y(n_591) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_561), .B(n_310), .C(n_302), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_526), .B(n_161), .C(n_292), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_493), .B(n_35), .Y(n_594) );
OAI21xp33_ASAP7_75t_SL g595 ( .A1(n_497), .A2(n_310), .B(n_282), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_545), .B(n_213), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_508), .B(n_296), .C(n_301), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_520), .B(n_36), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_521), .A2(n_319), .B1(n_222), .B2(n_294), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g600 ( .A(n_511), .B(n_282), .C(n_38), .D(n_40), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_523), .B(n_37), .Y(n_601) );
NAND3xp33_ASAP7_75t_L g602 ( .A(n_506), .B(n_301), .C(n_213), .Y(n_602) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_552), .B(n_319), .C(n_301), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_523), .B(n_38), .Y(n_604) );
AND2x2_ASAP7_75t_SL g605 ( .A(n_530), .B(n_252), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_519), .B(n_319), .C(n_252), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_531), .B(n_40), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_493), .B(n_319), .C(n_294), .Y(n_608) );
OAI221xp5_ASAP7_75t_SL g609 ( .A1(n_498), .A2(n_305), .B1(n_304), .B2(n_319), .C(n_224), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_515), .B(n_303), .C(n_294), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_513), .B(n_303), .C(n_294), .Y(n_611) );
OAI221xp5_ASAP7_75t_SL g612 ( .A1(n_543), .A2(n_305), .B1(n_304), .B2(n_229), .C(n_208), .Y(n_612) );
OAI21xp5_ASAP7_75t_SL g613 ( .A1(n_522), .A2(n_303), .B(n_294), .Y(n_613) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_517), .A2(n_303), .B(n_294), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_501), .B(n_44), .Y(n_615) );
OAI21xp5_ASAP7_75t_SL g616 ( .A1(n_502), .A2(n_304), .B(n_46), .Y(n_616) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_534), .B(n_45), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_543), .A2(n_244), .B1(n_228), .B2(n_48), .C(n_51), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_530), .B(n_52), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_525), .A2(n_54), .B1(n_56), .B2(n_58), .C(n_61), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_537), .B(n_63), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_525), .A2(n_64), .B1(n_70), .B2(n_71), .C(n_72), .Y(n_622) );
OA21x2_ASAP7_75t_L g623 ( .A1(n_530), .A2(n_74), .B(n_75), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g624 ( .A1(n_524), .A2(n_222), .B1(n_77), .B2(n_81), .Y(n_624) );
NOR2xp33_ASAP7_75t_SL g625 ( .A(n_539), .B(n_524), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_505), .A2(n_222), .B1(n_86), .B2(n_88), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_562), .B(n_85), .Y(n_627) );
OAI21xp5_ASAP7_75t_SL g628 ( .A1(n_549), .A2(n_89), .B(n_91), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_537), .A2(n_92), .B1(n_532), .B2(n_536), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_563), .A2(n_560), .B(n_494), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g631 ( .A(n_557), .B(n_538), .C(n_540), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_563), .B(n_527), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_550), .B(n_551), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_541), .B(n_528), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_571), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_581), .B(n_546), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_594), .B(n_546), .C(n_558), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_565), .B(n_544), .C(n_547), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_574), .B(n_559), .C(n_548), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_594), .B(n_535), .C(n_564), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_574), .B(n_553), .C(n_554), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_582), .B(n_567), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_582), .B(n_567), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_601), .B(n_604), .Y(n_644) );
OA211x2_ASAP7_75t_L g645 ( .A1(n_576), .A2(n_570), .B(n_625), .C(n_578), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_607), .B(n_572), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_614), .A2(n_584), .B1(n_573), .B2(n_630), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_572), .B(n_573), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_566), .B(n_575), .Y(n_649) );
NAND4xp75_ASAP7_75t_L g650 ( .A(n_605), .B(n_577), .C(n_595), .D(n_568), .Y(n_650) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_629), .B(n_632), .C(n_612), .D(n_588), .Y(n_651) );
AND2x4_ASAP7_75t_L g652 ( .A(n_619), .B(n_631), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_583), .B(n_591), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_583), .B(n_586), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_633), .B(n_605), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_598), .B(n_585), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_580), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g658 ( .A1(n_579), .A2(n_608), .B1(n_632), .B2(n_623), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_599), .B(n_624), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_624), .B(n_599), .C(n_631), .Y(n_660) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_596), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_634), .A2(n_600), .B1(n_629), .B2(n_593), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_613), .A2(n_588), .B1(n_587), .B2(n_621), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_620), .B(n_622), .C(n_628), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_589), .B(n_609), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_617), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_592), .A2(n_610), .B1(n_611), .B2(n_603), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_615), .B(n_627), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_592), .B(n_603), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_590), .B(n_602), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_597), .B(n_606), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_626), .B(n_581), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_616), .B(n_594), .C(n_618), .Y(n_673) );
OAI211xp5_ASAP7_75t_SL g674 ( .A1(n_616), .A2(n_404), .B(n_576), .C(n_574), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_616), .B(n_594), .C(n_618), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_565), .B(n_616), .C(n_576), .Y(n_676) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_616), .B(n_594), .C(n_618), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_571), .B(n_509), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g679 ( .A(n_575), .B(n_481), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g680 ( .A1(n_574), .A2(n_576), .B1(n_605), .B2(n_569), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_565), .B(n_616), .C(n_576), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_632), .A2(n_574), .B1(n_576), .B2(n_577), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_565), .B(n_616), .C(n_576), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_565), .B(n_616), .C(n_576), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_565), .B(n_616), .C(n_576), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_616), .A2(n_565), .B(n_516), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_616), .B(n_594), .C(n_618), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_605), .B(n_516), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_635), .Y(n_689) );
NAND4xp75_ASAP7_75t_L g690 ( .A(n_645), .B(n_659), .C(n_686), .D(n_647), .Y(n_690) );
INVx1_ASAP7_75t_SL g691 ( .A(n_666), .Y(n_691) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_678), .Y(n_692) );
AO22x2_ASAP7_75t_L g693 ( .A1(n_642), .A2(n_643), .B1(n_652), .B2(n_681), .Y(n_693) );
NAND4xp75_ASAP7_75t_L g694 ( .A(n_659), .B(n_688), .C(n_669), .D(n_668), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_658), .B(n_660), .C(n_680), .Y(n_695) );
NAND4xp75_ASAP7_75t_L g696 ( .A(n_688), .B(n_665), .C(n_663), .D(n_654), .Y(n_696) );
INVx1_ASAP7_75t_SL g697 ( .A(n_666), .Y(n_697) );
INVx2_ASAP7_75t_SL g698 ( .A(n_649), .Y(n_698) );
XOR2x1_ASAP7_75t_L g699 ( .A(n_652), .B(n_649), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_636), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_676), .B(n_685), .C(n_684), .Y(n_701) );
INVx1_ASAP7_75t_SL g702 ( .A(n_666), .Y(n_702) );
INVxp67_ASAP7_75t_L g703 ( .A(n_648), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_648), .B(n_651), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_683), .B(n_664), .C(n_674), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_657), .Y(n_706) );
XNOR2x2_ASAP7_75t_L g707 ( .A(n_650), .B(n_638), .Y(n_707) );
XOR2x2_ASAP7_75t_L g708 ( .A(n_673), .B(n_687), .Y(n_708) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_675), .B(n_677), .C(n_667), .Y(n_709) );
BUFx2_ASAP7_75t_L g710 ( .A(n_679), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_667), .A2(n_661), .B1(n_682), .B2(n_655), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_646), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_644), .B(n_656), .Y(n_713) );
CKINVDCx8_ASAP7_75t_R g714 ( .A(n_679), .Y(n_714) );
XNOR2xp5_ASAP7_75t_L g715 ( .A(n_708), .B(n_662), .Y(n_715) );
BUFx3_ASAP7_75t_L g716 ( .A(n_706), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_689), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_692), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_704), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_706), .Y(n_720) );
INVx1_ASAP7_75t_SL g721 ( .A(n_691), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_697), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_700), .B(n_656), .Y(n_723) );
AO22x2_ASAP7_75t_L g724 ( .A1(n_694), .A2(n_641), .B1(n_672), .B2(n_653), .Y(n_724) );
OAI22x1_ASAP7_75t_L g725 ( .A1(n_709), .A2(n_653), .B1(n_672), .B2(n_639), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_700), .B(n_637), .Y(n_726) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_712), .Y(n_727) );
INVxp67_ASAP7_75t_L g728 ( .A(n_709), .Y(n_728) );
XNOR2x2_ASAP7_75t_L g729 ( .A(n_707), .B(n_671), .Y(n_729) );
XNOR2xp5_ASAP7_75t_L g730 ( .A(n_708), .B(n_662), .Y(n_730) );
XNOR2x1_ASAP7_75t_L g731 ( .A(n_696), .B(n_670), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_703), .B(n_682), .Y(n_732) );
INVx2_ASAP7_75t_SL g733 ( .A(n_698), .Y(n_733) );
XOR2x2_ASAP7_75t_L g734 ( .A(n_696), .B(n_640), .Y(n_734) );
XNOR2x1_ASAP7_75t_L g735 ( .A(n_707), .B(n_694), .Y(n_735) );
INVxp33_ASAP7_75t_L g736 ( .A(n_690), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_727), .Y(n_737) );
OA22x2_ASAP7_75t_L g738 ( .A1(n_725), .A2(n_702), .B1(n_711), .B2(n_710), .Y(n_738) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_720), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_716), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_716), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_718), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_735), .A2(n_705), .B1(n_695), .B2(n_701), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_733), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_717), .Y(n_745) );
XNOR2x1_ASAP7_75t_L g746 ( .A(n_715), .B(n_690), .Y(n_746) );
AOI22x1_ASAP7_75t_L g747 ( .A1(n_724), .A2(n_693), .B1(n_714), .B2(n_699), .Y(n_747) );
AOI22x1_ASAP7_75t_L g748 ( .A1(n_724), .A2(n_693), .B1(n_714), .B2(n_699), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_739), .Y(n_749) );
INVx2_ASAP7_75t_SL g750 ( .A(n_740), .Y(n_750) );
INVx2_ASAP7_75t_SL g751 ( .A(n_740), .Y(n_751) );
INVx1_ASAP7_75t_SL g752 ( .A(n_741), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_737), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_748), .A2(n_724), .B1(n_735), .B2(n_731), .Y(n_754) );
OA22x2_ASAP7_75t_L g755 ( .A1(n_743), .A2(n_728), .B1(n_730), .B2(n_719), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_737), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_742), .Y(n_757) );
OA22x2_ASAP7_75t_L g758 ( .A1(n_754), .A2(n_730), .B1(n_729), .B2(n_748), .Y(n_758) );
AND4x1_ASAP7_75t_L g759 ( .A(n_749), .B(n_736), .C(n_746), .D(n_729), .Y(n_759) );
AOI22x1_ASAP7_75t_L g760 ( .A1(n_752), .A2(n_724), .B1(n_746), .B2(n_736), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_754), .A2(n_734), .B1(n_731), .B2(n_738), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_752), .Y(n_762) );
INVxp67_ASAP7_75t_L g763 ( .A(n_762), .Y(n_763) );
INVx2_ASAP7_75t_SL g764 ( .A(n_758), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_759), .Y(n_765) );
AO22x2_ASAP7_75t_L g766 ( .A1(n_764), .A2(n_750), .B1(n_751), .B2(n_756), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_764), .A2(n_761), .B1(n_755), .B2(n_753), .C(n_760), .Y(n_767) );
AO22x2_ASAP7_75t_L g768 ( .A1(n_766), .A2(n_765), .B1(n_763), .B2(n_760), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_767), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_769), .B(n_744), .Y(n_770) );
NOR2xp67_ASAP7_75t_L g771 ( .A(n_768), .B(n_757), .Y(n_771) );
INVx4_ASAP7_75t_L g772 ( .A(n_770), .Y(n_772) );
INVx2_ASAP7_75t_L g773 ( .A(n_771), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_772), .A2(n_768), .B1(n_734), .B2(n_738), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_774), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_775), .A2(n_772), .B1(n_773), .B2(n_747), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_776), .Y(n_777) );
AO22x2_ASAP7_75t_L g778 ( .A1(n_777), .A2(n_744), .B1(n_732), .B2(n_745), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_779), .A2(n_745), .B1(n_721), .B2(n_722), .C(n_726), .Y(n_780) );
AOI211xp5_ASAP7_75t_L g781 ( .A1(n_780), .A2(n_713), .B(n_733), .C(n_723), .Y(n_781) );
endmodule