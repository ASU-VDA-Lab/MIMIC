module fake_jpeg_2535_n_573 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_573);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_573;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_59),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_17),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_87),
.Y(n_132)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_63),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_79),
.Y(n_162)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_80),
.Y(n_126)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_18),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_16),
.Y(n_117)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_40),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_19),
.Y(n_146)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_97),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_27),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_105),
.Y(n_135)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_102),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_23),
.B(n_18),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_36),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_107),
.B(n_71),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_36),
.B1(n_81),
.B2(n_27),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_110),
.B(n_144),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_23),
.B(n_47),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_149),
.B(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_117),
.B(n_131),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_53),
.A2(n_28),
.B1(n_47),
.B2(n_44),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_119),
.A2(n_141),
.B1(n_155),
.B2(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_28),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_55),
.A2(n_19),
.B1(n_39),
.B2(n_34),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_45),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_98),
.B(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_79),
.B(n_45),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_54),
.A2(n_65),
.B1(n_57),
.B2(n_64),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_82),
.B(n_15),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_69),
.B(n_15),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_73),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_63),
.A2(n_19),
.B1(n_39),
.B2(n_34),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_56),
.A2(n_34),
.B1(n_31),
.B2(n_39),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_31),
.B1(n_50),
.B2(n_46),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_132),
.A2(n_68),
.B1(n_66),
.B2(n_88),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_171),
.A2(n_215),
.B1(n_167),
.B2(n_125),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_172),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_173),
.Y(n_269)
);

OA22x2_ASAP7_75t_L g268 ( 
.A1(n_175),
.A2(n_195),
.B1(n_128),
.B2(n_30),
.Y(n_268)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_176),
.Y(n_275)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_124),
.Y(n_177)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_177),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_107),
.A2(n_38),
.B1(n_32),
.B2(n_50),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_197),
.Y(n_248)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_179),
.Y(n_283)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_180),
.Y(n_281)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_181),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_182),
.B(n_184),
.Y(n_243)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_93),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_152),
.A2(n_103),
.B(n_99),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_185),
.A2(n_190),
.B(n_143),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_186),
.B(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_133),
.Y(n_189)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

O2A1O1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_42),
.B(n_32),
.C(n_33),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_135),
.B(n_93),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_194),
.B(n_216),
.Y(n_262)
);

OAI22xp33_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_90),
.B1(n_94),
.B2(n_136),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_148),
.Y(n_196)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_198),
.Y(n_257)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_199),
.Y(n_286)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_200),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_148),
.A2(n_31),
.B1(n_50),
.B2(n_46),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_202),
.A2(n_217),
.B1(n_222),
.B2(n_227),
.Y(n_252)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_154),
.Y(n_203)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_127),
.B(n_46),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_224),
.Y(n_239)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_208),
.B(n_209),
.Y(n_265)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_166),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_210),
.B(n_223),
.Y(n_261)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_109),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_211),
.Y(n_250)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_212),
.B(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_214),
.Y(n_235)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_162),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_127),
.A2(n_159),
.B1(n_126),
.B2(n_134),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_135),
.B(n_70),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_140),
.A2(n_42),
.B1(n_38),
.B2(n_37),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_225),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_220),
.Y(n_272)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_221),
.Y(n_273)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_124),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_158),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_137),
.B(n_42),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_37),
.C(n_33),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_226),
.B(n_30),
.C(n_3),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_118),
.A2(n_38),
.B1(n_37),
.B2(n_33),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_123),
.B(n_32),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_162),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_138),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_125),
.B(n_29),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_231),
.B(n_232),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_166),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_233),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_282),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_121),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_238),
.B(n_244),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_172),
.B(n_157),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_259),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_251),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_192),
.A2(n_160),
.B1(n_157),
.B2(n_156),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_253),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_156),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_254),
.B(n_280),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_187),
.B(n_129),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_187),
.B(n_129),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_274),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_224),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_271),
.B(n_173),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_128),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_230),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_178),
.B1(n_173),
.B2(n_231),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_197),
.A2(n_30),
.B1(n_1),
.B2(n_3),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_277),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_193),
.B(n_201),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_226),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_197),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_174),
.B(n_0),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_175),
.A2(n_30),
.B1(n_6),
.B2(n_8),
.Y(n_282)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_288),
.A2(n_297),
.B1(n_298),
.B2(n_305),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_290),
.B(n_285),
.Y(n_375)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_292),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_183),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_294),
.B(n_296),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_222),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_238),
.A2(n_201),
.B1(n_195),
.B2(n_202),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_238),
.A2(n_196),
.B1(n_223),
.B2(n_225),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_242),
.A2(n_244),
.B1(n_259),
.B2(n_263),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_299),
.A2(n_318),
.B1(n_330),
.B2(n_331),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_265),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_300),
.B(n_303),
.Y(n_358)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_301),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_302),
.B(n_313),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_265),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_239),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_307),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_239),
.B1(n_248),
.B2(n_245),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_248),
.B(n_207),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_306),
.B(n_241),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_209),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_261),
.Y(n_308)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_308),
.Y(n_365)
);

INVx8_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_309),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_238),
.B(n_190),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_310),
.B(n_311),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_200),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_314),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_260),
.B(n_203),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_320),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_199),
.B1(n_208),
.B2(n_220),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_316),
.A2(n_325),
.B1(n_298),
.B2(n_297),
.Y(n_354)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_317),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_248),
.A2(n_252),
.B1(n_268),
.B2(n_282),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_279),
.B(n_214),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_275),
.B(n_212),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_229),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_326),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_257),
.B(n_221),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_329),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_246),
.B(n_211),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_268),
.A2(n_282),
.B1(n_250),
.B2(n_273),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_282),
.A2(n_180),
.B1(n_219),
.B2(n_177),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_250),
.A2(n_219),
.B1(n_6),
.B2(n_9),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_336),
.A2(n_272),
.B1(n_270),
.B2(n_273),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_334),
.A2(n_249),
.B(n_235),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_363),
.B(n_349),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_342),
.B(n_361),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_375),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_322),
.A2(n_272),
.B1(n_258),
.B2(n_270),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_347),
.A2(n_300),
.B1(n_292),
.B2(n_319),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_325),
.A2(n_281),
.B1(n_286),
.B2(n_255),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_348),
.A2(n_355),
.B1(n_368),
.B2(n_301),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_286),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_352),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_266),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_354),
.A2(n_360),
.B1(n_331),
.B2(n_324),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_295),
.A2(n_266),
.B1(n_247),
.B2(n_240),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_308),
.A2(n_247),
.B1(n_240),
.B2(n_236),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_304),
.B(n_237),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_334),
.A2(n_267),
.B(n_237),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_307),
.B(n_236),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_370),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_295),
.A2(n_287),
.B1(n_267),
.B2(n_256),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_293),
.B(n_287),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_318),
.A2(n_335),
.B1(n_299),
.B2(n_330),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_371),
.Y(n_380)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_373),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_293),
.B(n_5),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_378),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_320),
.B(n_302),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_321),
.Y(n_379)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_376),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_383),
.Y(n_417)
);

AO21x2_ASAP7_75t_SL g384 ( 
.A1(n_337),
.A2(n_332),
.B(n_303),
.Y(n_384)
);

AOI22x1_ASAP7_75t_L g441 ( 
.A1(n_384),
.A2(n_347),
.B1(n_377),
.B2(n_376),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_388),
.B(n_392),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_349),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_290),
.C(n_306),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_391),
.B(n_403),
.C(n_409),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_340),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_351),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_393),
.B(n_394),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_357),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_327),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_395),
.B(n_404),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_340),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_397),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_341),
.B(n_361),
.Y(n_398)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_399),
.A2(n_355),
.B1(n_350),
.B2(n_373),
.Y(n_440)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_400),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_372),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_401),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_341),
.B(n_312),
.Y(n_402)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_291),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_327),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_405),
.Y(n_433)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_359),
.B(n_289),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_407),
.B(n_357),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_345),
.A2(n_335),
.B(n_311),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_408),
.A2(n_414),
.B(n_358),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_289),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_367),
.B(n_315),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_410),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_362),
.B(n_314),
.C(n_332),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_415),
.C(n_339),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_370),
.B(n_336),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_413),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_351),
.B(n_309),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_337),
.A2(n_333),
.B1(n_285),
.B2(n_9),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_416),
.A2(n_342),
.B1(n_350),
.B2(n_379),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_409),
.B(n_338),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_434),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_387),
.A2(n_346),
.B1(n_345),
.B2(n_371),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_424),
.A2(n_431),
.B1(n_436),
.B2(n_399),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_426),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_428),
.A2(n_445),
.B(n_446),
.Y(n_451)
);

XOR2x1_ASAP7_75t_SL g471 ( 
.A(n_430),
.B(n_388),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_387),
.A2(n_380),
.B1(n_384),
.B2(n_408),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_432),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_382),
.B(n_352),
.C(n_356),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_380),
.A2(n_348),
.B1(n_368),
.B2(n_356),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_352),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_437),
.B(n_439),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_382),
.B(n_374),
.Y(n_439)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_440),
.Y(n_453)
);

A2O1A1Ixp33_ASAP7_75t_SL g460 ( 
.A1(n_441),
.A2(n_411),
.B(n_390),
.C(n_410),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_443),
.B(n_396),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_403),
.B(n_366),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_444),
.B(n_415),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_384),
.A2(n_365),
.B(n_377),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_369),
.B(n_333),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_384),
.A2(n_369),
.B(n_6),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_449),
.A2(n_400),
.B(n_386),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_423),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_450),
.B(n_460),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_452),
.A2(n_427),
.B1(n_429),
.B2(n_440),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_454),
.B(n_422),
.Y(n_495)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_419),
.Y(n_455)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_448),
.A2(n_398),
.B1(n_390),
.B2(n_402),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_457),
.A2(n_470),
.B1(n_472),
.B2(n_477),
.Y(n_483)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_458),
.Y(n_481)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_459),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_461),
.B(n_467),
.Y(n_479)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_417),
.Y(n_464)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_412),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g480 ( 
.A(n_465),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_425),
.B(n_396),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_466),
.Y(n_491)
);

AOI322xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_389),
.A3(n_413),
.B1(n_411),
.B2(n_397),
.C1(n_392),
.C2(n_401),
.Y(n_467)
);

INVx13_ASAP7_75t_L g468 ( 
.A(n_421),
.Y(n_468)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_468),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_414),
.Y(n_469)
);

AOI21xp33_ASAP7_75t_L g499 ( 
.A1(n_469),
.A2(n_10),
.B(n_11),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_448),
.A2(n_424),
.B1(n_438),
.B2(n_449),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_420),
.B1(n_430),
.B2(n_445),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_406),
.B1(n_416),
.B2(n_381),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_426),
.B(n_383),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_473),
.B(n_474),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_428),
.B(n_405),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_475),
.A2(n_476),
.B(n_447),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_386),
.B(n_385),
.Y(n_476)
);

INVx13_ASAP7_75t_L g477 ( 
.A(n_417),
.Y(n_477)
);

CKINVDCx14_ASAP7_75t_R g514 ( 
.A(n_482),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_484),
.A2(n_489),
.B1(n_456),
.B2(n_476),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_495),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_452),
.A2(n_420),
.B1(n_436),
.B2(n_441),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_418),
.C(n_437),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_494),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_456),
.A2(n_432),
.B1(n_441),
.B2(n_446),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_493),
.A2(n_470),
.B1(n_456),
.B2(n_472),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_418),
.C(n_434),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_478),
.B(n_444),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_496),
.B(n_500),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_463),
.B(n_439),
.C(n_385),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_498),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_5),
.C(n_10),
.Y(n_498)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_459),
.B(n_10),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_490),
.B(n_453),
.C(n_451),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_505),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_497),
.C(n_496),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_506),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_486),
.Y(n_507)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_507),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_480),
.B(n_453),
.C(n_451),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_486),
.C(n_492),
.Y(n_528)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_501),
.Y(n_510)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_510),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_511),
.Y(n_527)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_487),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_513),
.B(n_500),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_469),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_482),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_450),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_516),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_479),
.B(n_461),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_517),
.B(n_518),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_520),
.A2(n_521),
.B1(n_485),
.B2(n_460),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_483),
.A2(n_475),
.B1(n_457),
.B2(n_460),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_523),
.B(n_519),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_492),
.B(n_488),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_524),
.B(n_481),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_484),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_528),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_529),
.B(n_530),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_509),
.B(n_493),
.C(n_489),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_532),
.A2(n_534),
.B1(n_460),
.B2(n_512),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_503),
.A2(n_520),
.B1(n_508),
.B2(n_516),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_535),
.B(n_505),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_485),
.C(n_464),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_526),
.Y(n_541)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_511),
.C(n_507),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_539),
.B(n_540),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_521),
.C(n_512),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_543),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_542),
.A2(n_547),
.B1(n_524),
.B2(n_532),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_533),
.A2(n_460),
.B1(n_498),
.B2(n_468),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_528),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_527),
.A2(n_481),
.B1(n_502),
.B2(n_458),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_519),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_548),
.B(n_523),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_529),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_550),
.B(n_551),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_527),
.C(n_525),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_552),
.A2(n_539),
.B(n_536),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_553),
.A2(n_543),
.B1(n_549),
.B2(n_522),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_545),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_557),
.A2(n_546),
.B(n_544),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_558),
.A2(n_551),
.B(n_550),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_559),
.B(n_560),
.Y(n_564)
);

AOI31xp33_ASAP7_75t_L g565 ( 
.A1(n_562),
.A2(n_561),
.A3(n_555),
.B(n_554),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_563),
.A2(n_565),
.B(n_564),
.Y(n_566)
);

OAI211xp5_ASAP7_75t_L g568 ( 
.A1(n_566),
.A2(n_567),
.B(n_455),
.C(n_12),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_563),
.A2(n_559),
.B(n_477),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_568),
.A2(n_11),
.B(n_12),
.Y(n_569)
);

AOI21x1_ASAP7_75t_L g570 ( 
.A1(n_569),
.A2(n_11),
.B(n_12),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_13),
.C(n_14),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_13),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_13),
.B(n_14),
.Y(n_573)
);


endmodule