module real_jpeg_27064_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_0),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_0),
.A2(n_93),
.B(n_167),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_1),
.A2(n_80),
.B1(n_81),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_1),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_152),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_152),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_1),
.A2(n_33),
.B1(n_36),
.B2(n_152),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_2),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_3),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_47),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_3),
.A2(n_47),
.B(n_190),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_150),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_3),
.A2(n_10),
.B(n_33),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_3),
.B(n_99),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_3),
.A2(n_63),
.B1(n_122),
.B2(n_238),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_5),
.A2(n_80),
.B1(n_81),
.B2(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_5),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_132),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_132),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_5),
.A2(n_33),
.B1(n_36),
.B2(n_132),
.Y(n_230)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_6),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_7),
.A2(n_27),
.B1(n_30),
.B2(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_33),
.B1(n_36),
.B2(n_58),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_29),
.B1(n_33),
.B2(n_36),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_29),
.B1(n_80),
.B2(n_81),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_8),
.A2(n_29),
.B1(n_47),
.B2(n_48),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_43),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_43),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_9),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_101)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_11),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_56),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_11),
.A2(n_33),
.B1(n_36),
.B2(n_56),
.Y(n_167)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_46)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_52),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_14),
.A2(n_80),
.B1(n_81),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_14),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_106),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_14),
.A2(n_27),
.B1(n_30),
.B2(n_106),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_14),
.A2(n_33),
.B1(n_36),
.B2(n_106),
.Y(n_225)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_134),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_20),
.B(n_109),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_89),
.B2(n_108),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_44),
.B(n_59),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_44),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_25),
.A2(n_40),
.B(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_26),
.Y(n_143)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_27),
.B(n_53),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_27),
.A2(n_35),
.B(n_150),
.C(n_217),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_30),
.A2(n_48),
.A3(n_52),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_31),
.B(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_32),
.A2(n_40),
.B1(n_72),
.B2(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_32),
.A2(n_38),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_32),
.A2(n_40),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_32),
.A2(n_40),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_32),
.A2(n_40),
.B1(n_197),
.B2(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_32),
.B(n_150),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_36),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_40),
.A2(n_73),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_45),
.A2(n_51),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_45),
.A2(n_51),
.B1(n_146),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_45),
.A2(n_51),
.B1(n_176),
.B2(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_48),
.B1(n_78),
.B2(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_47),
.B(n_78),
.Y(n_164)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_48),
.A2(n_82),
.B1(n_149),
.B2(n_164),
.Y(n_163)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_51),
.B(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_51),
.B(n_127),
.Y(n_161)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_74),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_71),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_75),
.B1(n_76),
.B2(n_88),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_71),
.B1(n_88),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_66),
.B(n_69),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_63),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_63),
.A2(n_119),
.B1(n_122),
.B2(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_63),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_63),
.A2(n_95),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_63),
.A2(n_68),
.B1(n_230),
.B2(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_64),
.B(n_150),
.Y(n_242)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_67),
.A2(n_188),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_70),
.A2(n_121),
.B(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_85),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_77),
.A2(n_83),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_80),
.Y(n_82)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_80),
.B(n_150),
.CON(n_149),
.SN(n_149)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_104),
.B1(n_105),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_86),
.A2(n_104),
.B1(n_131),
.B2(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_86),
.B(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_102),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_91),
.B(n_96),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_114),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_116),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_124),
.C(n_129),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_117),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_123),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_123),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_124),
.A2(n_129),
.B1(n_130),
.B2(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_124),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_128),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_275),
.B(n_280),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_180),
.B(n_261),
.C(n_274),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_168),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_137),
.B(n_168),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_153),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_139),
.B(n_140),
.C(n_153),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_148),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_151),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_162),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_155),
.B(n_159),
.C(n_162),
.Y(n_272)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_169),
.A2(n_170),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_178),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_203),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_177),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_260),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_253),
.B(n_259),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_208),
.B(n_252),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_199),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_184),
.B(n_199),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.C(n_195),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_185),
.A2(n_186),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_189),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_200),
.B(n_206),
.C(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_246),
.B(n_251),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_226),
.B(n_245),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_218),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_212),
.A2(n_213),
.B1(n_216),
.B2(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_225),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_244),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_232),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_232),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_239),
.B(n_243),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_247),
.B(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_254),
.B(n_255),
.Y(n_259)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_262),
.B(n_263),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_272),
.B2(n_273),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_269),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);


endmodule