module fake_jpeg_8841_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_27),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_18),
.B1(n_36),
.B2(n_32),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_42),
.B1(n_53),
.B2(n_36),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_18),
.B1(n_26),
.B2(n_22),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_49),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_20),
.B1(n_26),
.B2(n_22),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_37),
.B1(n_19),
.B2(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_20),
.B1(n_25),
.B2(n_24),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_62),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_31),
.B(n_39),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_43),
.B1(n_33),
.B2(n_35),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_65),
.B1(n_74),
.B2(n_32),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_61),
.B(n_70),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_68),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_45),
.B1(n_52),
.B2(n_43),
.Y(n_83)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_31),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_28),
.B(n_52),
.C(n_45),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_73),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_37),
.B1(n_32),
.B2(n_30),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_0),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_0),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_1),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_29),
.B1(n_21),
.B2(n_15),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_27),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_89),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_52),
.A3(n_28),
.B1(n_33),
.B2(n_35),
.Y(n_87)
);

NOR3xp33_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_66),
.C(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_23),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_97),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_104),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_33),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_102),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_57),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_68),
.B1(n_54),
.B2(n_77),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_56),
.B(n_33),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_108),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_114),
.B(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_82),
.A2(n_62),
.B1(n_75),
.B2(n_61),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_121),
.B1(n_126),
.B2(n_103),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_76),
.C(n_69),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_93),
.C(n_88),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_127),
.B1(n_80),
.B2(n_103),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_57),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_35),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_123),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_80),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_98),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_67),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_87),
.B(n_98),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_84),
.A2(n_33),
.B1(n_66),
.B2(n_30),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_132),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_143),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_110),
.B1(n_84),
.B2(n_112),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_136),
.A2(n_150),
.B1(n_148),
.B2(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_145),
.C(n_147),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_146),
.B1(n_99),
.B2(n_123),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_106),
.A2(n_89),
.B(n_102),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_149),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_118),
.CI(n_111),
.CON(n_143),
.SN(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_118),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_94),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_152),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_100),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_102),
.B1(n_94),
.B2(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_157),
.A2(n_166),
.B1(n_169),
.B2(n_171),
.Y(n_172)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_161),
.Y(n_173)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_170),
.B1(n_137),
.B2(n_149),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_105),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_129),
.C(n_143),
.Y(n_179)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_132),
.A2(n_125),
.B1(n_108),
.B2(n_104),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_147),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_181),
.Y(n_191)
);

AOI21x1_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_142),
.B(n_131),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_184),
.B(n_8),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_176),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_165),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_3),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_180),
.C(n_3),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_156),
.Y(n_180)
);

OAI322xp33_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_143),
.A3(n_158),
.B1(n_164),
.B2(n_168),
.C1(n_153),
.C2(n_170),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_139),
.B1(n_60),
.B2(n_66),
.Y(n_183)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_163),
.A2(n_60),
.B1(n_66),
.B2(n_21),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_2),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_8),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_186),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_160),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_193),
.B1(n_184),
.B2(n_178),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_7),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_195),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_8),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_180),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_191),
.C(n_194),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_192),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_205),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_198),
.B(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_213),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_210),
.B(n_199),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_199),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_197),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_219),
.A2(n_220),
.A3(n_221),
.B1(n_216),
.B2(n_200),
.C1(n_195),
.C2(n_12),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_214),
.A2(n_208),
.B1(n_191),
.B2(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_9),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_10),
.Y(n_228)
);


endmodule