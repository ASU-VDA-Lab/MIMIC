module fake_jpeg_28117_n_181 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_1),
.B(n_4),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_30),
.B(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_34),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_15),
.B1(n_26),
.B2(n_17),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_56),
.B1(n_41),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_32),
.A2(n_16),
.B1(n_15),
.B2(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_18),
.B1(n_27),
.B2(n_36),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_54),
.B(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_22),
.B2(n_18),
.Y(n_56)
);

AO22x1_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_16),
.B1(n_28),
.B2(n_31),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_59),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_63),
.Y(n_96)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_38),
.B1(n_37),
.B2(n_40),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_24),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_72),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_48),
.B(n_27),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_41),
.C(n_39),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_33),
.B1(n_43),
.B2(n_30),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_52),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_28),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_23),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_28),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_40),
.B1(n_41),
.B2(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_84),
.B1(n_45),
.B2(n_33),
.Y(n_90)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_100),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_45),
.B1(n_47),
.B2(n_39),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_77),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_28),
.B1(n_31),
.B2(n_30),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_80),
.B1(n_62),
.B2(n_61),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_29),
.B(n_33),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_65),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_29),
.Y(n_103)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_108),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_75),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_112),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_104),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_118),
.B1(n_119),
.B2(n_98),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_86),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_123),
.C(n_91),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_29),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_63),
.B1(n_62),
.B2(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_23),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_122),
.A2(n_87),
.B(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_131),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_103),
.C(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_29),
.C(n_73),
.Y(n_147)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_133),
.C(n_126),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_97),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_3),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_106),
.B1(n_114),
.B2(n_119),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_87),
.B1(n_85),
.B2(n_101),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_116),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_135),
.Y(n_157)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_144),
.B(n_132),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_138),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_146),
.Y(n_153)
);

AOI322xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_120),
.A3(n_116),
.B1(n_108),
.B2(n_33),
.C1(n_72),
.C2(n_101),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_145),
.A2(n_149),
.B1(n_137),
.B2(n_134),
.Y(n_151)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_147),
.B(n_148),
.C(n_125),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_71),
.C(n_9),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_130),
.B(n_131),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_154),
.B(n_155),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_148),
.C(n_10),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_139),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_5),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_145),
.A2(n_149),
.B1(n_141),
.B2(n_147),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_162),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_141),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_164),
.C(n_165),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_7),
.C(n_9),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_153),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_151),
.C(n_162),
.Y(n_172)
);

AOI31xp67_ASAP7_75t_L g169 ( 
.A1(n_165),
.A2(n_158),
.A3(n_156),
.B(n_159),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_170),
.B(n_171),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_163),
.B(n_6),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_173),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_175),
.B(n_12),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_13),
.B(n_7),
.Y(n_175)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_176),
.Y(n_178)
);

NOR2xp67_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_11),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_12),
.B(n_5),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_178),
.Y(n_181)
);


endmodule