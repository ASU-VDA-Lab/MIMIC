module fake_jpeg_11632_n_56 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_56);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_56;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_8),
.Y(n_20)
);

NAND2x1_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_17),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_8),
.A2(n_9),
.B1(n_1),
.B2(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_37),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_43)
);

OAI22x1_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_28),
.B1(n_21),
.B2(n_31),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_44),
.B(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_34),
.B1(n_7),
.B2(n_9),
.Y(n_48)
);

AO32x1_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_25),
.A3(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_R g44 ( 
.A(n_36),
.B(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_34),
.B1(n_10),
.B2(n_3),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.C(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_39),
.B(n_15),
.Y(n_50)
);

AO21x1_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_50),
.B(n_46),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_51),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_41),
.C(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_10),
.Y(n_56)
);


endmodule