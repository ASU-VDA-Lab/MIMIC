module fake_aes_2675_n_1267 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1267);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1267;
wire n_963;
wire n_1034;
wire n_949;
wire n_858;
wire n_646;
wire n_829;
wire n_1198;
wire n_667;
wire n_988;
wire n_311;
wire n_655;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_860;
wire n_1208;
wire n_305;
wire n_1201;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_830;
wire n_1112;
wire n_517;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_304;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_619;
wire n_501;
wire n_299;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_673;
wire n_1071;
wire n_1079;
wire n_315;
wire n_409;
wire n_295;
wire n_677;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_586;
wire n_1246;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_293;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_294;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_307;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_308;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_557;
wire n_842;
wire n_439;
wire n_614;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_306;
wire n_1007;
wire n_1117;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_867;
wire n_1070;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_287;
wire n_606;
wire n_332;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_284;
wire n_500;
wire n_607;
wire n_496;
wire n_801;
wire n_1059;
wire n_309;
wire n_701;
wire n_612;
wire n_1032;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_301;
wire n_609;
wire n_909;
wire n_366;
wire n_596;
wire n_1215;
wire n_286;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1254;
wire n_764;
wire n_426;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_427;
wire n_703;
wire n_415;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_285;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_300;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1043;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_290;
wire n_385;
wire n_1127;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_292;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_288;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_296;
wire n_765;
wire n_1177;
wire n_462;
wire n_783;
wire n_1074;
wire n_463;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_303;
wire n_326;
wire n_289;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_302;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_948;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_639;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_335;
wire n_700;
wire n_534;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_297;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_291;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1219;
wire n_1120;
wire n_595;
wire n_759;
wire n_559;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
INVxp67_ASAP7_75t_SL g284 ( .A(n_64), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_160), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_26), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_86), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_65), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_211), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_33), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_233), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_74), .Y(n_293) );
INVxp67_ASAP7_75t_SL g294 ( .A(n_221), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_73), .Y(n_295) );
BUFx5_ASAP7_75t_L g296 ( .A(n_245), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_59), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_250), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_224), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_238), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_172), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_157), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_28), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_260), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_31), .Y(n_307) );
BUFx10_ASAP7_75t_L g308 ( .A(n_141), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_198), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_165), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_66), .Y(n_311) );
NOR2xp67_ASAP7_75t_L g312 ( .A(n_115), .B(n_13), .Y(n_312) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_232), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_173), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_105), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_226), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_84), .Y(n_317) );
INVxp33_ASAP7_75t_L g318 ( .A(n_11), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_193), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_90), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_246), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_143), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_39), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_53), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_180), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_49), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_73), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_212), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_102), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_144), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_77), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_152), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_25), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_176), .Y(n_334) );
CKINVDCx14_ASAP7_75t_R g335 ( .A(n_162), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_145), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_39), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_108), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_32), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_147), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_65), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_49), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_239), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_2), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_137), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_87), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_251), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_130), .Y(n_348) );
INVxp67_ASAP7_75t_L g349 ( .A(n_2), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_80), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_253), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_266), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_79), .Y(n_353) );
BUFx8_ASAP7_75t_SL g354 ( .A(n_281), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_17), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_25), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_202), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_222), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_136), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_241), .Y(n_360) );
CKINVDCx14_ASAP7_75t_R g361 ( .A(n_37), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_278), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_142), .Y(n_363) );
NOR2xp67_ASAP7_75t_L g364 ( .A(n_169), .B(n_218), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_188), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_50), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_88), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_149), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_270), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_213), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_242), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_109), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_236), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_252), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_133), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_74), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_112), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_187), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_191), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_27), .Y(n_380) );
INVxp33_ASAP7_75t_SL g381 ( .A(n_163), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_216), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_186), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_33), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_272), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_129), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_7), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_125), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_215), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_29), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_199), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_139), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_13), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_282), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_106), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_124), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_189), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_228), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_257), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_127), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_117), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_263), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_42), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_177), .Y(n_404) );
INVx1_ASAP7_75t_SL g405 ( .A(n_71), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_91), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_244), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_60), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_94), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_230), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_52), .Y(n_411) );
CKINVDCx20_ASAP7_75t_R g412 ( .A(n_92), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_214), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_26), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g415 ( .A(n_37), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_219), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_63), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_43), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_17), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_267), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_227), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_113), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_93), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_290), .B(n_0), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_290), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_354), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_313), .Y(n_427) );
BUFx8_ASAP7_75t_L g428 ( .A(n_296), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_311), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_311), .Y(n_430) );
BUFx8_ASAP7_75t_L g431 ( .A(n_296), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_313), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_296), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_296), .Y(n_435) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_312), .B(n_0), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_313), .Y(n_437) );
OAI22x1_ASAP7_75t_R g438 ( .A1(n_341), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_393), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_323), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_318), .B(n_1), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_361), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_296), .Y(n_443) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_313), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_323), .B(n_5), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_324), .B(n_6), .Y(n_446) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_320), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_296), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_298), .B(n_6), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_296), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_343), .B(n_7), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_324), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_342), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_320), .Y(n_454) );
CKINVDCx11_ASAP7_75t_R g455 ( .A(n_341), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_318), .B(n_8), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_342), .Y(n_457) );
INVx5_ASAP7_75t_L g458 ( .A(n_320), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_308), .Y(n_459) );
BUFx2_ASAP7_75t_L g460 ( .A(n_428), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_434), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_459), .B(n_347), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_459), .B(n_356), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_424), .A2(n_295), .B1(n_307), .B2(n_288), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_434), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_459), .B(n_299), .Y(n_467) );
AND2x6_ASAP7_75t_L g468 ( .A(n_424), .B(n_377), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_459), .B(n_328), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_441), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_441), .B(n_335), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_425), .B(n_299), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_428), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_432), .B(n_301), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
INVx3_ASAP7_75t_L g478 ( .A(n_435), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_432), .B(n_301), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_443), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_432), .B(n_382), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_443), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_428), .B(n_382), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_431), .B(n_395), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_424), .Y(n_486) );
AND3x2_ASAP7_75t_L g487 ( .A(n_439), .B(n_284), .C(n_349), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_431), .B(n_308), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_427), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_448), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_431), .B(n_395), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_425), .B(n_401), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_431), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_427), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_456), .B(n_401), .Y(n_495) );
AOI22xp33_ASAP7_75t_SL g496 ( .A1(n_424), .A2(n_415), .B1(n_361), .B2(n_315), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_456), .B(n_422), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_445), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_427), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_427), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_448), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_426), .Y(n_502) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_445), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_448), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_427), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_433), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_463), .Y(n_508) );
O2A1O1Ixp5_ASAP7_75t_L g509 ( .A1(n_503), .A2(n_446), .B(n_445), .C(n_451), .Y(n_509) );
AOI22x1_ASAP7_75t_L g510 ( .A1(n_486), .A2(n_503), .B1(n_498), .B2(n_493), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_470), .B(n_426), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_472), .B(n_445), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_472), .B(n_446), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_495), .B(n_449), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_472), .B(n_446), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_460), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_497), .B(n_381), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_463), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_470), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_502), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_460), .B(n_374), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_498), .A2(n_450), .B1(n_430), .B2(n_440), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_497), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_468), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_463), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_469), .B(n_381), .Y(n_528) );
NAND3xp33_ASAP7_75t_SL g529 ( .A(n_496), .B(n_442), .C(n_305), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_498), .A2(n_450), .B1(n_430), .B2(n_440), .Y(n_530) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_475), .B(n_442), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_467), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_486), .B(n_374), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_486), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
AND2x6_ASAP7_75t_SL g536 ( .A(n_473), .B(n_455), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_475), .B(n_436), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_467), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_468), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_488), .B(n_378), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_462), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_468), .A2(n_315), .B1(n_345), .B2(n_291), .Y(n_542) );
AND2x4_ASAP7_75t_L g543 ( .A(n_493), .B(n_464), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_468), .A2(n_345), .B1(n_394), .B2(n_291), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_468), .B(n_398), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_466), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_468), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_468), .B(n_398), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_462), .B(n_429), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_493), .B(n_423), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_464), .B(n_436), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_484), .B(n_423), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g553 ( .A(n_473), .B(n_429), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_492), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_485), .B(n_452), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_485), .B(n_452), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g557 ( .A1(n_492), .A2(n_457), .B(n_453), .C(n_333), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_476), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_491), .B(n_453), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_491), .B(n_457), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_476), .B(n_287), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_479), .B(n_482), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_496), .A2(n_396), .B1(n_406), .B2(n_394), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_487), .B(n_293), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g565 ( .A(n_479), .B(n_308), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_466), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_461), .A2(n_337), .B1(n_339), .B2(n_326), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_482), .B(n_285), .Y(n_568) );
INVx8_ASAP7_75t_L g569 ( .A(n_466), .Y(n_569) );
AND2x6_ASAP7_75t_SL g570 ( .A(n_487), .B(n_438), .Y(n_570) );
INVx5_ASAP7_75t_L g571 ( .A(n_466), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_461), .A2(n_396), .B1(n_407), .B2(n_406), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_466), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_471), .A2(n_422), .B(n_321), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_471), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_477), .A2(n_344), .B1(n_384), .B2(n_376), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_480), .A2(n_407), .B1(n_413), .B2(n_412), .Y(n_577) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_480), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_481), .B(n_316), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_474), .B(n_289), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_481), .B(n_329), .Y(n_581) );
NAND2xp33_ASAP7_75t_L g582 ( .A(n_483), .B(n_330), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_483), .A2(n_408), .B1(n_418), .B2(n_387), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_504), .A2(n_413), .B1(n_412), .B2(n_355), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_504), .B(n_332), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_507), .B(n_474), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_474), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_507), .B(n_336), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_474), .B(n_338), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_474), .B(n_340), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_478), .Y(n_591) );
NOR2xp33_ASAP7_75t_R g592 ( .A(n_478), .B(n_415), .Y(n_592) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_478), .Y(n_593) );
OR2x6_ASAP7_75t_L g594 ( .A(n_478), .B(n_380), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_490), .A2(n_419), .B1(n_356), .B2(n_411), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_490), .A2(n_366), .B1(n_417), .B2(n_403), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_490), .B(n_390), .Y(n_597) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_509), .A2(n_501), .B(n_490), .C(n_411), .Y(n_598) );
BUFx2_ASAP7_75t_SL g599 ( .A(n_522), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_572), .B(n_286), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_525), .B(n_490), .Y(n_601) );
INVx4_ASAP7_75t_L g602 ( .A(n_569), .Y(n_602) );
INVx6_ASAP7_75t_L g603 ( .A(n_536), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_562), .A2(n_501), .B(n_294), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_529), .A2(n_501), .B1(n_297), .B2(n_300), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_538), .A2(n_501), .B1(n_390), .B2(n_414), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_529), .A2(n_405), .B(n_501), .C(n_303), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_512), .A2(n_304), .B(n_292), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_518), .B(n_350), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_521), .B(n_327), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_543), .A2(n_327), .B1(n_306), .B2(n_310), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_515), .B(n_354), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_511), .B(n_327), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g614 ( .A1(n_514), .A2(n_314), .B(n_309), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_515), .B(n_358), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_509), .A2(n_317), .B(n_322), .C(n_319), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_519), .B(n_302), .Y(n_617) );
INVx6_ASAP7_75t_L g618 ( .A(n_570), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_577), .B(n_327), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_519), .B(n_346), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_517), .A2(n_334), .B(n_325), .Y(n_621) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_569), .Y(n_622) );
OR2x6_ASAP7_75t_L g623 ( .A(n_594), .B(n_364), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_518), .B(n_359), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_555), .A2(n_351), .B(n_348), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_556), .A2(n_353), .B(n_352), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_541), .B(n_360), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_559), .A2(n_362), .B(n_357), .Y(n_628) );
BUFx2_ASAP7_75t_L g629 ( .A(n_592), .Y(n_629) );
INVx2_ASAP7_75t_SL g630 ( .A(n_594), .Y(n_630) );
AND2x2_ASAP7_75t_SL g631 ( .A(n_542), .B(n_363), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_539), .B(n_368), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_532), .B(n_369), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_528), .B(n_421), .Y(n_634) );
INVx6_ASAP7_75t_L g635 ( .A(n_597), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_584), .B(n_531), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_543), .A2(n_367), .B1(n_370), .B2(n_365), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g638 ( .A1(n_549), .A2(n_372), .B(n_373), .C(n_371), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_544), .A2(n_379), .B1(n_383), .B2(n_375), .Y(n_639) );
A2O1A1Ixp33_ASAP7_75t_L g640 ( .A1(n_549), .A2(n_386), .B(n_388), .C(n_385), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_SL g641 ( .A1(n_540), .A2(n_454), .B(n_494), .C(n_465), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g642 ( .A1(n_568), .A2(n_391), .B(n_392), .C(n_389), .Y(n_642) );
CKINVDCx5p33_ASAP7_75t_R g643 ( .A(n_594), .Y(n_643) );
AO21x1_ASAP7_75t_L g644 ( .A1(n_580), .A2(n_399), .B(n_397), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_539), .B(n_404), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_560), .A2(n_402), .B(n_400), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_568), .A2(n_410), .B(n_416), .C(n_409), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_578), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_563), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_526), .B(n_420), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_551), .B(n_8), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_558), .B(n_331), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_551), .B(n_9), .Y(n_653) );
INVx2_ASAP7_75t_SL g654 ( .A(n_569), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_596), .B(n_10), .Y(n_655) );
OAI21xp5_ASAP7_75t_L g656 ( .A1(n_535), .A2(n_506), .B(n_500), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_537), .B(n_11), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_575), .A2(n_454), .B1(n_331), .B2(n_458), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_571), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_547), .B(n_458), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_564), .B(n_12), .Y(n_661) );
OAI21xp33_ASAP7_75t_L g662 ( .A1(n_524), .A2(n_437), .B(n_433), .Y(n_662) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_574), .A2(n_500), .B(n_499), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_554), .B(n_12), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_508), .Y(n_665) );
INVx3_ASAP7_75t_L g666 ( .A(n_573), .Y(n_666) );
BUFx3_ASAP7_75t_L g667 ( .A(n_571), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_573), .Y(n_668) );
AO21x1_ASAP7_75t_L g669 ( .A1(n_580), .A2(n_500), .B(n_499), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_533), .A2(n_505), .B(n_499), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_513), .A2(n_516), .B1(n_527), .B2(n_520), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_593), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_593), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_552), .B(n_14), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_524), .A2(n_458), .B1(n_447), .B2(n_444), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_586), .Y(n_676) );
BUFx6f_ASAP7_75t_SL g677 ( .A(n_591), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g678 ( .A1(n_561), .A2(n_506), .B(n_505), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_530), .A2(n_458), .B1(n_447), .B2(n_444), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_553), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_565), .B(n_14), .Y(n_681) );
OAI21x1_ASAP7_75t_SL g682 ( .A1(n_510), .A2(n_506), .B(n_505), .Y(n_682) );
BUFx3_ASAP7_75t_L g683 ( .A(n_571), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_545), .B(n_548), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_530), .A2(n_447), .B(n_444), .C(n_437), .Y(n_685) );
OAI21x1_ASAP7_75t_L g686 ( .A1(n_546), .A2(n_489), .B(n_458), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_567), .B(n_458), .C(n_437), .Y(n_687) );
OR2x2_ASAP7_75t_L g688 ( .A(n_567), .B(n_15), .Y(n_688) );
A2O1A1Ixp33_ASAP7_75t_L g689 ( .A1(n_576), .A2(n_447), .B(n_444), .C(n_437), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_585), .A2(n_489), .B(n_437), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_566), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g692 ( .A1(n_588), .A2(n_489), .B(n_437), .Y(n_692) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_571), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_587), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_523), .B(n_15), .Y(n_695) );
A2O1A1Ixp33_ASAP7_75t_L g696 ( .A1(n_576), .A2(n_447), .B(n_444), .C(n_433), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_589), .Y(n_697) );
INVxp67_ASAP7_75t_SL g698 ( .A(n_582), .Y(n_698) );
NOR2xp33_ASAP7_75t_SL g699 ( .A(n_550), .B(n_433), .Y(n_699) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_590), .Y(n_700) );
NOR2xp33_ASAP7_75t_R g701 ( .A(n_583), .B(n_16), .Y(n_701) );
BUFx2_ASAP7_75t_L g702 ( .A(n_583), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_595), .B(n_16), .Y(n_703) );
BUFx12f_ASAP7_75t_L g704 ( .A(n_595), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_579), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_581), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_509), .A2(n_433), .B(n_489), .C(n_20), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_562), .A2(n_489), .B(n_78), .Y(n_708) );
O2A1O1Ixp33_ASAP7_75t_SL g709 ( .A1(n_557), .A2(n_138), .B(n_283), .C(n_280), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_562), .A2(n_489), .B(n_81), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_529), .A2(n_18), .B(n_19), .C(n_20), .Y(n_711) );
AND2x4_ASAP7_75t_L g712 ( .A(n_525), .B(n_18), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_538), .A2(n_19), .B1(n_21), .B2(n_22), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_525), .Y(n_714) );
INVx5_ASAP7_75t_L g715 ( .A(n_569), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_534), .Y(n_716) );
OAI21x1_ASAP7_75t_L g717 ( .A1(n_510), .A2(n_489), .B(n_82), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_525), .Y(n_718) );
OR2x6_ASAP7_75t_L g719 ( .A(n_572), .B(n_22), .Y(n_719) );
AOI21x1_ASAP7_75t_L g720 ( .A1(n_562), .A2(n_83), .B(n_76), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_534), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_525), .B(n_23), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_521), .B(n_23), .Y(n_723) );
O2A1O1Ixp5_ASAP7_75t_L g724 ( .A1(n_509), .A2(n_146), .B(n_277), .C(n_275), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_538), .A2(n_24), .B1(n_27), .B2(n_28), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g726 ( .A1(n_531), .A2(n_24), .B1(n_29), .B2(n_30), .Y(n_726) );
NAND3xp33_ASAP7_75t_SL g727 ( .A(n_522), .B(n_30), .C(n_31), .Y(n_727) );
O2A1O1Ixp33_ASAP7_75t_SL g728 ( .A1(n_598), .A2(n_150), .B(n_274), .C(n_271), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_648), .B(n_32), .Y(n_729) );
AO31x2_ASAP7_75t_L g730 ( .A1(n_669), .A2(n_34), .A3(n_35), .B(n_36), .Y(n_730) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_599), .Y(n_731) );
AOI221x1_ASAP7_75t_L g732 ( .A1(n_662), .A2(n_38), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g733 ( .A1(n_616), .A2(n_89), .B(n_85), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_631), .A2(n_38), .B1(n_40), .B2(n_41), .Y(n_734) );
INVx4_ASAP7_75t_L g735 ( .A(n_715), .Y(n_735) );
OAI21x1_ASAP7_75t_L g736 ( .A1(n_682), .A2(n_717), .B(n_686), .Y(n_736) );
AO31x2_ASAP7_75t_L g737 ( .A1(n_707), .A2(n_43), .A3(n_44), .B(n_45), .Y(n_737) );
INVx5_ASAP7_75t_L g738 ( .A(n_622), .Y(n_738) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_622), .Y(n_739) );
O2A1O1Ixp33_ASAP7_75t_SL g740 ( .A1(n_641), .A2(n_685), .B(n_696), .C(n_689), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_643), .Y(n_741) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_701), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_742) );
OAI22x1_ASAP7_75t_L g743 ( .A1(n_605), .A2(n_47), .B1(n_48), .B2(n_50), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_702), .A2(n_51), .B1(n_52), .B2(n_53), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_715), .B(n_51), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_670), .A2(n_692), .B(n_690), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_656), .A2(n_166), .B(n_269), .Y(n_747) );
OAI21xp5_ASAP7_75t_L g748 ( .A1(n_604), .A2(n_164), .B(n_268), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g749 ( .A1(n_726), .A2(n_54), .B1(n_55), .B2(n_56), .C1(n_57), .C2(n_58), .Y(n_749) );
BUFx2_ASAP7_75t_SL g750 ( .A(n_715), .Y(n_750) );
OAI22x1_ASAP7_75t_L g751 ( .A1(n_605), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_607), .A2(n_57), .B(n_58), .C(n_59), .Y(n_752) );
BUFx12f_ASAP7_75t_L g753 ( .A(n_603), .Y(n_753) );
NAND2x1p5_ASAP7_75t_L g754 ( .A(n_602), .B(n_60), .Y(n_754) );
AO32x2_ASAP7_75t_L g755 ( .A1(n_611), .A2(n_61), .A3(n_62), .B1(n_63), .B2(n_64), .Y(n_755) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_618), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_656), .A2(n_174), .B(n_264), .Y(n_757) );
CKINVDCx11_ASAP7_75t_R g758 ( .A(n_719), .Y(n_758) );
BUFx12f_ASAP7_75t_L g759 ( .A(n_603), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_678), .A2(n_175), .B(n_262), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g761 ( .A1(n_724), .A2(n_171), .B(n_261), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_613), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_712), .Y(n_763) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_726), .A2(n_67), .B1(n_68), .B2(n_69), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_676), .B(n_68), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_649), .B(n_612), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_627), .A2(n_170), .B(n_259), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_602), .Y(n_768) );
OA21x2_ASAP7_75t_L g769 ( .A1(n_662), .A2(n_168), .B(n_258), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_714), .B(n_69), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_712), .Y(n_771) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_651), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_708), .A2(n_178), .B(n_256), .Y(n_773) );
INVx2_ASAP7_75t_SL g774 ( .A(n_622), .Y(n_774) );
A2O1A1Ixp33_ASAP7_75t_L g775 ( .A1(n_608), .A2(n_75), .B(n_95), .C(n_96), .Y(n_775) );
INVx4_ASAP7_75t_L g776 ( .A(n_659), .Y(n_776) );
AO31x2_ASAP7_75t_L g777 ( .A1(n_644), .A2(n_97), .A3(n_98), .B(n_99), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_718), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_SL g779 ( .A1(n_647), .A2(n_100), .B(n_101), .C(n_103), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_630), .Y(n_780) );
A2O1A1Ixp33_ASAP7_75t_L g781 ( .A1(n_614), .A2(n_104), .B(n_107), .C(n_110), .Y(n_781) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_654), .B(n_111), .Y(n_782) );
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_719), .A2(n_114), .B1(n_116), .B2(n_118), .Y(n_783) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_615), .A2(n_119), .B(n_120), .Y(n_784) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_659), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g786 ( .A1(n_719), .A2(n_121), .B1(n_122), .B2(n_123), .Y(n_786) );
BUFx2_ASAP7_75t_L g787 ( .A(n_704), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_618), .B(n_126), .Y(n_788) );
OAI22xp33_ASAP7_75t_L g789 ( .A1(n_653), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_789) );
OAI22xp33_ASAP7_75t_SL g790 ( .A1(n_600), .A2(n_134), .B1(n_135), .B2(n_140), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_664), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_637), .B(n_148), .Y(n_792) );
INVx3_ASAP7_75t_L g793 ( .A(n_659), .Y(n_793) );
NOR2xp33_ASAP7_75t_SL g794 ( .A(n_629), .B(n_151), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_610), .Y(n_795) );
O2A1O1Ixp33_ASAP7_75t_SL g796 ( .A1(n_674), .A2(n_153), .B(n_154), .C(n_155), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_688), .Y(n_797) );
OAI22x1_ASAP7_75t_L g798 ( .A1(n_681), .A2(n_156), .B1(n_158), .B2(n_159), .Y(n_798) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_601), .Y(n_799) );
INVxp67_ASAP7_75t_L g800 ( .A(n_723), .Y(n_800) );
CKINVDCx9p33_ASAP7_75t_R g801 ( .A(n_657), .Y(n_801) );
NAND2xp33_ASAP7_75t_L g802 ( .A(n_672), .B(n_161), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_716), .Y(n_803) );
CKINVDCx6p67_ASAP7_75t_R g804 ( .A(n_623), .Y(n_804) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_635), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_660), .A2(n_167), .B(n_179), .Y(n_806) );
AO31x2_ASAP7_75t_L g807 ( .A1(n_710), .A2(n_181), .A3(n_182), .B(n_183), .Y(n_807) );
BUFx10_ASAP7_75t_L g808 ( .A(n_681), .Y(n_808) );
NAND2xp33_ASAP7_75t_L g809 ( .A(n_673), .B(n_184), .Y(n_809) );
O2A1O1Ixp33_ASAP7_75t_L g810 ( .A1(n_711), .A2(n_185), .B(n_190), .C(n_192), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_721), .Y(n_811) );
AO31x2_ASAP7_75t_L g812 ( .A1(n_675), .A2(n_194), .A3(n_195), .B(n_196), .Y(n_812) );
A2O1A1Ixp33_ASAP7_75t_L g813 ( .A1(n_621), .A2(n_197), .B(n_200), .C(n_201), .Y(n_813) );
OAI21x1_ASAP7_75t_L g814 ( .A1(n_720), .A2(n_203), .B(n_204), .Y(n_814) );
BUFx3_ASAP7_75t_L g815 ( .A(n_667), .Y(n_815) );
O2A1O1Ixp33_ASAP7_75t_SL g816 ( .A1(n_652), .A2(n_205), .B(n_206), .C(n_207), .Y(n_816) );
OAI21x1_ASAP7_75t_L g817 ( .A1(n_663), .A2(n_208), .B(n_209), .Y(n_817) );
NOR2xp33_ASAP7_75t_SL g818 ( .A(n_636), .B(n_210), .Y(n_818) );
INVx3_ASAP7_75t_L g819 ( .A(n_683), .Y(n_819) );
AO31x2_ASAP7_75t_L g820 ( .A1(n_679), .A2(n_217), .A3(n_220), .B(n_223), .Y(n_820) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_625), .A2(n_225), .B(n_229), .Y(n_821) );
NAND2xp33_ASAP7_75t_L g822 ( .A(n_697), .B(n_231), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_635), .A2(n_234), .B1(n_235), .B2(n_237), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_671), .B(n_240), .Y(n_824) );
OA22x2_ASAP7_75t_L g825 ( .A1(n_623), .A2(n_243), .B1(n_247), .B2(n_248), .Y(n_825) );
INVx2_ASAP7_75t_L g826 ( .A(n_665), .Y(n_826) );
AOI21x1_ASAP7_75t_L g827 ( .A1(n_626), .A2(n_249), .B(n_254), .Y(n_827) );
AO31x2_ASAP7_75t_L g828 ( .A1(n_713), .A2(n_725), .A3(n_606), .B(n_703), .Y(n_828) );
CKINVDCx11_ASAP7_75t_R g829 ( .A(n_623), .Y(n_829) );
OA21x2_ASAP7_75t_L g830 ( .A1(n_687), .A2(n_255), .B(n_279), .Y(n_830) );
INVx2_ASAP7_75t_L g831 ( .A(n_691), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_661), .A2(n_639), .B1(n_617), .B2(n_620), .C(n_619), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_628), .A2(n_646), .B(n_698), .Y(n_833) );
OAI21xp5_ASAP7_75t_L g834 ( .A1(n_687), .A2(n_694), .B(n_680), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_655), .B(n_633), .Y(n_835) );
AND2x4_ASAP7_75t_L g836 ( .A(n_705), .B(n_706), .Y(n_836) );
AO31x2_ASAP7_75t_L g837 ( .A1(n_658), .A2(n_695), .A3(n_722), .B(n_634), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_609), .B(n_624), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_668), .A2(n_650), .B(n_645), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_693), .A2(n_666), .B1(n_700), .B2(n_677), .Y(n_840) );
NOR4xp25_ASAP7_75t_L g841 ( .A(n_727), .B(n_709), .C(n_666), .D(n_632), .Y(n_841) );
INVx3_ASAP7_75t_L g842 ( .A(n_677), .Y(n_842) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_699), .A2(n_493), .B(n_684), .Y(n_843) );
O2A1O1Ixp33_ASAP7_75t_L g844 ( .A1(n_700), .A2(n_640), .B(n_638), .C(n_607), .Y(n_844) );
AO31x2_ASAP7_75t_L g845 ( .A1(n_669), .A2(n_707), .A3(n_644), .B(n_598), .Y(n_845) );
OAI21x1_ASAP7_75t_SL g846 ( .A1(n_644), .A2(n_518), .B(n_664), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_648), .B(n_525), .Y(n_847) );
OAI21x1_ASAP7_75t_L g848 ( .A1(n_682), .A2(n_717), .B(n_686), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_702), .A2(n_653), .B1(n_651), .B2(n_543), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_613), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_649), .B(n_531), .Y(n_851) );
INVx3_ASAP7_75t_L g852 ( .A(n_715), .Y(n_852) );
CKINVDCx11_ASAP7_75t_R g853 ( .A(n_719), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_648), .B(n_525), .Y(n_854) );
O2A1O1Ixp33_ASAP7_75t_L g855 ( .A1(n_638), .A2(n_640), .B(n_607), .C(n_642), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g856 ( .A(n_599), .Y(n_856) );
O2A1O1Ixp33_ASAP7_75t_SL g857 ( .A1(n_598), .A2(n_707), .B(n_616), .C(n_641), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_649), .B(n_531), .Y(n_858) );
CKINVDCx11_ASAP7_75t_R g859 ( .A(n_719), .Y(n_859) );
OR2x2_ASAP7_75t_L g860 ( .A(n_599), .B(n_572), .Y(n_860) );
AO21x2_ASAP7_75t_L g861 ( .A1(n_669), .A2(n_682), .B(n_662), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_649), .B(n_531), .Y(n_862) );
INVx3_ASAP7_75t_L g863 ( .A(n_735), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g864 ( .A1(n_746), .A2(n_857), .B(n_833), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_787), .B(n_758), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g866 ( .A1(n_855), .A2(n_844), .B(n_846), .Y(n_866) );
OAI221xp5_ASAP7_75t_L g867 ( .A1(n_835), .A2(n_832), .B1(n_766), .B2(n_800), .C(n_862), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_788), .A2(n_860), .B1(n_754), .B2(n_818), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_853), .A2(n_859), .B1(n_851), .B2(n_858), .Y(n_869) );
INVx2_ASAP7_75t_SL g870 ( .A(n_738), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_797), .B(n_849), .Y(n_871) );
NAND2x1p5_ASAP7_75t_L g872 ( .A(n_738), .B(n_735), .Y(n_872) );
AND2x2_ASAP7_75t_L g873 ( .A(n_749), .B(n_847), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_741), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_764), .A2(n_829), .B1(n_791), .B2(n_804), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_854), .B(n_826), .Y(n_876) );
NOR2xp67_ASAP7_75t_L g877 ( .A(n_738), .B(n_753), .Y(n_877) );
AND2x2_ASAP7_75t_L g878 ( .A(n_808), .B(n_750), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_778), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_799), .A2(n_734), .B1(n_788), .B2(n_742), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_761), .A2(n_822), .B(n_809), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_729), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_770), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_808), .B(n_745), .Y(n_884) );
AND2x6_ASAP7_75t_L g885 ( .A(n_745), .B(n_852), .Y(n_885) );
OAI21xp33_ASAP7_75t_SL g886 ( .A1(n_825), .A2(n_733), .B(n_817), .Y(n_886) );
INVx1_ASAP7_75t_L g887 ( .A(n_765), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_736), .A2(n_848), .B(n_814), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_763), .B(n_771), .Y(n_889) );
BUFx2_ASAP7_75t_L g890 ( .A(n_731), .Y(n_890) );
OA21x2_ASAP7_75t_L g891 ( .A1(n_732), .A2(n_773), .B(n_748), .Y(n_891) );
AOI21xp5_ASAP7_75t_L g892 ( .A1(n_802), .A2(n_740), .B(n_861), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_815), .B(n_805), .Y(n_893) );
AOI221x1_ASAP7_75t_SL g894 ( .A1(n_772), .A2(n_783), .B1(n_836), .B2(n_838), .C(n_789), .Y(n_894) );
AND2x2_ASAP7_75t_L g895 ( .A(n_836), .B(n_780), .Y(n_895) );
AND2x4_ASAP7_75t_L g896 ( .A(n_768), .B(n_852), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_762), .A2(n_850), .B1(n_795), .B2(n_751), .Y(n_897) );
AOI21xp33_ASAP7_75t_SL g898 ( .A1(n_756), .A2(n_856), .B(n_743), .Y(n_898) );
AO21x2_ASAP7_75t_L g899 ( .A1(n_841), .A2(n_834), .B(n_728), .Y(n_899) );
BUFx12f_ASAP7_75t_L g900 ( .A(n_759), .Y(n_900) );
AOI21xp5_ASAP7_75t_L g901 ( .A1(n_843), .A2(n_839), .B(n_796), .Y(n_901) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_794), .A2(n_842), .B1(n_790), .B2(n_782), .Y(n_902) );
O2A1O1Ixp33_ASAP7_75t_L g903 ( .A1(n_775), .A2(n_840), .B(n_792), .C(n_781), .Y(n_903) );
AO22x2_ASAP7_75t_L g904 ( .A1(n_776), .A2(n_842), .B1(n_768), .B2(n_819), .Y(n_904) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_744), .A2(n_798), .B1(n_779), .B2(n_786), .C(n_821), .Y(n_905) );
OAI21xp5_ASAP7_75t_L g906 ( .A1(n_824), .A2(n_784), .B(n_767), .Y(n_906) );
AO31x2_ASAP7_75t_L g907 ( .A1(n_813), .A2(n_747), .A3(n_757), .B(n_760), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_828), .B(n_774), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_819), .B(n_831), .Y(n_909) );
INVx4_ASAP7_75t_L g910 ( .A(n_739), .Y(n_910) );
INVxp67_ASAP7_75t_L g911 ( .A(n_803), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_776), .B(n_793), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g913 ( .A1(n_823), .A2(n_811), .B1(n_816), .B2(n_801), .C(n_806), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_827), .A2(n_845), .B(n_777), .Y(n_914) );
OAI21xp5_ASAP7_75t_L g915 ( .A1(n_830), .A2(n_769), .B(n_793), .Y(n_915) );
INVxp33_ASAP7_75t_L g916 ( .A(n_785), .Y(n_916) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_785), .A2(n_828), .B1(n_755), .B2(n_837), .Y(n_917) );
INVxp67_ASAP7_75t_L g918 ( .A(n_730), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_837), .A2(n_845), .B(n_807), .Y(n_919) );
A2O1A1Ixp33_ASAP7_75t_L g920 ( .A1(n_828), .A2(n_737), .B(n_777), .C(n_730), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_730), .Y(n_921) );
INVx1_ASAP7_75t_SL g922 ( .A(n_807), .Y(n_922) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_737), .A2(n_812), .B1(n_820), .B2(n_777), .Y(n_923) );
OR2x2_ASAP7_75t_L g924 ( .A(n_737), .B(n_812), .Y(n_924) );
AO21x1_ASAP7_75t_L g925 ( .A1(n_820), .A2(n_812), .B(n_807), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_746), .A2(n_692), .B(n_690), .Y(n_926) );
OAI221xp5_ASAP7_75t_L g927 ( .A1(n_835), .A2(n_496), .B1(n_832), .B2(n_563), .C(n_766), .Y(n_927) );
OR2x6_ASAP7_75t_L g928 ( .A(n_750), .B(n_602), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_847), .Y(n_929) );
NAND2xp5_ASAP7_75t_SL g930 ( .A(n_739), .B(n_592), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_787), .B(n_636), .Y(n_931) );
BUFx3_ASAP7_75t_L g932 ( .A(n_738), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g933 ( .A1(n_849), .A2(n_702), .B1(n_653), .B2(n_651), .Y(n_933) );
BUFx8_ASAP7_75t_L g934 ( .A(n_753), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_847), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_746), .A2(n_692), .B(n_690), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_787), .B(n_636), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_847), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_746), .A2(n_692), .B(n_690), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_797), .B(n_525), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_797), .B(n_525), .Y(n_941) );
AOI21xp33_ASAP7_75t_L g942 ( .A1(n_855), .A2(n_844), .B(n_846), .Y(n_942) );
AOI21x1_ASAP7_75t_L g943 ( .A1(n_746), .A2(n_848), .B(n_736), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_797), .B(n_525), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g945 ( .A(n_810), .B(n_732), .C(n_752), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_847), .Y(n_946) );
OR2x2_ASAP7_75t_L g947 ( .A(n_787), .B(n_572), .Y(n_947) );
HB1xp67_ASAP7_75t_L g948 ( .A(n_738), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_797), .B(n_525), .Y(n_949) );
BUFx2_ASAP7_75t_L g950 ( .A(n_738), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_797), .B(n_525), .Y(n_951) );
OAI222xp33_ASAP7_75t_L g952 ( .A1(n_788), .A2(n_719), .B1(n_563), .B2(n_742), .C1(n_577), .C2(n_572), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g953 ( .A1(n_849), .A2(n_702), .B1(n_653), .B2(n_651), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_847), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_797), .B(n_525), .Y(n_955) );
NAND2xp5_ASAP7_75t_SL g956 ( .A(n_739), .B(n_592), .Y(n_956) );
INVx2_ASAP7_75t_SL g957 ( .A(n_738), .Y(n_957) );
INVx1_ASAP7_75t_L g958 ( .A(n_847), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_787), .B(n_636), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_787), .B(n_636), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_746), .A2(n_692), .B(n_690), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_847), .Y(n_962) );
AOI21x1_ASAP7_75t_L g963 ( .A1(n_746), .A2(n_848), .B(n_736), .Y(n_963) );
INVx2_ASAP7_75t_SL g964 ( .A(n_738), .Y(n_964) );
AO31x2_ASAP7_75t_L g965 ( .A1(n_732), .A2(n_669), .A3(n_746), .B(n_644), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_758), .A2(n_529), .B1(n_859), .B2(n_853), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_849), .A2(n_702), .B1(n_653), .B2(n_651), .Y(n_967) );
INVx3_ASAP7_75t_L g968 ( .A(n_735), .Y(n_968) );
CKINVDCx14_ASAP7_75t_R g969 ( .A(n_758), .Y(n_969) );
BUFx3_ASAP7_75t_L g970 ( .A(n_738), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_928), .Y(n_971) );
OA21x2_ASAP7_75t_L g972 ( .A1(n_919), .A2(n_920), .B(n_864), .Y(n_972) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_928), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_908), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_921), .Y(n_975) );
INVx2_ASAP7_75t_L g976 ( .A(n_943), .Y(n_976) );
INVx2_ASAP7_75t_L g977 ( .A(n_963), .Y(n_977) );
HB1xp67_ASAP7_75t_L g978 ( .A(n_928), .Y(n_978) );
BUFx3_ASAP7_75t_L g979 ( .A(n_872), .Y(n_979) );
INVxp67_ASAP7_75t_L g980 ( .A(n_948), .Y(n_980) );
AO21x2_ASAP7_75t_L g981 ( .A1(n_923), .A2(n_892), .B(n_925), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_924), .Y(n_982) );
OR2x2_ASAP7_75t_L g983 ( .A(n_871), .B(n_876), .Y(n_983) );
HB1xp67_ASAP7_75t_L g984 ( .A(n_950), .Y(n_984) );
AOI21x1_ASAP7_75t_L g985 ( .A1(n_923), .A2(n_881), .B(n_917), .Y(n_985) );
BUFx2_ASAP7_75t_L g986 ( .A(n_885), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_885), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_933), .B(n_953), .Y(n_988) );
AO21x2_ASAP7_75t_L g989 ( .A1(n_915), .A2(n_942), .B(n_866), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_873), .B(n_929), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_935), .B(n_938), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_879), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_918), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_880), .A2(n_867), .B1(n_927), .B2(n_933), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_953), .B(n_967), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_889), .Y(n_996) );
BUFx2_ASAP7_75t_L g997 ( .A(n_885), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_888), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_946), .B(n_954), .Y(n_999) );
BUFx2_ASAP7_75t_L g1000 ( .A(n_885), .Y(n_1000) );
INVx1_ASAP7_75t_L g1001 ( .A(n_965), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_958), .B(n_962), .Y(n_1002) );
OR2x2_ASAP7_75t_SL g1003 ( .A(n_868), .B(n_969), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_887), .B(n_882), .Y(n_1004) );
AND2x2_ASAP7_75t_L g1005 ( .A(n_883), .B(n_897), .Y(n_1005) );
INVx3_ASAP7_75t_L g1006 ( .A(n_910), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_904), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_904), .Y(n_1008) );
OA21x2_ASAP7_75t_L g1009 ( .A1(n_915), .A2(n_922), .B(n_942), .Y(n_1009) );
AND2x4_ASAP7_75t_SL g1010 ( .A(n_863), .B(n_968), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_914), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_911), .B(n_931), .Y(n_1012) );
INVx3_ASAP7_75t_L g1013 ( .A(n_910), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_937), .B(n_960), .Y(n_1014) );
INVx2_ASAP7_75t_SL g1015 ( .A(n_872), .Y(n_1015) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_952), .B(n_947), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_959), .B(n_863), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_968), .B(n_967), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_932), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_886), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_909), .B(n_884), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_886), .Y(n_1022) );
AO21x2_ASAP7_75t_L g1023 ( .A1(n_926), .A2(n_961), .B(n_936), .Y(n_1023) );
INVxp67_ASAP7_75t_L g1024 ( .A(n_877), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_880), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_939), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_970), .Y(n_1027) );
AOI21xp5_ASAP7_75t_SL g1028 ( .A1(n_905), .A2(n_891), .B(n_903), .Y(n_1028) );
OA21x2_ASAP7_75t_L g1029 ( .A1(n_945), .A2(n_901), .B(n_906), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_940), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_896), .B(n_916), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_941), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_896), .B(n_912), .Y(n_1033) );
OR2x6_ASAP7_75t_L g1034 ( .A(n_870), .B(n_964), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_899), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_944), .B(n_951), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_966), .A2(n_902), .B1(n_875), .B2(n_869), .Y(n_1037) );
OAI211xp5_ASAP7_75t_L g1038 ( .A1(n_898), .A2(n_930), .B(n_956), .C(n_949), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_955), .Y(n_1039) );
OR2x2_ASAP7_75t_L g1040 ( .A(n_957), .B(n_895), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1041 ( .A1(n_865), .A2(n_945), .B1(n_878), .B2(n_893), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_890), .B(n_907), .Y(n_1042) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_907), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_907), .B(n_894), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_913), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_874), .B(n_934), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_998), .Y(n_1047) );
BUFx3_ASAP7_75t_L g1048 ( .A(n_979), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_988), .B(n_934), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_988), .B(n_900), .Y(n_1050) );
BUFx3_ASAP7_75t_L g1051 ( .A(n_979), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1020), .B(n_1022), .Y(n_1052) );
HB1xp67_ASAP7_75t_L g1053 ( .A(n_974), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_975), .Y(n_1054) );
OR2x2_ASAP7_75t_L g1055 ( .A(n_995), .B(n_1042), .Y(n_1055) );
INVx4_ASAP7_75t_L g1056 ( .A(n_986), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1020), .B(n_1022), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1058 ( .A1(n_994), .A2(n_1016), .B1(n_1025), .B2(n_995), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_974), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1060 ( .A(n_982), .B(n_1044), .Y(n_1060) );
AOI33xp33_ASAP7_75t_L g1061 ( .A1(n_1004), .A2(n_991), .A3(n_1002), .B1(n_1005), .B2(n_1014), .B3(n_1012), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_982), .B(n_1044), .Y(n_1062) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_1037), .A2(n_990), .B1(n_1018), .B2(n_1005), .Y(n_1063) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_993), .Y(n_1064) );
AND2x2_ASAP7_75t_L g1065 ( .A(n_989), .B(n_1043), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_993), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_989), .B(n_1043), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_989), .B(n_1001), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1001), .B(n_1026), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_1042), .B(n_983), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1023), .B(n_981), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_1018), .Y(n_1072) );
OR2x2_ASAP7_75t_L g1073 ( .A(n_983), .B(n_1007), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_981), .B(n_1011), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_1008), .Y(n_1075) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_1003), .B(n_1041), .Y(n_1076) );
BUFx2_ASAP7_75t_L g1077 ( .A(n_986), .Y(n_1077) );
OR2x2_ASAP7_75t_L g1078 ( .A(n_1003), .B(n_1041), .Y(n_1078) );
INVx2_ASAP7_75t_SL g1079 ( .A(n_1010), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_992), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_992), .Y(n_1081) );
AO21x2_ASAP7_75t_L g1082 ( .A1(n_1028), .A2(n_977), .B(n_976), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_987), .Y(n_1083) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_987), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_997), .A2(n_1000), .B1(n_996), .B2(n_973), .Y(n_1085) );
NOR2x1_ASAP7_75t_SL g1086 ( .A(n_979), .B(n_1015), .Y(n_1086) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1054), .Y(n_1087) );
NAND2xp5_ASAP7_75t_SL g1088 ( .A(n_1079), .B(n_1015), .Y(n_1088) );
NAND2xp5_ASAP7_75t_L g1089 ( .A(n_1061), .B(n_1004), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1054), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1052), .B(n_1057), .Y(n_1091) );
OR2x2_ASAP7_75t_L g1092 ( .A(n_1070), .B(n_1014), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1047), .Y(n_1093) );
HB1xp67_ASAP7_75t_L g1094 ( .A(n_1053), .Y(n_1094) );
INVx1_ASAP7_75t_SL g1095 ( .A(n_1048), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1072), .B(n_1009), .Y(n_1096) );
AND2x2_ASAP7_75t_L g1097 ( .A(n_1072), .B(n_1009), .Y(n_1097) );
INVx2_ASAP7_75t_SL g1098 ( .A(n_1048), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1099 ( .A(n_1049), .B(n_1046), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_1063), .B(n_991), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1060), .B(n_1009), .Y(n_1101) );
OR2x2_ASAP7_75t_L g1102 ( .A(n_1070), .B(n_1012), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1103 ( .A(n_1053), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_1060), .B(n_1009), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1058), .B(n_1002), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_1060), .B(n_972), .Y(n_1106) );
INVx1_ASAP7_75t_SL g1107 ( .A(n_1048), .Y(n_1107) );
NAND2xp5_ASAP7_75t_SL g1108 ( .A(n_1079), .B(n_997), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1062), .B(n_972), .Y(n_1109) );
INVxp67_ASAP7_75t_L g1110 ( .A(n_1049), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1111 ( .A(n_1070), .B(n_972), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1062), .B(n_972), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1113 ( .A(n_1055), .B(n_1029), .Y(n_1113) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_1076), .A2(n_1000), .B1(n_971), .B2(n_978), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1062), .B(n_985), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1058), .B(n_1032), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1080), .B(n_1032), .Y(n_1117) );
NAND2x1p5_ASAP7_75t_L g1118 ( .A(n_1051), .B(n_1079), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1074), .B(n_1029), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1081), .B(n_1030), .Y(n_1120) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1074), .B(n_1029), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1081), .B(n_1039), .Y(n_1122) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_1069), .B(n_1029), .Y(n_1123) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_1055), .B(n_1035), .Y(n_1124) );
INVxp67_ASAP7_75t_L g1125 ( .A(n_1049), .Y(n_1125) );
INVx3_ASAP7_75t_L g1126 ( .A(n_1082), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1127 ( .A(n_1050), .B(n_1046), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1087), .Y(n_1128) );
NOR2x1_ASAP7_75t_L g1129 ( .A(n_1099), .B(n_1051), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_1091), .B(n_1055), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_1110), .B(n_1050), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1091), .B(n_1065), .Y(n_1132) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1116), .B(n_1073), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_1105), .B(n_1073), .Y(n_1134) );
INVx1_ASAP7_75t_SL g1135 ( .A(n_1092), .Y(n_1135) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_1098), .Y(n_1136) );
OR2x6_ASAP7_75t_SL g1137 ( .A(n_1092), .B(n_1076), .Y(n_1137) );
NOR2x1p5_ASAP7_75t_SL g1138 ( .A(n_1113), .B(n_1076), .Y(n_1138) );
INVx2_ASAP7_75t_SL g1139 ( .A(n_1098), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1093), .Y(n_1140) );
OR2x2_ASAP7_75t_L g1141 ( .A(n_1102), .B(n_1073), .Y(n_1141) );
OR2x2_ASAP7_75t_L g1142 ( .A(n_1111), .B(n_1059), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1089), .B(n_1059), .Y(n_1143) );
OAI21xp33_ASAP7_75t_L g1144 ( .A1(n_1127), .A2(n_1078), .B(n_1071), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1106), .B(n_1065), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1087), .Y(n_1146) );
INVxp67_ASAP7_75t_L g1147 ( .A(n_1094), .Y(n_1147) );
OR2x2_ASAP7_75t_L g1148 ( .A(n_1102), .B(n_1064), .Y(n_1148) );
HB1xp67_ASAP7_75t_L g1149 ( .A(n_1103), .Y(n_1149) );
NOR2xp67_ASAP7_75t_L g1150 ( .A(n_1125), .B(n_1078), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1100), .B(n_1064), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1152 ( .A(n_1111), .B(n_1075), .Y(n_1152) );
NAND4xp25_ASAP7_75t_SL g1153 ( .A(n_1107), .B(n_1078), .C(n_1050), .D(n_1038), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1106), .B(n_1065), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_1114), .A2(n_1085), .B1(n_1017), .B2(n_1036), .Y(n_1155) );
INVx1_ASAP7_75t_SL g1156 ( .A(n_1095), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1109), .B(n_1067), .Y(n_1157) );
INVx1_ASAP7_75t_SL g1158 ( .A(n_1107), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1109), .B(n_1067), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1090), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1161 ( .A(n_1123), .B(n_1067), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1112), .B(n_1068), .Y(n_1162) );
INVxp67_ASAP7_75t_L g1163 ( .A(n_1117), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1113), .B(n_1075), .Y(n_1164) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_1124), .B(n_1066), .Y(n_1165) );
AND2x2_ASAP7_75t_SL g1166 ( .A(n_1096), .B(n_1056), .Y(n_1166) );
INVx3_ASAP7_75t_SL g1167 ( .A(n_1088), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1168 ( .A(n_1143), .B(n_1123), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1162), .B(n_1119), .Y(n_1169) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1135), .B(n_1119), .Y(n_1170) );
NAND2xp5_ASAP7_75t_SL g1171 ( .A(n_1166), .B(n_1118), .Y(n_1171) );
CKINVDCx16_ASAP7_75t_R g1172 ( .A(n_1137), .Y(n_1172) );
INVx1_ASAP7_75t_SL g1173 ( .A(n_1156), .Y(n_1173) );
NOR2xp67_ASAP7_75t_SL g1174 ( .A(n_1136), .B(n_1051), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1140), .Y(n_1175) );
INVxp33_ASAP7_75t_L g1176 ( .A(n_1129), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1177 ( .A(n_1130), .B(n_1121), .Y(n_1177) );
NAND2xp5_ASAP7_75t_L g1178 ( .A(n_1163), .B(n_1121), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1179 ( .A(n_1130), .B(n_1124), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1162), .B(n_1112), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1164), .Y(n_1181) );
INVxp67_ASAP7_75t_L g1182 ( .A(n_1149), .Y(n_1182) );
NAND2xp5_ASAP7_75t_SL g1183 ( .A(n_1166), .B(n_1118), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1151), .B(n_1101), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_1132), .B(n_1101), .Y(n_1185) );
NOR2xp33_ASAP7_75t_L g1186 ( .A(n_1131), .B(n_1024), .Y(n_1186) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1164), .Y(n_1187) );
NAND2x1p5_ASAP7_75t_L g1188 ( .A(n_1136), .B(n_1056), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1161), .B(n_1104), .Y(n_1189) );
NOR2xp33_ASAP7_75t_L g1190 ( .A(n_1131), .B(n_1019), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1128), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1146), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1160), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1194 ( .A(n_1132), .B(n_1104), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1195 ( .A(n_1147), .B(n_1027), .Y(n_1195) );
AOI21xp5_ASAP7_75t_L g1196 ( .A1(n_1171), .A2(n_1153), .B(n_1139), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1197 ( .A1(n_1183), .A2(n_1139), .B(n_1108), .Y(n_1197) );
AND2x4_ASAP7_75t_L g1198 ( .A(n_1181), .B(n_1138), .Y(n_1198) );
OAI222xp33_ASAP7_75t_L g1199 ( .A1(n_1172), .A2(n_1155), .B1(n_1148), .B2(n_1137), .C1(n_1141), .C2(n_1158), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1181), .Y(n_1200) );
INVxp67_ASAP7_75t_L g1201 ( .A(n_1173), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1187), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1189), .B(n_1161), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1187), .Y(n_1204) );
AND2x4_ASAP7_75t_L g1205 ( .A(n_1189), .B(n_1161), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1179), .Y(n_1206) );
AOI22xp5_ASAP7_75t_L g1207 ( .A1(n_1172), .A2(n_1144), .B1(n_1150), .B2(n_1134), .Y(n_1207) );
CKINVDCx16_ASAP7_75t_R g1208 ( .A(n_1190), .Y(n_1208) );
OAI31xp33_ASAP7_75t_L g1209 ( .A1(n_1176), .A2(n_1085), .A3(n_1118), .B(n_1142), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_1188), .A2(n_1167), .B1(n_1056), .B2(n_1142), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1169), .B(n_1145), .Y(n_1211) );
OAI21xp33_ASAP7_75t_L g1212 ( .A1(n_1168), .A2(n_1159), .B(n_1157), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1178), .B(n_1145), .Y(n_1213) );
INVx2_ASAP7_75t_L g1214 ( .A(n_1175), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_1186), .A2(n_1017), .B1(n_1021), .B2(n_1115), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1179), .Y(n_1216) );
AOI322xp5_ASAP7_75t_L g1217 ( .A1(n_1212), .A2(n_1169), .A3(n_1180), .B1(n_1195), .B2(n_1194), .C1(n_1185), .C2(n_1182), .Y(n_1217) );
AOI21xp5_ASAP7_75t_L g1218 ( .A1(n_1199), .A2(n_1188), .B(n_1086), .Y(n_1218) );
OAI22xp33_ASAP7_75t_L g1219 ( .A1(n_1207), .A2(n_1167), .B1(n_1188), .B2(n_1177), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1206), .B(n_1177), .Y(n_1220) );
OAI221xp5_ASAP7_75t_L g1221 ( .A1(n_1209), .A2(n_1133), .B1(n_1170), .B2(n_1184), .C(n_1174), .Y(n_1221) );
AOI322xp5_ASAP7_75t_L g1222 ( .A1(n_1208), .A2(n_1180), .A3(n_1154), .B1(n_1157), .B2(n_1159), .C1(n_1097), .C2(n_1096), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1200), .Y(n_1223) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1214), .Y(n_1224) );
OAI211xp5_ASAP7_75t_L g1225 ( .A1(n_1196), .A2(n_1056), .B(n_1152), .C(n_980), .Y(n_1225) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1202), .Y(n_1226) );
NAND2xp5_ASAP7_75t_SL g1227 ( .A(n_1198), .B(n_1175), .Y(n_1227) );
OAI22xp5_ASAP7_75t_SL g1228 ( .A1(n_1201), .A2(n_1056), .B1(n_1084), .B2(n_1077), .Y(n_1228) );
OAI21xp5_ASAP7_75t_SL g1229 ( .A1(n_1210), .A2(n_1010), .B(n_1083), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1230 ( .A1(n_1215), .A2(n_1154), .B1(n_1174), .B2(n_1191), .Y(n_1230) );
AOI22xp5_ASAP7_75t_L g1231 ( .A1(n_1225), .A2(n_1198), .B1(n_1215), .B2(n_1216), .Y(n_1231) );
NAND2xp33_ASAP7_75t_R g1232 ( .A(n_1218), .B(n_1198), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1217), .B(n_1204), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_1221), .A2(n_1205), .B1(n_1203), .B2(n_1211), .Y(n_1234) );
AOI311xp33_ASAP7_75t_L g1235 ( .A1(n_1219), .A2(n_1197), .A3(n_1213), .B(n_1192), .C(n_1193), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_1228), .A2(n_1205), .B1(n_1115), .B2(n_1203), .Y(n_1236) );
NOR2x1_ASAP7_75t_L g1237 ( .A(n_1229), .B(n_1205), .Y(n_1237) );
OAI22xp5_ASAP7_75t_L g1238 ( .A1(n_1229), .A2(n_1211), .B1(n_1214), .B2(n_1165), .Y(n_1238) );
INVxp67_ASAP7_75t_L g1239 ( .A(n_1230), .Y(n_1239) );
NOR3xp33_ASAP7_75t_L g1240 ( .A(n_1233), .B(n_1227), .C(n_1039), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1239), .Y(n_1241) );
NAND4xp75_ASAP7_75t_L g1242 ( .A(n_1237), .B(n_1226), .C(n_1223), .D(n_999), .Y(n_1242) );
XOR2x2_ASAP7_75t_L g1243 ( .A(n_1234), .B(n_1220), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_1238), .A2(n_1224), .B1(n_1191), .B2(n_1193), .C(n_1192), .Y(n_1244) );
NAND3xp33_ASAP7_75t_L g1245 ( .A(n_1235), .B(n_1222), .C(n_984), .Y(n_1245) );
NOR2x1_ASAP7_75t_L g1246 ( .A(n_1232), .B(n_1034), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_1245), .A2(n_1236), .B1(n_1231), .B2(n_1083), .C(n_1077), .Y(n_1247) );
NAND2xp5_ASAP7_75t_SL g1248 ( .A(n_1246), .B(n_1126), .Y(n_1248) );
AND3x2_ASAP7_75t_L g1249 ( .A(n_1241), .B(n_1084), .C(n_1036), .Y(n_1249) );
OAI22xp5_ASAP7_75t_SL g1250 ( .A1(n_1242), .A2(n_1034), .B1(n_1040), .B2(n_1006), .Y(n_1250) );
NOR3xp33_ASAP7_75t_L g1251 ( .A(n_1240), .B(n_1013), .C(n_1006), .Y(n_1251) );
NAND5xp2_ASAP7_75t_L g1252 ( .A(n_1247), .B(n_1244), .C(n_1243), .D(n_1045), .E(n_1031), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1249), .Y(n_1253) );
INVx3_ASAP7_75t_L g1254 ( .A(n_1248), .Y(n_1254) );
NAND3xp33_ASAP7_75t_L g1255 ( .A(n_1251), .B(n_1034), .C(n_1040), .Y(n_1255) );
INVx2_ASAP7_75t_L g1256 ( .A(n_1254), .Y(n_1256) );
BUFx6f_ASAP7_75t_L g1257 ( .A(n_1253), .Y(n_1257) );
OAI21xp5_ASAP7_75t_SL g1258 ( .A1(n_1255), .A2(n_1250), .B(n_1010), .Y(n_1258) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1257), .Y(n_1259) );
INVx1_ASAP7_75t_SL g1260 ( .A(n_1257), .Y(n_1260) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1256), .Y(n_1261) );
OAI21x1_ASAP7_75t_L g1262 ( .A1(n_1259), .A2(n_1254), .B(n_1258), .Y(n_1262) );
XNOR2xp5_ASAP7_75t_L g1263 ( .A(n_1260), .B(n_1252), .Y(n_1263) );
OAI222xp33_ASAP7_75t_L g1264 ( .A1(n_1263), .A2(n_1261), .B1(n_1259), .B2(n_1034), .C1(n_996), .C2(n_1033), .Y(n_1264) );
OA21x2_ASAP7_75t_L g1265 ( .A1(n_1262), .A2(n_1122), .B(n_1120), .Y(n_1265) );
AOI21xp5_ASAP7_75t_L g1266 ( .A1(n_1264), .A2(n_1262), .B(n_1034), .Y(n_1266) );
AOI22xp5_ASAP7_75t_L g1267 ( .A1(n_1266), .A2(n_1265), .B1(n_1033), .B2(n_1021), .Y(n_1267) );
endmodule