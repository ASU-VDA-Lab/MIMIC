module real_aes_1516_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_782, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_782;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_0), .B(n_125), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_1), .A2(n_134), .B(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_2), .B(n_778), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_3), .B(n_125), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_4), .B(n_141), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_5), .B(n_141), .Y(n_480) );
INVx1_ASAP7_75t_L g132 ( .A(n_6), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_7), .B(n_141), .Y(n_550) );
CKINVDCx16_ASAP7_75t_R g778 ( .A(n_8), .Y(n_778) );
NAND2xp33_ASAP7_75t_L g535 ( .A(n_9), .B(n_143), .Y(n_535) );
AND2x2_ASAP7_75t_L g161 ( .A(n_10), .B(n_150), .Y(n_161) );
AND2x2_ASAP7_75t_L g172 ( .A(n_11), .B(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
AOI221x1_ASAP7_75t_L g484 ( .A1(n_13), .A2(n_24), .B1(n_125), .B2(n_134), .C(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_14), .B(n_141), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_15), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_16), .B(n_125), .Y(n_531) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_17), .A2(n_150), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_18), .B(n_145), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_19), .B(n_141), .Y(n_524) );
AO21x1_ASAP7_75t_L g475 ( .A1(n_20), .A2(n_125), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_21), .B(n_125), .Y(n_229) );
INVx1_ASAP7_75t_L g451 ( .A(n_22), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_23), .A2(n_91), .B1(n_125), .B2(n_178), .Y(n_177) );
NAND2x1_ASAP7_75t_L g495 ( .A(n_25), .B(n_141), .Y(n_495) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_26), .B(n_143), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_27), .Y(n_457) );
OR2x2_ASAP7_75t_L g148 ( .A(n_28), .B(n_88), .Y(n_148) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_28), .A2(n_88), .B(n_147), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_29), .B(n_143), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_30), .B(n_141), .Y(n_534) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_31), .A2(n_173), .B(n_220), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_32), .A2(n_105), .B1(n_772), .B2(n_779), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_33), .B(n_143), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_34), .A2(n_134), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_35), .B(n_141), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_36), .A2(n_134), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g131 ( .A(n_37), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g135 ( .A(n_37), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g186 ( .A(n_37), .Y(n_186) );
OR2x6_ASAP7_75t_L g449 ( .A(n_38), .B(n_450), .Y(n_449) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_38), .B(n_447), .C(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_39), .B(n_125), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_40), .B(n_125), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_41), .B(n_141), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_42), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_43), .B(n_143), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_44), .B(n_125), .Y(n_124) );
AOI22xp5_ASAP7_75t_SL g463 ( .A1(n_45), .A2(n_67), .B1(n_464), .B2(n_465), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_45), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_46), .A2(n_86), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_46), .Y(n_437) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_47), .A2(n_134), .B(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_48), .A2(n_134), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_49), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_50), .B(n_143), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_51), .B(n_125), .Y(n_221) );
XNOR2xp5_ASAP7_75t_L g462 ( .A(n_52), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g128 ( .A(n_53), .Y(n_128) );
INVx1_ASAP7_75t_L g138 ( .A(n_53), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_54), .B(n_141), .Y(n_170) );
AND2x2_ASAP7_75t_L g210 ( .A(n_55), .B(n_145), .Y(n_210) );
XOR2xp5_ASAP7_75t_L g461 ( .A(n_56), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_57), .B(n_143), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_58), .B(n_141), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_59), .B(n_143), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_60), .A2(n_134), .B(n_494), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_61), .B(n_125), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_62), .B(n_125), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_63), .A2(n_134), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g235 ( .A(n_64), .B(n_146), .Y(n_235) );
AO21x1_ASAP7_75t_L g477 ( .A1(n_65), .A2(n_134), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_66), .B(n_125), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_67), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_68), .B(n_143), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_69), .B(n_125), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_70), .B(n_143), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_71), .A2(n_95), .B1(n_134), .B2(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_72), .B(n_141), .Y(n_232) );
AND2x2_ASAP7_75t_L g508 ( .A(n_73), .B(n_146), .Y(n_508) );
INVx1_ASAP7_75t_L g130 ( .A(n_74), .Y(n_130) );
INVx1_ASAP7_75t_L g136 ( .A(n_74), .Y(n_136) );
AND2x2_ASAP7_75t_L g552 ( .A(n_75), .B(n_173), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_76), .B(n_143), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_77), .A2(n_134), .B(n_214), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_78), .A2(n_134), .B(n_139), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_79), .A2(n_134), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g246 ( .A(n_80), .B(n_146), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_81), .B(n_145), .Y(n_175) );
INVx1_ASAP7_75t_L g452 ( .A(n_82), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_82), .B(n_451), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_83), .B(n_125), .Y(n_526) );
AND2x2_ASAP7_75t_L g538 ( .A(n_84), .B(n_173), .Y(n_538) );
AND2x2_ASAP7_75t_L g149 ( .A(n_85), .B(n_150), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_86), .Y(n_436) );
AND2x2_ASAP7_75t_L g476 ( .A(n_87), .B(n_217), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_89), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_89), .B(n_112), .C(n_442), .Y(n_454) );
AND2x2_ASAP7_75t_L g498 ( .A(n_89), .B(n_173), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_90), .B(n_143), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_92), .B(n_141), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_93), .B(n_143), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_94), .A2(n_134), .B(n_523), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_96), .A2(n_134), .B(n_231), .Y(n_230) );
OAI22xp5_ASAP7_75t_SL g433 ( .A1(n_97), .A2(n_434), .B1(n_435), .B2(n_438), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_97), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_98), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_99), .B(n_141), .Y(n_543) );
BUFx2_ASAP7_75t_L g234 ( .A(n_100), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_101), .A2(n_449), .B1(n_460), .B2(n_767), .Y(n_459) );
BUFx2_ASAP7_75t_L g110 ( .A(n_102), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_103), .A2(n_134), .B(n_533), .Y(n_532) );
OA21x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_458), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_108), .B(n_456), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
OAI211xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_441), .B(n_454), .C(n_455), .Y(n_111) );
AOI22x1_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_433), .B1(n_439), .B2(n_440), .Y(n_112) );
INVx3_ASAP7_75t_L g440 ( .A(n_113), .Y(n_440) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_113), .A2(n_467), .B1(n_765), .B2(n_766), .Y(n_466) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_346), .Y(n_113) );
NOR4xp75_ASAP7_75t_L g114 ( .A(n_115), .B(n_269), .C(n_294), .D(n_321), .Y(n_114) );
OAI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_205), .B(n_247), .Y(n_115) );
NOR4xp25_ASAP7_75t_L g116 ( .A(n_117), .B(n_189), .C(n_196), .D(n_200), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_162), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_152), .Y(n_120) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_121), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_121), .B(n_193), .Y(n_340) );
AND2x2_ASAP7_75t_L g365 ( .A(n_121), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g390 ( .A(n_121), .B(n_174), .Y(n_390) );
AND2x2_ASAP7_75t_L g431 ( .A(n_121), .B(n_198), .Y(n_431) );
INVx4_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_SL g202 ( .A(n_122), .B(n_195), .Y(n_202) );
AND2x2_ASAP7_75t_L g204 ( .A(n_122), .B(n_164), .Y(n_204) );
NOR2x1_ASAP7_75t_L g255 ( .A(n_122), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g266 ( .A(n_122), .Y(n_266) );
AND2x2_ASAP7_75t_L g272 ( .A(n_122), .B(n_198), .Y(n_272) );
BUFx2_ASAP7_75t_L g285 ( .A(n_122), .Y(n_285) );
AND2x4_ASAP7_75t_L g316 ( .A(n_122), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g363 ( .A(n_122), .B(n_364), .Y(n_363) );
OR2x6_ASAP7_75t_L g122 ( .A(n_123), .B(n_149), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_133), .B(n_145), .Y(n_123) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_131), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_127), .B(n_129), .Y(n_126) );
AND2x6_ASAP7_75t_L g143 ( .A(n_127), .B(n_136), .Y(n_143) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g141 ( .A(n_129), .B(n_138), .Y(n_141) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx5_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
AND2x2_ASAP7_75t_L g137 ( .A(n_132), .B(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
AND2x6_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
BUFx3_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
INVx2_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
AND2x4_ASAP7_75t_L g184 ( .A(n_137), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g180 ( .A(n_138), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_142), .B(n_144), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_143), .B(n_234), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_144), .A2(n_158), .B(n_159), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_144), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_144), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_144), .A2(n_224), .B(n_225), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_144), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_144), .A2(n_243), .B(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_144), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_144), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_144), .A2(n_495), .B(n_496), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_144), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_144), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_144), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_144), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_144), .A2(n_549), .B(n_550), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_145), .Y(n_154) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_145), .A2(n_177), .B(n_183), .Y(n_176) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_145), .A2(n_484), .B(n_488), .Y(n_483) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_145), .A2(n_484), .B(n_488), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_145), .A2(n_540), .B(n_541), .Y(n_539) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_147), .B(n_148), .Y(n_146) );
AND2x4_ASAP7_75t_L g217 ( .A(n_147), .B(n_148), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_150), .A2(n_229), .B(n_230), .Y(n_228) );
BUFx4f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
INVx1_ASAP7_75t_L g357 ( .A(n_152), .Y(n_357) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
AND2x2_ASAP7_75t_L g198 ( .A(n_153), .B(n_164), .Y(n_198) );
AOI21x1_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_161), .Y(n_153) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_154), .A2(n_546), .B(n_552), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_162), .B(n_375), .Y(n_428) );
INVx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g265 ( .A(n_163), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_174), .Y(n_163) );
INVx2_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
INVx2_ASAP7_75t_L g256 ( .A(n_164), .Y(n_256) );
AND2x2_ASAP7_75t_L g366 ( .A(n_164), .B(n_195), .Y(n_366) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_172), .Y(n_164) );
INVx4_ASAP7_75t_L g173 ( .A(n_165), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
INVx3_ASAP7_75t_L g239 ( .A(n_173), .Y(n_239) );
INVx2_ASAP7_75t_L g254 ( .A(n_174), .Y(n_254) );
BUFx3_ASAP7_75t_L g271 ( .A(n_174), .Y(n_271) );
AND2x2_ASAP7_75t_L g298 ( .A(n_174), .B(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AND2x4_ASAP7_75t_L g191 ( .A(n_175), .B(n_176), .Y(n_191) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_182), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2x1p5_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NOR2x1_ASAP7_75t_L g189 ( .A(n_190), .B(n_192), .Y(n_189) );
INVx2_ASAP7_75t_L g199 ( .A(n_190), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_190), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g369 ( .A(n_190), .B(n_309), .Y(n_369) );
AND2x2_ASAP7_75t_L g393 ( .A(n_190), .B(n_202), .Y(n_393) );
INVx3_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g289 ( .A(n_191), .B(n_194), .Y(n_289) );
AND2x2_ASAP7_75t_L g371 ( .A(n_191), .B(n_364), .Y(n_371) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_SL g414 ( .A(n_193), .Y(n_414) );
AND2x2_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g299 ( .A(n_194), .Y(n_299) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_195), .Y(n_303) );
INVx2_ASAP7_75t_L g311 ( .A(n_195), .Y(n_311) );
INVx1_ASAP7_75t_L g317 ( .A(n_195), .Y(n_317) );
AOI222xp33_ASAP7_75t_SL g247 ( .A1(n_196), .A2(n_248), .B1(n_252), .B2(n_257), .C1(n_264), .C2(n_267), .Y(n_247) );
INVx1_ASAP7_75t_SL g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g324 ( .A(n_198), .Y(n_324) );
BUFx2_ASAP7_75t_L g353 ( .A(n_198), .Y(n_353) );
OAI211xp5_ASAP7_75t_L g347 ( .A1(n_199), .A2(n_348), .B(n_352), .C(n_360), .Y(n_347) );
OR2x2_ASAP7_75t_L g418 ( .A(n_199), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g426 ( .A(n_199), .B(n_331), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_203), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_202), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g401 ( .A(n_202), .B(n_289), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_202), .B(n_381), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_203), .B(n_271), .Y(n_409) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g331 ( .A(n_204), .B(n_303), .Y(n_331) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_226), .Y(n_206) );
INVx1_ASAP7_75t_L g425 ( .A(n_207), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AND2x2_ASAP7_75t_L g268 ( .A(n_208), .B(n_227), .Y(n_268) );
INVx1_ASAP7_75t_L g345 ( .A(n_208), .Y(n_345) );
OR2x2_ASAP7_75t_L g404 ( .A(n_208), .B(n_227), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_208), .B(n_276), .Y(n_410) );
INVx4_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
OR2x2_ASAP7_75t_L g283 ( .A(n_209), .B(n_237), .Y(n_283) );
AND2x2_ASAP7_75t_L g292 ( .A(n_209), .B(n_219), .Y(n_292) );
NAND2x1_ASAP7_75t_L g320 ( .A(n_209), .B(n_227), .Y(n_320) );
AND2x2_ASAP7_75t_L g367 ( .A(n_209), .B(n_262), .Y(n_367) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_217), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_217), .A2(n_221), .B(n_222), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_217), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g520 ( .A(n_217), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_217), .A2(n_531), .B(n_532), .Y(n_530) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
INVx1_ASAP7_75t_L g260 ( .A(n_219), .Y(n_260) );
AND2x2_ASAP7_75t_L g276 ( .A(n_219), .B(n_263), .Y(n_276) );
INVx2_ASAP7_75t_L g281 ( .A(n_219), .Y(n_281) );
OR2x2_ASAP7_75t_L g377 ( .A(n_219), .B(n_227), .Y(n_377) );
AND2x2_ASAP7_75t_L g226 ( .A(n_227), .B(n_236), .Y(n_226) );
NOR2x1_ASAP7_75t_SL g262 ( .A(n_227), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g280 ( .A(n_227), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g293 ( .A(n_227), .B(n_237), .Y(n_293) );
BUFx2_ASAP7_75t_L g312 ( .A(n_227), .Y(n_312) );
INVx2_ASAP7_75t_SL g339 ( .A(n_227), .Y(n_339) );
OR2x6_ASAP7_75t_L g227 ( .A(n_228), .B(n_235), .Y(n_227) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g249 ( .A(n_237), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g395 ( .A(n_237), .B(n_337), .Y(n_395) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_246), .Y(n_238) );
AO21x1_ASAP7_75t_SL g263 ( .A1(n_239), .A2(n_240), .B(n_246), .Y(n_263) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_239), .A2(n_492), .B(n_498), .Y(n_491) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_239), .A2(n_502), .B(n_508), .Y(n_501) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_239), .A2(n_492), .B(n_498), .Y(n_513) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_239), .A2(n_502), .B(n_508), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_245), .Y(n_240) );
AOI211xp5_ASAP7_75t_L g411 ( .A1(n_248), .A2(n_272), .B(n_412), .C(n_416), .Y(n_411) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_249), .B(n_327), .Y(n_362) );
BUFx2_ASAP7_75t_L g326 ( .A(n_250), .Y(n_326) );
OR2x2_ASAP7_75t_L g274 ( .A(n_251), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g359 ( .A(n_251), .B(n_293), .Y(n_359) );
AND2x2_ASAP7_75t_L g380 ( .A(n_251), .B(n_336), .Y(n_380) );
INVx2_ASAP7_75t_L g387 ( .A(n_251), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g392 ( .A1(n_252), .A2(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g334 ( .A(n_253), .B(n_316), .Y(n_334) );
OR2x2_ASAP7_75t_L g413 ( .A(n_253), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_254), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_256), .Y(n_287) );
AND2x2_ASAP7_75t_L g364 ( .A(n_256), .B(n_311), .Y(n_364) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
AND2x2_ASAP7_75t_L g349 ( .A(n_259), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_SL g358 ( .A(n_259), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_259), .B(n_268), .Y(n_391) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g267 ( .A(n_260), .B(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g386 ( .A(n_261), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g336 ( .A(n_262), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g306 ( .A(n_263), .B(n_281), .Y(n_306) );
OAI31xp33_ASAP7_75t_L g313 ( .A1(n_264), .A2(n_314), .A3(n_316), .B(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_266), .B(n_289), .Y(n_315) );
AO21x1_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_273), .B(n_277), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
OR2x2_ASAP7_75t_L g325 ( .A(n_271), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g430 ( .A(n_271), .Y(n_430) );
INVx2_ASAP7_75t_SL g415 ( .A(n_272), .Y(n_415) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g319 ( .A(n_275), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g403 ( .A(n_275), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_276), .B(n_339), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_284), .B1(n_288), .B2(n_290), .Y(n_277) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_278), .A2(n_397), .B(n_398), .Y(n_396) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_L g337 ( .A(n_281), .Y(n_337) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g351 ( .A(n_283), .B(n_312), .Y(n_351) );
OR2x2_ASAP7_75t_L g376 ( .A(n_283), .B(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_285), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_285), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g375 ( .A(n_285), .Y(n_375) );
INVx2_ASAP7_75t_L g304 ( .A(n_286), .Y(n_304) );
INVx1_ASAP7_75t_L g384 ( .A(n_287), .Y(n_384) );
AND2x2_ASAP7_75t_L g307 ( .A(n_289), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g381 ( .A(n_289), .Y(n_381) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_295), .B(n_313), .Y(n_294) );
OAI321xp33_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .A3(n_305), .B1(n_306), .B2(n_307), .C(n_312), .Y(n_295) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_296), .A2(n_327), .A3(n_422), .B1(n_424), .B2(n_426), .C1(n_427), .C2(n_432), .Y(n_421) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g374 ( .A(n_299), .Y(n_374) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_301), .B(n_381), .Y(n_398) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g406 ( .A(n_304), .Y(n_406) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp33_ASAP7_75t_SL g338 ( .A(n_306), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI21xp33_ASAP7_75t_SL g405 ( .A1(n_309), .A2(n_315), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx3_ASAP7_75t_L g327 ( .A(n_320), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_341), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_327), .B1(n_328), .B2(n_329), .C(n_332), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
AND2x2_ASAP7_75t_L g328 ( .A(n_326), .B(n_327), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI22xp33_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_335), .B1(n_338), .B2(n_340), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g344 ( .A(n_336), .B(n_345), .Y(n_344) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_339), .A2(n_428), .B(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NOR3xp33_ASAP7_75t_SL g346 ( .A(n_347), .B(n_378), .C(n_399), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_351), .A2(n_386), .B1(n_413), .B2(n_415), .Y(n_412) );
OAI21xp33_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_354), .B(n_358), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_353), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_359), .A2(n_401), .B1(n_402), .B2(n_405), .C(n_407), .Y(n_400) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B1(n_365), .B2(n_367), .C(n_368), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g397 ( .A(n_363), .Y(n_397) );
INVx1_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
INVx1_ASAP7_75t_SL g417 ( .A(n_365), .Y(n_417) );
AOI31xp33_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .A3(n_372), .B(n_376), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_369), .A2(n_379), .B1(n_381), .B2(n_382), .C(n_782), .Y(n_378) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI211xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .B(n_388), .C(n_396), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g394 ( .A(n_387), .B(n_395), .Y(n_394) );
OAI21xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_391), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g423 ( .A(n_395), .Y(n_423) );
BUFx2_ASAP7_75t_SL g432 ( .A(n_395), .Y(n_432) );
NAND3xp33_ASAP7_75t_SL g399 ( .A(n_400), .B(n_411), .C(n_421), .Y(n_399) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B(n_410), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_420), .Y(n_416) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g439 ( .A(n_433), .Y(n_439) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_442), .B(n_453), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_444), .B(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
CKINVDCx16_ASAP7_75t_R g766 ( .A(n_447), .Y(n_766) );
OR2x2_ASAP7_75t_L g770 ( .A(n_447), .B(n_449), .Y(n_770) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_771), .Y(n_458) );
XNOR2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_466), .Y(n_460) );
AND2x4_ASAP7_75t_L g467 ( .A(n_468), .B(n_664), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_601), .C(n_624), .Y(n_468) );
NAND3xp33_ASAP7_75t_SL g469 ( .A(n_470), .B(n_553), .C(n_570), .Y(n_469) );
OAI31xp33_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_489), .A3(n_509), .B(n_516), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_471), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_483), .Y(n_472) );
AND2x4_ASAP7_75t_L g556 ( .A(n_473), .B(n_483), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_473), .B(n_500), .Y(n_585) );
AND2x4_ASAP7_75t_L g587 ( .A(n_473), .B(n_581), .Y(n_587) );
AND2x2_ASAP7_75t_L g718 ( .A(n_473), .B(n_513), .Y(n_718) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g563 ( .A(n_474), .Y(n_563) );
OAI21x1_ASAP7_75t_SL g474 ( .A1(n_475), .A2(n_477), .B(n_481), .Y(n_474) );
INVx1_ASAP7_75t_L g482 ( .A(n_476), .Y(n_482) );
AND2x2_ASAP7_75t_L g499 ( .A(n_483), .B(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_SL g654 ( .A(n_483), .B(n_562), .Y(n_654) );
AND2x2_ASAP7_75t_L g660 ( .A(n_483), .B(n_501), .Y(n_660) );
AND2x2_ASAP7_75t_L g749 ( .A(n_483), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g731 ( .A(n_489), .Y(n_731) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
BUFx2_ASAP7_75t_L g560 ( .A(n_490), .Y(n_560) );
AND2x2_ASAP7_75t_L g594 ( .A(n_490), .B(n_500), .Y(n_594) );
AND2x2_ASAP7_75t_L g643 ( .A(n_490), .B(n_501), .Y(n_643) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g600 ( .A(n_491), .B(n_501), .Y(n_600) );
INVxp67_ASAP7_75t_L g612 ( .A(n_491), .Y(n_612) );
BUFx3_ASAP7_75t_L g657 ( .A(n_491), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
OAI31xp33_ASAP7_75t_L g553 ( .A1(n_499), .A2(n_554), .A3(n_559), .B(n_564), .Y(n_553) );
AND2x2_ASAP7_75t_L g561 ( .A(n_500), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g580 ( .A(n_501), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_507), .Y(n_502) );
AOI322xp5_ASAP7_75t_L g754 ( .A1(n_509), .A2(n_629), .A3(n_658), .B1(n_663), .B2(n_755), .C1(n_758), .C2(n_759), .Y(n_754) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_510), .B(n_600), .Y(n_605) );
NAND2x1_ASAP7_75t_L g642 ( .A(n_510), .B(n_643), .Y(n_642) );
AND2x4_ASAP7_75t_L g686 ( .A(n_510), .B(n_590), .Y(n_686) );
INVx1_ASAP7_75t_SL g700 ( .A(n_510), .Y(n_700) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g581 ( .A(n_511), .Y(n_581) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_511), .Y(n_724) );
AND2x2_ASAP7_75t_L g653 ( .A(n_512), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_512), .B(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_SL g512 ( .A(n_513), .B(n_514), .Y(n_512) );
BUFx2_ASAP7_75t_L g558 ( .A(n_513), .Y(n_558) );
INVx1_ASAP7_75t_L g750 ( .A(n_513), .Y(n_750) );
OR2x2_ASAP7_75t_L g617 ( .A(n_514), .B(n_562), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_514), .B(n_587), .Y(n_651) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g590 ( .A(n_515), .B(n_562), .Y(n_590) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_536), .Y(n_516) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g646 ( .A(n_518), .Y(n_646) );
OR2x2_ASAP7_75t_L g673 ( .A(n_518), .B(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_529), .Y(n_518) );
NOR2x1_ASAP7_75t_SL g567 ( .A(n_519), .B(n_537), .Y(n_567) );
AND2x2_ASAP7_75t_L g574 ( .A(n_519), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g746 ( .A(n_519), .B(n_608), .Y(n_746) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_527), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_520), .B(n_528), .Y(n_527) );
AO21x2_ASAP7_75t_L g623 ( .A1(n_520), .A2(n_521), .B(n_527), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
OR2x2_ASAP7_75t_L g568 ( .A(n_529), .B(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g577 ( .A(n_529), .Y(n_577) );
INVx2_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
INVx1_ASAP7_75t_L g649 ( .A(n_529), .Y(n_649) );
AND2x2_ASAP7_75t_L g680 ( .A(n_529), .B(n_537), .Y(n_680) );
AND2x2_ASAP7_75t_L g711 ( .A(n_529), .B(n_638), .Y(n_711) );
AND2x2_ASAP7_75t_L g607 ( .A(n_536), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_536), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_SL g710 ( .A(n_536), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g715 ( .A(n_536), .B(n_577), .Y(n_715) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_545), .Y(n_536) );
INVx5_ASAP7_75t_L g575 ( .A(n_537), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_537), .B(n_569), .Y(n_647) );
BUFx2_ASAP7_75t_L g707 ( .A(n_537), .Y(n_707) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx4_ASAP7_75t_L g569 ( .A(n_545), .Y(n_569) );
AND2x2_ASAP7_75t_L g692 ( .A(n_545), .B(n_575), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_555), .A2(n_682), .B1(n_685), .B2(n_687), .C(n_688), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AND2x2_ASAP7_75t_L g703 ( .A(n_556), .B(n_594), .Y(n_703) );
INVx1_ASAP7_75t_SL g729 ( .A(n_556), .Y(n_729) );
AND2x2_ASAP7_75t_L g714 ( .A(n_557), .B(n_686), .Y(n_714) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_558), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g583 ( .A(n_560), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g589 ( .A(n_560), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g613 ( .A(n_561), .Y(n_613) );
AND2x2_ASAP7_75t_L g671 ( .A(n_561), .B(n_599), .Y(n_671) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g596 ( .A(n_563), .Y(n_596) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g592 ( .A(n_568), .Y(n_592) );
OR2x2_ASAP7_75t_L g760 ( .A(n_568), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g576 ( .A(n_569), .Y(n_576) );
AND2x4_ASAP7_75t_L g632 ( .A(n_569), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_569), .B(n_637), .Y(n_636) );
NAND2x1p5_ASAP7_75t_L g674 ( .A(n_569), .B(n_575), .Y(n_674) );
AND2x2_ASAP7_75t_L g734 ( .A(n_569), .B(n_637), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_578), .B1(n_591), .B2(n_593), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_571), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND3x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .C(n_577), .Y(n_573) );
AND2x4_ASAP7_75t_L g591 ( .A(n_574), .B(n_592), .Y(n_591) );
INVx4_ASAP7_75t_L g631 ( .A(n_575), .Y(n_631) );
AND2x2_ASAP7_75t_SL g764 ( .A(n_575), .B(n_632), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_576), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g676 ( .A(n_577), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g741 ( .A1(n_577), .A2(n_706), .A3(n_742), .B1(n_744), .B2(n_747), .C1(n_751), .C2(n_752), .Y(n_741) );
NAND4xp25_ASAP7_75t_SL g578 ( .A(n_579), .B(n_582), .C(n_586), .D(n_588), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_580), .B(n_596), .Y(n_708) );
BUFx2_ASAP7_75t_L g599 ( .A(n_581), .Y(n_599) );
INVx1_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g723 ( .A(n_584), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g737 ( .A(n_585), .B(n_612), .Y(n_737) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g603 ( .A(n_587), .B(n_604), .Y(n_603) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_587), .A2(n_656), .B(n_658), .C(n_661), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_587), .B(n_594), .Y(n_713) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_589), .A2(n_671), .B1(n_672), .B2(n_675), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_590), .A2(n_626), .B1(n_630), .B2(n_634), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_590), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_590), .B(n_727), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_590), .B(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g757 ( .A(n_590), .Y(n_757) );
INVx1_ASAP7_75t_L g696 ( .A(n_591), .Y(n_696) );
OAI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_595), .B(n_597), .Y(n_593) );
INVx1_ASAP7_75t_L g604 ( .A(n_594), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_594), .B(n_599), .Y(n_753) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g689 ( .A(n_596), .B(n_600), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_598), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g756 ( .A(n_599), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g730 ( .A(n_600), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B(n_606), .C(n_609), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI22xp33_ASAP7_75t_SL g716 ( .A1(n_604), .A2(n_635), .B1(n_682), .B2(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_608), .B(n_631), .Y(n_639) );
OR2x2_ASAP7_75t_L g668 ( .A(n_608), .B(n_669), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g609 ( .A1(n_610), .A2(n_614), .B(n_618), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g629 ( .A(n_612), .Y(n_629) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_615), .A2(n_668), .B(n_670), .C(n_678), .Y(n_667) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2xp67_ASAP7_75t_SL g701 ( .A(n_620), .B(n_647), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_620), .Y(n_704) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_622), .B(n_631), .Y(n_761) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g633 ( .A(n_623), .Y(n_633) );
INVx2_ASAP7_75t_L g638 ( .A(n_623), .Y(n_638) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_640), .C(n_652), .D(n_655), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_628), .A2(n_760), .B1(n_762), .B2(n_763), .Y(n_759) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x4_ASAP7_75t_L g727 ( .A(n_631), .B(n_657), .Y(n_727) );
AND2x2_ASAP7_75t_L g648 ( .A(n_632), .B(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g669 ( .A(n_632), .Y(n_669) );
AND2x2_ASAP7_75t_L g679 ( .A(n_632), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_639), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_638), .Y(n_693) );
INVx1_ASAP7_75t_L g683 ( .A(n_639), .Y(n_683) );
AOI32xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .A3(n_647), .B1(n_648), .B2(n_650), .Y(n_640) );
OAI21xp33_ASAP7_75t_L g688 ( .A1(n_641), .A2(n_689), .B(n_690), .Y(n_688) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_644), .A2(n_721), .B1(n_723), .B2(n_725), .C(n_728), .Y(n_720) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g705 ( .A(n_646), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g663 ( .A(n_647), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_648), .A2(n_686), .B1(n_736), .B2(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g662 ( .A(n_649), .Y(n_662) );
AND2x2_ASAP7_75t_L g740 ( .A(n_649), .B(n_693), .Y(n_740) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_656), .B(n_708), .Y(n_743) );
INVx1_ASAP7_75t_L g762 ( .A(n_656), .Y(n_762) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NOR2xp67_ASAP7_75t_L g664 ( .A(n_665), .B(n_719), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_709), .Y(n_665) );
NOR3xp33_ASAP7_75t_SL g666 ( .A(n_667), .B(n_681), .C(n_694), .Y(n_666) );
INVx1_ASAP7_75t_L g684 ( .A(n_669), .Y(n_684) );
INVx1_ASAP7_75t_SL g695 ( .A(n_671), .Y(n_695) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g677 ( .A(n_674), .Y(n_677) );
INVx2_ASAP7_75t_L g687 ( .A(n_675), .Y(n_687) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AND2x4_ASAP7_75t_L g733 ( .A(n_676), .B(n_734), .Y(n_733) );
AND2x4_ASAP7_75t_L g751 ( .A(n_680), .B(n_734), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
AOI32xp33_ASAP7_75t_L g702 ( .A1(n_691), .A2(n_703), .A3(n_704), .B1(n_705), .B2(n_708), .Y(n_702) );
NOR2xp33_ASAP7_75t_SL g721 ( .A(n_691), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_SL g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g722 ( .A(n_693), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_696), .B(n_697), .C(n_702), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g758 ( .A(n_706), .B(n_746), .Y(n_758) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_707), .B(n_746), .Y(n_745) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B1(n_714), .B2(n_715), .C(n_716), .Y(n_709) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
CKINVDCx16_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
NAND4xp25_ASAP7_75t_L g719 ( .A(n_720), .B(n_735), .C(n_741), .D(n_754), .Y(n_719) );
INVxp33_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
O2A1O1Ixp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B(n_731), .C(n_732), .Y(n_728) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx3_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
CKINVDCx5p33_ASAP7_75t_R g768 ( .A(n_769), .Y(n_768) );
INVx3_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_773), .Y(n_780) );
INVx3_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_SL g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_SL g779 ( .A(n_780), .Y(n_779) );
endmodule