module fake_ariane_1550_n_1004 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1004);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1004;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_985;
wire n_245;
wire n_421;
wire n_549;
wire n_760;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_898;
wire n_857;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_758;
wire n_738;
wire n_339;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_721;
wire n_600;
wire n_840;
wire n_398;
wire n_210;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_277;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_644;
wire n_536;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_981;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_34),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_95),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_31),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_40),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_30),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_75),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_201),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_113),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_32),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_8),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_10),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_14),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_20),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_109),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_157),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_72),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_104),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_64),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_15),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_195),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_147),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_69),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_74),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_19),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_165),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_114),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_36),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_129),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

BUFx2_ASAP7_75t_SL g240 ( 
.A(n_152),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_90),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_82),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_163),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_139),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_103),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_146),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_181),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_61),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_48),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_43),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_140),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_98),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_186),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_16),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_117),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_183),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_131),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_51),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_36),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_102),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_71),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_160),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_20),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_87),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_168),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_76),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_53),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_58),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_200),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_107),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_62),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_149),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_46),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_132),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_127),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_77),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_108),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_59),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_27),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_142),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_174),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_17),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_23),
.Y(n_294)
);

CKINVDCx6p67_ASAP7_75t_R g295 ( 
.A(n_222),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_0),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_222),
.B(n_0),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_1),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_2),
.Y(n_300)
);

AND2x4_ASAP7_75t_SL g301 ( 
.A(n_222),
.B(n_3),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_221),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_230),
.B(n_3),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_234),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_242),
.B(n_4),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_243),
.B(n_4),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_215),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_220),
.B(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_245),
.B(n_5),
.Y(n_313)
);

BUFx8_ASAP7_75t_SL g314 ( 
.A(n_206),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_268),
.B(n_214),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_206),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_212),
.B(n_6),
.Y(n_319)
);

AND2x4_ASAP7_75t_L g320 ( 
.A(n_268),
.B(n_6),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_212),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_246),
.B(n_7),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_236),
.B(n_7),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g324 ( 
.A(n_244),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_247),
.B(n_8),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_228),
.Y(n_326)
);

BUFx8_ASAP7_75t_SL g327 ( 
.A(n_207),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_214),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_224),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_249),
.B(n_256),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_260),
.B(n_9),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_267),
.B(n_10),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g333 ( 
.A(n_244),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_224),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_236),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_237),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_255),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_202),
.Y(n_338)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_228),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_228),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_258),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_228),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

BUFx8_ASAP7_75t_L g345 ( 
.A(n_228),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_272),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_283),
.B(n_11),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_L g349 ( 
.A1(n_295),
.A2(n_232),
.B1(n_280),
.B2(n_207),
.Y(n_349)
);

NAND2xp33_ASAP7_75t_SL g350 ( 
.A(n_319),
.B(n_232),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_286),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_296),
.A2(n_330),
.B1(n_306),
.B2(n_297),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_226),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_302),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_319),
.A2(n_280),
.B1(n_229),
.B2(n_290),
.Y(n_355)
);

OA22x2_ASAP7_75t_L g356 ( 
.A1(n_342),
.A2(n_294),
.B1(n_213),
.B2(n_216),
.Y(n_356)
);

AO22x2_ASAP7_75t_L g357 ( 
.A1(n_323),
.A2(n_203),
.B1(n_252),
.B2(n_240),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_312),
.A2(n_204),
.B1(n_211),
.B2(n_217),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_233),
.B1(n_264),
.B2(n_291),
.Y(n_359)
);

AO22x2_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_289),
.B1(n_12),
.B2(n_13),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_301),
.A2(n_288),
.B1(n_287),
.B2(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_295),
.A2(n_284),
.B1(n_281),
.B2(n_279),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g364 ( 
.A(n_301),
.B(n_205),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_321),
.A2(n_277),
.B1(n_275),
.B2(n_274),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_302),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_R g367 ( 
.A1(n_305),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_208),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_338),
.B(n_209),
.Y(n_369)
);

AO22x2_ASAP7_75t_L g370 ( 
.A1(n_312),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_301),
.A2(n_273),
.B1(n_271),
.B2(n_270),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_324),
.A2(n_269),
.B1(n_266),
.B2(n_263),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_302),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_298),
.A2(n_262),
.B1(n_261),
.B2(n_259),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_336),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_304),
.A2(n_238),
.B1(n_254),
.B2(n_253),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_317),
.B(n_210),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_218),
.Y(n_379)
);

AO22x2_ASAP7_75t_L g380 ( 
.A1(n_312),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_309),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_298),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

AO22x2_ASAP7_75t_L g386 ( 
.A1(n_298),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_309),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

AO22x2_ASAP7_75t_L g389 ( 
.A1(n_298),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_389)
);

OR2x6_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_24),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_317),
.B(n_219),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_223),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_300),
.A2(n_257),
.B1(n_251),
.B2(n_250),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_L g397 ( 
.A1(n_324),
.A2(n_248),
.B1(n_241),
.B2(n_239),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_25),
.Y(n_398)
);

AOI22x1_ASAP7_75t_L g399 ( 
.A1(n_320),
.A2(n_235),
.B1(n_227),
.B2(n_225),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_317),
.B(n_26),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_333),
.B(n_342),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_329),
.Y(n_403)
);

OAI22xp33_ASAP7_75t_L g404 ( 
.A1(n_333),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_L g405 ( 
.A1(n_333),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_362),
.A2(n_318),
.B(n_303),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_388),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_354),
.A2(n_313),
.B(n_307),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

NAND2x1p5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_315),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_336),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_310),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_375),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_346),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_355),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_393),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_384),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_379),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_355),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_395),
.B(n_335),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_385),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_376),
.B(n_327),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_392),
.A2(n_331),
.B(n_325),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_391),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_376),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_401),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_377),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_377),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_390),
.B(n_300),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_374),
.B(n_346),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_369),
.B(n_336),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_359),
.B(n_346),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_403),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_359),
.B(n_347),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_400),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_390),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_349),
.B(n_314),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_351),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_349),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_394),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_352),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_361),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_352),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_356),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_356),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_364),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_396),
.B(n_300),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_335),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_360),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_382),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_361),
.B(n_316),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_371),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_386),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_371),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_378),
.A2(n_318),
.B(n_303),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_389),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_363),
.B(n_315),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_372),
.B(n_337),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_358),
.B(n_300),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_363),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_357),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_370),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_365),
.A2(n_318),
.B(n_303),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_412),
.B(n_357),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_412),
.B(n_370),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_372),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_439),
.B(n_380),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_416),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_407),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_438),
.B(n_397),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_413),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_437),
.B(n_397),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_407),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_480),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_438),
.B(n_358),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_449),
.B(n_404),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_415),
.B(n_315),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_461),
.A2(n_380),
.B1(n_367),
.B2(n_405),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_417),
.B(n_320),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_444),
.B(n_347),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_444),
.B(n_347),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_480),
.Y(n_501)
);

AND2x4_ASAP7_75t_SL g502 ( 
.A(n_480),
.B(n_320),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_472),
.A2(n_332),
.B(n_348),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_449),
.B(n_453),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_419),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_409),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_437),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_461),
.B(n_347),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_406),
.A2(n_326),
.B(n_341),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_480),
.B(n_320),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_417),
.B(n_308),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_436),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_462),
.B(n_322),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_404),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_428),
.A2(n_326),
.B(n_343),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_436),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_459),
.B(n_328),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_455),
.B(n_328),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_462),
.B(n_334),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_425),
.B(n_334),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_334),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_426),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_430),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_451),
.B(n_334),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_433),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_410),
.B(n_340),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_440),
.B(n_340),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_477),
.B(n_340),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_435),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_477),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_445),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_460),
.B(n_405),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_477),
.B(n_340),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_441),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_463),
.B(n_340),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_443),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_474),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_421),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_464),
.B(n_340),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_448),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_458),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_452),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_420),
.B(n_335),
.Y(n_552)
);

CKINVDCx16_ASAP7_75t_R g553 ( 
.A(n_478),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_481),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_452),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_408),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_423),
.B(n_335),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_424),
.A2(n_326),
.B(n_343),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_456),
.B(n_335),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_457),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_442),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_465),
.B(n_344),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_R g563 ( 
.A(n_431),
.B(n_345),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_460),
.B(n_335),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_466),
.B(n_344),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_470),
.B(n_344),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_492),
.B(n_499),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_473),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_554),
.B(n_476),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_489),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_492),
.B(n_468),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_560),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_504),
.B(n_479),
.Y(n_573)
);

BUFx12f_ASAP7_75t_L g574 ( 
.A(n_561),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_488),
.B(n_469),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_507),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_501),
.B(n_450),
.Y(n_577)
);

BUFx4f_ASAP7_75t_L g578 ( 
.A(n_561),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_489),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_560),
.Y(n_580)
);

NAND2x1_ASAP7_75t_L g581 ( 
.A(n_520),
.B(n_341),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_539),
.B(n_344),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_491),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_560),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_494),
.B(n_454),
.Y(n_585)
);

OR2x6_ASAP7_75t_L g586 ( 
.A(n_539),
.B(n_467),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_517),
.B(n_446),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_517),
.B(n_446),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_539),
.B(n_344),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_512),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_521),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_512),
.B(n_454),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_512),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_483),
.B(n_431),
.Y(n_595)
);

CKINVDCx10_ASAP7_75t_R g596 ( 
.A(n_553),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_471),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_512),
.B(n_471),
.Y(n_599)
);

NAND2x1_ASAP7_75t_L g600 ( 
.A(n_520),
.B(n_341),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_560),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_483),
.B(n_447),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_508),
.B(n_418),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_539),
.B(n_418),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_561),
.B(n_422),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_521),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_485),
.B(n_482),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_563),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_498),
.B(n_343),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_491),
.B(n_344),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_498),
.B(n_345),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_515),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_500),
.B(n_345),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_502),
.Y(n_616)
);

NOR2x1_ASAP7_75t_L g617 ( 
.A(n_490),
.B(n_427),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_561),
.B(n_422),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_522),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_485),
.B(n_482),
.Y(n_620)
);

BUFx8_ASAP7_75t_L g621 ( 
.A(n_526),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_541),
.B(n_31),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_500),
.B(n_311),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_549),
.B(n_345),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_311),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_516),
.B(n_32),
.Y(n_626)
);

BUFx12f_ASAP7_75t_L g627 ( 
.A(n_522),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_553),
.B(n_311),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_532),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_486),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_546),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_502),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_496),
.B(n_311),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_590),
.Y(n_634)
);

BUFx6f_ASAP7_75t_SL g635 ( 
.A(n_606),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_574),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_585),
.A2(n_496),
.B1(n_484),
.B2(n_547),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_630),
.Y(n_638)
);

OR2x6_ASAP7_75t_SL g639 ( 
.A(n_610),
.B(n_495),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_594),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_616),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_575),
.B(n_549),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_578),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_570),
.Y(n_644)
);

CKINVDCx6p67_ASAP7_75t_R g645 ( 
.A(n_596),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_590),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_621),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_568),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_587),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_616),
.B(n_502),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_572),
.B(n_565),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_629),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_571),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_632),
.Y(n_654)
);

BUFx4f_ASAP7_75t_SL g655 ( 
.A(n_621),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_632),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_579),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_575),
.B(n_535),
.Y(n_658)
);

INVx1_ASAP7_75t_SL g659 ( 
.A(n_607),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_607),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_614),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_585),
.B(n_535),
.Y(n_662)
);

BUFx12f_ASAP7_75t_L g663 ( 
.A(n_586),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_614),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_568),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_569),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_578),
.Y(n_667)
);

BUFx4f_ASAP7_75t_L g668 ( 
.A(n_619),
.Y(n_668)
);

BUFx2_ASAP7_75t_SL g669 ( 
.A(n_594),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_588),
.Y(n_670)
);

BUFx2_ASAP7_75t_SL g671 ( 
.A(n_601),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_586),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_569),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_567),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_586),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_614),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_601),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_598),
.B(n_526),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_593),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_627),
.Y(n_682)
);

CKINVDCx8_ASAP7_75t_R g683 ( 
.A(n_606),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_591),
.Y(n_684)
);

INVx6_ASAP7_75t_L g685 ( 
.A(n_597),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_598),
.A2(n_550),
.B1(n_565),
.B2(n_544),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_609),
.B(n_537),
.Y(n_687)
);

INVx6_ASAP7_75t_SL g688 ( 
.A(n_618),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_597),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_628),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_567),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_637),
.A2(n_622),
.B1(n_626),
.B2(n_617),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_642),
.A2(n_622),
.B1(n_633),
.B2(n_604),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_638),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_644),
.Y(n_695)
);

BUFx4f_ASAP7_75t_SL g696 ( 
.A(n_645),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_662),
.A2(n_626),
.B1(n_605),
.B2(n_599),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_643),
.Y(n_698)
);

INVx6_ASAP7_75t_L g699 ( 
.A(n_643),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_679),
.A2(n_605),
.B1(n_592),
.B2(n_599),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_644),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_681),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_691),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_657),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_649),
.A2(n_514),
.B1(n_503),
.B2(n_540),
.Y(n_705)
);

CKINVDCx6p67_ASAP7_75t_R g706 ( 
.A(n_645),
.Y(n_706)
);

INVx6_ASAP7_75t_L g707 ( 
.A(n_654),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_681),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_657),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_L g710 ( 
.A1(n_658),
.A2(n_540),
.B1(n_486),
.B2(n_505),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_670),
.A2(n_595),
.B1(n_592),
.B2(n_603),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_635),
.A2(n_573),
.B1(n_618),
.B2(n_620),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_684),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_684),
.Y(n_714)
);

BUFx2_ASAP7_75t_L g715 ( 
.A(n_691),
.Y(n_715)
);

CKINVDCx6p67_ASAP7_75t_R g716 ( 
.A(n_682),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_648),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_647),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_665),
.Y(n_719)
);

INVx6_ASAP7_75t_L g720 ( 
.A(n_654),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_635),
.A2(n_573),
.B1(n_577),
.B2(n_506),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_683),
.A2(n_618),
.B1(n_505),
.B2(n_550),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_666),
.B(n_577),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_SL g724 ( 
.A1(n_635),
.A2(n_550),
.B1(n_615),
.B2(n_613),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_668),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_686),
.A2(n_602),
.B1(n_584),
.B2(n_580),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_652),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_659),
.A2(n_510),
.B1(n_506),
.B2(n_537),
.Y(n_728)
);

BUFx8_ASAP7_75t_L g729 ( 
.A(n_636),
.Y(n_729)
);

INVx5_ASAP7_75t_L g730 ( 
.A(n_651),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_655),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_653),
.B(n_576),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_634),
.A2(n_497),
.B1(n_487),
.B2(n_583),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_673),
.Y(n_734)
);

BUFx10_ASAP7_75t_L g735 ( 
.A(n_647),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_678),
.Y(n_736)
);

BUFx8_ASAP7_75t_L g737 ( 
.A(n_636),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_675),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_660),
.A2(n_510),
.B1(n_542),
.B2(n_523),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_674),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_682),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_SL g742 ( 
.A1(n_675),
.A2(n_613),
.B1(n_615),
.B2(n_542),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_651),
.A2(n_571),
.B1(n_565),
.B2(n_544),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_641),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_687),
.A2(n_523),
.B1(n_529),
.B2(n_528),
.Y(n_745)
);

INVx1_ASAP7_75t_SL g746 ( 
.A(n_727),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_696),
.Y(n_747)
);

INVx5_ASAP7_75t_SL g748 ( 
.A(n_706),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_692),
.A2(n_639),
.B1(n_683),
.B2(n_674),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_694),
.Y(n_750)
);

OAI21xp33_ASAP7_75t_L g751 ( 
.A1(n_692),
.A2(n_556),
.B(n_530),
.Y(n_751)
);

OAI21xp5_ASAP7_75t_L g752 ( 
.A1(n_705),
.A2(n_624),
.B(n_611),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_697),
.A2(n_639),
.B1(n_646),
.B2(n_668),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_736),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_695),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_693),
.A2(n_687),
.B1(n_663),
.B2(n_688),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_693),
.A2(n_663),
.B1(n_688),
.B2(n_531),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_740),
.B(n_672),
.Y(n_758)
);

BUFx3_ASAP7_75t_L g759 ( 
.A(n_729),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_SL g760 ( 
.A1(n_730),
.A2(n_672),
.B1(n_668),
.B2(n_690),
.Y(n_760)
);

OAI22xp33_ASAP7_75t_L g761 ( 
.A1(n_743),
.A2(n_688),
.B1(n_677),
.B2(n_667),
.Y(n_761)
);

NAND2x1p5_ASAP7_75t_L g762 ( 
.A(n_730),
.B(n_654),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_717),
.Y(n_763)
);

NAND2x1p5_ASAP7_75t_L g764 ( 
.A(n_730),
.B(n_654),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_730),
.A2(n_525),
.B1(n_651),
.B2(n_671),
.Y(n_765)
);

OAI21xp33_ASAP7_75t_L g766 ( 
.A1(n_697),
.A2(n_556),
.B(n_527),
.Y(n_766)
);

AO22x1_ASAP7_75t_L g767 ( 
.A1(n_729),
.A2(n_680),
.B1(n_667),
.B2(n_677),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_700),
.A2(n_531),
.B1(n_528),
.B2(n_529),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_732),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_700),
.A2(n_624),
.B1(n_651),
.B2(n_608),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_711),
.B(n_680),
.Y(n_771)
);

BUFx12f_ASAP7_75t_L g772 ( 
.A(n_718),
.Y(n_772)
);

INVx1_ASAP7_75t_SL g773 ( 
.A(n_738),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_710),
.A2(n_611),
.B(n_518),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_742),
.A2(n_651),
.B1(n_623),
.B2(n_544),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_742),
.A2(n_651),
.B1(n_544),
.B2(n_522),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_703),
.B(n_548),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_745),
.A2(n_589),
.B1(n_582),
.B2(n_671),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_SL g779 ( 
.A1(n_722),
.A2(n_656),
.B(n_589),
.Y(n_779)
);

INVx1_ASAP7_75t_SL g780 ( 
.A(n_741),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_745),
.A2(n_582),
.B1(n_641),
.B2(n_656),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_723),
.A2(n_545),
.B(n_543),
.Y(n_782)
);

AOI22xp33_ASAP7_75t_L g783 ( 
.A1(n_739),
.A2(n_534),
.B1(n_562),
.B2(n_566),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_721),
.A2(n_534),
.B1(n_562),
.B2(n_566),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_721),
.A2(n_548),
.B1(n_551),
.B2(n_545),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_722),
.A2(n_551),
.B1(n_543),
.B2(n_538),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_712),
.A2(n_538),
.B1(n_536),
.B2(n_533),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_719),
.Y(n_788)
);

INVxp33_ASAP7_75t_L g789 ( 
.A(n_698),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_734),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_712),
.A2(n_551),
.B1(n_536),
.B2(n_533),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_728),
.A2(n_551),
.B1(n_524),
.B2(n_519),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_715),
.B(n_689),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_724),
.A2(n_551),
.B1(n_524),
.B2(n_519),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_701),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_725),
.A2(n_641),
.B1(n_656),
.B2(n_487),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_737),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_704),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_698),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_713),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_724),
.A2(n_513),
.B1(n_511),
.B2(n_669),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_SL g802 ( 
.A1(n_744),
.A2(n_650),
.B(n_640),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_726),
.A2(n_487),
.B1(n_583),
.B2(n_669),
.Y(n_803)
);

INVx4_ASAP7_75t_L g804 ( 
.A(n_716),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_757),
.A2(n_709),
.B1(n_714),
.B2(n_511),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_756),
.A2(n_744),
.B1(n_699),
.B2(n_702),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_757),
.A2(n_513),
.B1(n_625),
.B2(n_555),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_771),
.A2(n_625),
.B1(n_555),
.B2(n_640),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_750),
.B(n_33),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_756),
.A2(n_699),
.B1(n_733),
.B2(n_708),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_769),
.B(n_698),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_SL g812 ( 
.A1(n_749),
.A2(n_720),
.B1(n_707),
.B2(n_699),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_754),
.B(n_33),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_746),
.B(n_698),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_758),
.B(n_689),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_770),
.A2(n_625),
.B1(n_555),
.B2(n_640),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_763),
.B(n_737),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_795),
.B(n_34),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_799),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_SL g820 ( 
.A1(n_753),
.A2(n_720),
.B1(n_707),
.B2(n_640),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_SL g821 ( 
.A1(n_803),
.A2(n_720),
.B1(n_707),
.B2(n_640),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_798),
.Y(n_822)
);

BUFx4f_ASAP7_75t_SL g823 ( 
.A(n_747),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_802),
.B(n_664),
.C(n_661),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_SL g825 ( 
.A1(n_782),
.A2(n_764),
.B(n_762),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_786),
.A2(n_696),
.B1(n_731),
.B2(n_654),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_779),
.A2(n_597),
.B1(n_685),
.B2(n_676),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_770),
.A2(n_625),
.B1(n_555),
.B2(n_311),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_788),
.B(n_661),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_776),
.A2(n_311),
.B1(n_329),
.B2(n_552),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_SL g831 ( 
.A1(n_778),
.A2(n_685),
.B1(n_329),
.B2(n_676),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_776),
.A2(n_329),
.B1(n_557),
.B2(n_685),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_786),
.A2(n_661),
.B1(n_664),
.B2(n_676),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_790),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_766),
.A2(n_329),
.B1(n_685),
.B2(n_515),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_787),
.A2(n_515),
.B1(n_564),
.B2(n_520),
.Y(n_836)
);

OAI21xp33_ASAP7_75t_L g837 ( 
.A1(n_752),
.A2(n_299),
.B(n_664),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_SL g838 ( 
.A1(n_781),
.A2(n_735),
.B1(n_612),
.B2(n_515),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_775),
.A2(n_515),
.B1(n_520),
.B2(n_487),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_775),
.A2(n_559),
.B1(n_299),
.B2(n_612),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_SL g841 ( 
.A1(n_777),
.A2(n_735),
.B1(n_339),
.B2(n_509),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_791),
.A2(n_558),
.B1(n_581),
.B2(n_600),
.Y(n_842)
);

OAI222xp33_ASAP7_75t_L g843 ( 
.A1(n_760),
.A2(n_339),
.B1(n_37),
.B2(n_38),
.C1(n_39),
.C2(n_35),
.Y(n_843)
);

OAI222xp33_ASAP7_75t_L g844 ( 
.A1(n_801),
.A2(n_339),
.B1(n_37),
.B2(n_38),
.C1(n_39),
.C2(n_35),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_791),
.A2(n_768),
.B1(n_751),
.B2(n_785),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_768),
.A2(n_785),
.B1(n_801),
.B2(n_792),
.Y(n_846)
);

AOI221xp5_ASAP7_75t_L g847 ( 
.A1(n_773),
.A2(n_339),
.B1(n_42),
.B2(n_44),
.C(n_45),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_774),
.A2(n_339),
.B1(n_509),
.B2(n_50),
.Y(n_848)
);

NAND3xp33_ASAP7_75t_L g849 ( 
.A(n_794),
.B(n_339),
.C(n_47),
.Y(n_849)
);

NOR3xp33_ASAP7_75t_L g850 ( 
.A(n_843),
.B(n_844),
.C(n_810),
.Y(n_850)
);

NAND3xp33_ASAP7_75t_L g851 ( 
.A(n_849),
.B(n_767),
.C(n_794),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_811),
.B(n_793),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_822),
.B(n_793),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_822),
.B(n_789),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_834),
.A2(n_800),
.B(n_755),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_845),
.A2(n_792),
.B1(n_784),
.B2(n_783),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_827),
.B(n_761),
.Y(n_857)
);

NAND3xp33_ASAP7_75t_L g858 ( 
.A(n_849),
.B(n_804),
.C(n_796),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_819),
.B(n_780),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_809),
.B(n_804),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_SL g861 ( 
.A(n_809),
.B(n_765),
.C(n_783),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_813),
.B(n_759),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_813),
.B(n_818),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_818),
.B(n_748),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_834),
.B(n_797),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_846),
.A2(n_826),
.B1(n_812),
.B2(n_837),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_815),
.B(n_748),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_814),
.B(n_748),
.Y(n_868)
);

OAI221xp5_ASAP7_75t_L g869 ( 
.A1(n_817),
.A2(n_784),
.B1(n_764),
.B2(n_762),
.C(n_772),
.Y(n_869)
);

OAI221xp5_ASAP7_75t_SL g870 ( 
.A1(n_837),
.A2(n_41),
.B1(n_52),
.B2(n_54),
.C(n_55),
.Y(n_870)
);

NAND3xp33_ASAP7_75t_L g871 ( 
.A(n_847),
.B(n_56),
.C(n_57),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_829),
.B(n_60),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_824),
.B(n_63),
.Y(n_873)
);

OAI221xp5_ASAP7_75t_SL g874 ( 
.A1(n_820),
.A2(n_816),
.B1(n_838),
.B2(n_831),
.C(n_828),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_833),
.B(n_821),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_65),
.Y(n_876)
);

AOI221xp5_ASAP7_75t_L g877 ( 
.A1(n_806),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.C(n_73),
.Y(n_877)
);

OAI221xp5_ASAP7_75t_SL g878 ( 
.A1(n_805),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_833),
.Y(n_879)
);

AOI221xp5_ASAP7_75t_L g880 ( 
.A1(n_850),
.A2(n_832),
.B1(n_835),
.B2(n_830),
.C(n_848),
.Y(n_880)
);

OAI211xp5_ASAP7_75t_SL g881 ( 
.A1(n_860),
.A2(n_841),
.B(n_808),
.C(n_825),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_851),
.B(n_839),
.C(n_807),
.Y(n_882)
);

OR2x2_ASAP7_75t_L g883 ( 
.A(n_863),
.B(n_853),
.Y(n_883)
);

NAND4xp75_ASAP7_75t_L g884 ( 
.A(n_875),
.B(n_825),
.C(n_836),
.D(n_840),
.Y(n_884)
);

NOR2x1_ASAP7_75t_L g885 ( 
.A(n_867),
.B(n_842),
.Y(n_885)
);

OA211x2_ASAP7_75t_L g886 ( 
.A1(n_858),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_859),
.B(n_86),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_852),
.B(n_88),
.Y(n_888)
);

AO21x2_ASAP7_75t_L g889 ( 
.A1(n_851),
.A2(n_89),
.B(n_91),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_859),
.B(n_92),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_879),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_891)
);

NAND4xp25_ASAP7_75t_L g892 ( 
.A(n_858),
.B(n_97),
.C(n_99),
.D(n_100),
.Y(n_892)
);

OAI211xp5_ASAP7_75t_SL g893 ( 
.A1(n_867),
.A2(n_864),
.B(n_868),
.C(n_876),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_854),
.B(n_101),
.Y(n_894)
);

OR2x2_ASAP7_75t_SL g895 ( 
.A(n_861),
.B(n_105),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_855),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_866),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_862),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_871),
.B(n_870),
.C(n_878),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_854),
.B(n_112),
.Y(n_900)
);

BUFx2_ASAP7_75t_L g901 ( 
.A(n_898),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_883),
.Y(n_902)
);

AO22x2_ASAP7_75t_L g903 ( 
.A1(n_896),
.A2(n_865),
.B1(n_879),
.B2(n_862),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_885),
.B(n_865),
.Y(n_904)
);

XNOR2xp5_ASAP7_75t_L g905 ( 
.A(n_887),
.B(n_869),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_890),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_894),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_900),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_893),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_899),
.A2(n_857),
.B1(n_871),
.B2(n_856),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_889),
.B(n_855),
.Y(n_911)
);

NAND4xp75_ASAP7_75t_L g912 ( 
.A(n_886),
.B(n_877),
.C(n_873),
.D(n_872),
.Y(n_912)
);

NOR2x1_ASAP7_75t_L g913 ( 
.A(n_892),
.B(n_872),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_909),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_903),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_902),
.B(n_889),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_902),
.Y(n_917)
);

CKINVDCx16_ASAP7_75t_R g918 ( 
.A(n_904),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_913),
.A2(n_892),
.B1(n_882),
.B2(n_897),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_908),
.Y(n_920)
);

XOR2x2_ASAP7_75t_L g921 ( 
.A(n_905),
.B(n_884),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_914),
.A2(n_911),
.B1(n_907),
.B2(n_904),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_917),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_915),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_918),
.Y(n_925)
);

AOI22x1_ASAP7_75t_L g926 ( 
.A1(n_920),
.A2(n_903),
.B1(n_906),
.B2(n_901),
.Y(n_926)
);

INVx2_ASAP7_75t_SL g927 ( 
.A(n_920),
.Y(n_927)
);

OA22x2_ASAP7_75t_L g928 ( 
.A1(n_915),
.A2(n_910),
.B1(n_906),
.B2(n_911),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_916),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_919),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_923),
.Y(n_931)
);

INVxp33_ASAP7_75t_L g932 ( 
.A(n_925),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_927),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_927),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_924),
.Y(n_935)
);

NAND4xp25_ASAP7_75t_SL g936 ( 
.A(n_933),
.B(n_930),
.C(n_928),
.D(n_922),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_931),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_932),
.A2(n_926),
.B1(n_922),
.B2(n_928),
.Y(n_938)
);

NOR4xp25_ASAP7_75t_L g939 ( 
.A(n_936),
.B(n_934),
.C(n_935),
.D(n_924),
.Y(n_939)
);

HB1xp67_ASAP7_75t_L g940 ( 
.A(n_937),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_938),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_937),
.Y(n_942)
);

AO22x1_ASAP7_75t_L g943 ( 
.A1(n_941),
.A2(n_932),
.B1(n_929),
.B2(n_921),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_939),
.A2(n_922),
.B1(n_942),
.B2(n_940),
.Y(n_944)
);

OAI22xp33_ASAP7_75t_SL g945 ( 
.A1(n_942),
.A2(n_874),
.B1(n_895),
.B2(n_888),
.Y(n_945)
);

OA22x2_ASAP7_75t_L g946 ( 
.A1(n_942),
.A2(n_903),
.B1(n_912),
.B2(n_881),
.Y(n_946)
);

NOR2x1_ASAP7_75t_L g947 ( 
.A(n_942),
.B(n_882),
.Y(n_947)
);

OA22x2_ASAP7_75t_L g948 ( 
.A1(n_941),
.A2(n_880),
.B1(n_891),
.B2(n_855),
.Y(n_948)
);

INVxp67_ASAP7_75t_SL g949 ( 
.A(n_942),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_944),
.B(n_115),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_949),
.B(n_118),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_947),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_943),
.B(n_120),
.Y(n_953)
);

NOR2x1_ASAP7_75t_L g954 ( 
.A(n_946),
.B(n_945),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_948),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_949),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_956),
.Y(n_957)
);

NAND5xp2_ASAP7_75t_L g958 ( 
.A(n_952),
.B(n_121),
.C(n_123),
.D(n_124),
.E(n_125),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_955),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_950),
.A2(n_855),
.B1(n_128),
.B2(n_130),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_951),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_954),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_953),
.A2(n_126),
.B1(n_134),
.B2(n_136),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_957),
.Y(n_964)
);

INVxp67_ASAP7_75t_SL g965 ( 
.A(n_962),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_961),
.B(n_137),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_959),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_958),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_963),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_960),
.Y(n_970)
);

AOI22x1_ASAP7_75t_L g971 ( 
.A1(n_957),
.A2(n_138),
.B1(n_141),
.B2(n_143),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_957),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_957),
.B(n_144),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_965),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_SL g975 ( 
.A1(n_964),
.A2(n_145),
.B1(n_148),
.B2(n_151),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_973),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_972),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_967),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_968),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_966),
.Y(n_980)
);

OAI22x1_ASAP7_75t_L g981 ( 
.A1(n_969),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_970),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_969),
.A2(n_161),
.B1(n_166),
.B2(n_167),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_SL g984 ( 
.A1(n_971),
.A2(n_169),
.B1(n_170),
.B2(n_171),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_974),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_976),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_977),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_981),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_978),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_980),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_979),
.Y(n_991)
);

AO22x2_ASAP7_75t_L g992 ( 
.A1(n_986),
.A2(n_975),
.B1(n_984),
.B2(n_983),
.Y(n_992)
);

AOI221xp5_ASAP7_75t_L g993 ( 
.A1(n_991),
.A2(n_982),
.B1(n_173),
.B2(n_175),
.C(n_176),
.Y(n_993)
);

AO22x2_ASAP7_75t_L g994 ( 
.A1(n_987),
.A2(n_172),
.B1(n_177),
.B2(n_178),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_992),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_994),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_996),
.A2(n_985),
.B1(n_988),
.B2(n_989),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_995),
.A2(n_990),
.B1(n_993),
.B2(n_182),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_995),
.A2(n_179),
.B1(n_180),
.B2(n_185),
.Y(n_999)
);

INVxp67_ASAP7_75t_SL g1000 ( 
.A(n_997),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_998),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_999),
.Y(n_1002)
);

OAI221xp5_ASAP7_75t_L g1003 ( 
.A1(n_1000),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.C(n_192),
.Y(n_1003)
);

AOI211xp5_ASAP7_75t_L g1004 ( 
.A1(n_1003),
.A2(n_1001),
.B(n_1002),
.C(n_193),
.Y(n_1004)
);


endmodule