module fake_jpeg_30776_n_541 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_541);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_541;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g140 ( 
.A(n_55),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_89),
.Y(n_106)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_59),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_32),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_0),
.B(n_2),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_47),
.C(n_45),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_83),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_0),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_93),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_2),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_2),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_103),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_100),
.Y(n_148)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_101),
.Y(n_133)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_24),
.B(n_35),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_118),
.B(n_48),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_86),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_122),
.B(n_137),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_57),
.B(n_45),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_34),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_81),
.A2(n_41),
.B1(n_44),
.B2(n_48),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_126),
.A2(n_158),
.B1(n_36),
.B2(n_23),
.Y(n_178)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_55),
.B(n_51),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_55),
.B(n_37),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_138),
.B(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_53),
.A2(n_21),
.B1(n_51),
.B2(n_35),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_150),
.B1(n_26),
.B2(n_30),
.Y(n_189)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_63),
.A2(n_37),
.B1(n_47),
.B2(n_49),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_59),
.Y(n_157)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_71),
.A2(n_50),
.B1(n_34),
.B2(n_39),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_162),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_93),
.B(n_50),
.Y(n_164)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_169),
.B(n_170),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_39),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_171),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_117),
.B(n_87),
.C(n_69),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_172),
.B(n_212),
.Y(n_258)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_115),
.A2(n_36),
.B1(n_76),
.B2(n_30),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_173),
.B(n_194),
.Y(n_255)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_178),
.A2(n_218),
.B1(n_166),
.B2(n_132),
.Y(n_251)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_179),
.Y(n_249)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_100),
.B1(n_98),
.B2(n_97),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_183),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_244)
);

INVx3_ASAP7_75t_SL g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_184),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_192),
.Y(n_235)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_104),
.Y(n_188)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_131),
.A2(n_96),
.B1(n_95),
.B2(n_88),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_77),
.B1(n_78),
.B2(n_84),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_139),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_105),
.A2(n_30),
.B(n_26),
.Y(n_193)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_129),
.B(n_143),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_116),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_139),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_198),
.B(n_221),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_109),
.Y(n_199)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_199),
.Y(n_278)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_200),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_131),
.A2(n_80),
.B1(n_145),
.B2(n_148),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_201),
.A2(n_216),
.B1(n_166),
.B2(n_143),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_204),
.Y(n_261)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_136),
.Y(n_205)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_206),
.Y(n_276)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_154),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

NAND3xp33_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_26),
.C(n_23),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_108),
.B(n_23),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_210),
.B(n_209),
.Y(n_254)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_112),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_105),
.B(n_48),
.C(n_44),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_126),
.A2(n_36),
.B1(n_76),
.B2(n_93),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_213),
.B(n_214),
.Y(n_266)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_110),
.Y(n_215)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_215),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_108),
.A2(n_48),
.B1(n_44),
.B2(n_41),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_127),
.A2(n_44),
.B1(n_41),
.B2(n_22),
.Y(n_218)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_222),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_134),
.Y(n_223)
);

BUFx4f_ASAP7_75t_SL g241 ( 
.A(n_223),
.Y(n_241)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_119),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_225),
.Y(n_253)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_111),
.B(n_22),
.C(n_4),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_226),
.A2(n_22),
.B(n_4),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g227 ( 
.A(n_114),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_132),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_228),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_229),
.Y(n_272)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_193),
.A2(n_160),
.B(n_135),
.C(n_163),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_230),
.B(n_231),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_165),
.B1(n_152),
.B2(n_167),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_234),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_310)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_22),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_243),
.B(n_254),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_245),
.A2(n_262),
.B1(n_263),
.B2(n_270),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_223),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_173),
.B(n_149),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_257),
.B(n_227),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g313 ( 
.A(n_259),
.B(n_16),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_196),
.B(n_3),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_268),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_173),
.A2(n_149),
.B1(n_134),
.B2(n_22),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_183),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_195),
.B(n_6),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_213),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_213),
.A2(n_16),
.B1(n_9),
.B2(n_10),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_275),
.A2(n_218),
.B1(n_184),
.B2(n_180),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_174),
.B(n_8),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_8),
.Y(n_306)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_298),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_181),
.C(n_175),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_283),
.B(n_320),
.Y(n_342)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_280),
.Y(n_284)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_285),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_286),
.B(n_291),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_185),
.B1(n_168),
.B2(n_176),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_287),
.A2(n_272),
.B1(n_271),
.B2(n_232),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_295),
.Y(n_329)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_266),
.A2(n_182),
.B(n_186),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_290),
.A2(n_292),
.B(n_278),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_266),
.A2(n_171),
.B(n_215),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_293),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_203),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_248),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_258),
.B(n_197),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_299),
.B(n_308),
.Y(n_353)
);

AO22x1_ASAP7_75t_SL g300 ( 
.A1(n_257),
.A2(n_208),
.B1(n_201),
.B2(n_190),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_309),
.Y(n_339)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_250),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_224),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

AOI32xp33_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_229),
.A3(n_199),
.B1(n_188),
.B2(n_219),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_SL g346 ( 
.A(n_305),
.B(n_313),
.C(n_241),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_317),
.Y(n_341)
);

BUFx24_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_307),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_240),
.B(n_222),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_179),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_239),
.B1(n_267),
.B2(n_272),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_230),
.B(n_11),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_311),
.B(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_254),
.B(n_277),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_243),
.B(n_12),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_315),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_12),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_253),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_247),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_318),
.B(n_319),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_12),
.C(n_13),
.Y(n_320)
);

OAI32xp33_ASAP7_75t_L g321 ( 
.A1(n_251),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_323),
.Y(n_359)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_322),
.Y(n_366)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_325),
.Y(n_365)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_261),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_237),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_239),
.B1(n_237),
.B2(n_249),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_328),
.A2(n_349),
.B1(n_364),
.B2(n_295),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_291),
.A2(n_303),
.B1(n_317),
.B2(n_282),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_333),
.A2(n_360),
.B1(n_335),
.B2(n_337),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_294),
.A2(n_265),
.B1(n_232),
.B2(n_256),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_335),
.A2(n_337),
.B1(n_344),
.B2(n_354),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_294),
.A2(n_265),
.B1(n_256),
.B2(n_271),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_288),
.A2(n_252),
.B1(n_276),
.B2(n_269),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_346),
.A2(n_351),
.B(n_357),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_291),
.A2(n_276),
.B1(n_252),
.B2(n_242),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_297),
.A2(n_242),
.B(n_260),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_307),
.B(n_330),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_303),
.A2(n_321),
.B1(n_297),
.B2(n_286),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_311),
.A2(n_249),
.B1(n_274),
.B2(n_233),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_299),
.B(n_238),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_283),
.C(n_314),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_324),
.A2(n_274),
.B1(n_233),
.B2(n_264),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_308),
.B(n_264),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_285),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_300),
.A2(n_241),
.B1(n_13),
.B2(n_15),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_397),
.Y(n_427)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_368),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_380),
.B1(n_387),
.B2(n_391),
.Y(n_412)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_332),
.B(n_296),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_372),
.B(n_375),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_353),
.B(n_356),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_341),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_343),
.B(n_312),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_351),
.A2(n_309),
.B(n_292),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_376),
.A2(n_382),
.B(n_398),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_361),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_396),
.Y(n_411)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_343),
.B(n_315),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_395),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_339),
.A2(n_304),
.B1(n_300),
.B2(n_290),
.Y(n_380)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_361),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_389),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_346),
.A2(n_313),
.B(n_320),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_313),
.C(n_319),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_384),
.B(n_394),
.C(n_347),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_385),
.Y(n_425)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_386),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_339),
.A2(n_310),
.B1(n_302),
.B2(n_301),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_360),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_344),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_352),
.A2(n_322),
.B1(n_325),
.B2(n_316),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_359),
.A2(n_241),
.B1(n_307),
.B2(n_364),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_392),
.A2(n_336),
.B1(n_365),
.B2(n_358),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_393),
.A2(n_401),
.B(n_388),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_363),
.C(n_342),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_332),
.Y(n_395)
);

NAND2x1p5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_329),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_329),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_360),
.A2(n_359),
.B(n_350),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_399),
.A2(n_349),
.B1(n_328),
.B2(n_348),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_347),
.A2(n_348),
.B(n_341),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_403),
.A2(n_412),
.B1(n_428),
.B2(n_419),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_404),
.B(n_405),
.Y(n_458)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_406),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_345),
.Y(n_408)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_345),
.Y(n_409)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_340),
.Y(n_410)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_410),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_377),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_432),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_401),
.B(n_334),
.Y(n_415)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_415),
.Y(n_452)
);

AOI22x1_ASAP7_75t_L g419 ( 
.A1(n_396),
.A2(n_366),
.B1(n_333),
.B2(n_358),
.Y(n_419)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_419),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_340),
.C(n_334),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_423),
.C(n_424),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_421),
.A2(n_383),
.B1(n_370),
.B2(n_386),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_383),
.A2(n_336),
.B1(n_365),
.B2(n_362),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_422),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_397),
.B(n_374),
.C(n_384),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_367),
.B(n_362),
.C(n_388),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_429),
.B(n_382),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_393),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_378),
.C(n_368),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_373),
.A2(n_389),
.B(n_400),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_385),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_387),
.Y(n_435)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_435),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_417),
.A2(n_400),
.B(n_376),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_436),
.A2(n_438),
.B(n_446),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_399),
.Y(n_438)
);

OAI22x1_ASAP7_75t_L g442 ( 
.A1(n_411),
.A2(n_369),
.B1(n_373),
.B2(n_396),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_442),
.A2(n_402),
.B(n_429),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_411),
.B(n_392),
.Y(n_443)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_444),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_417),
.A2(n_369),
.B(n_391),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_445),
.A2(n_431),
.B(n_430),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_371),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_450),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_448),
.B(n_457),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_409),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_437),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_453),
.A2(n_412),
.B1(n_421),
.B2(n_406),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_427),
.B(n_420),
.C(n_405),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_427),
.C(n_424),
.Y(n_469)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_425),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_425),
.Y(n_479)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_452),
.B(n_410),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_460),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_461),
.A2(n_456),
.B1(n_434),
.B2(n_449),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_435),
.B(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_462),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_457),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_464),
.B(n_469),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_440),
.A2(n_419),
.B1(n_402),
.B2(n_426),
.Y(n_466)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_466),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_407),
.Y(n_467)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_467),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_471),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_449),
.B(n_416),
.Y(n_470)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_470),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_423),
.C(n_404),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_480),
.C(n_451),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_430),
.Y(n_473)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_431),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_478),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_479),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_437),
.B(n_413),
.C(n_458),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_466),
.A2(n_442),
.B1(n_440),
.B2(n_438),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_492),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_483),
.B(n_493),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_475),
.A2(n_456),
.B1(n_453),
.B2(n_443),
.Y(n_486)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_461),
.A2(n_438),
.B1(n_448),
.B2(n_445),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_460),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_494),
.A2(n_463),
.B1(n_474),
.B2(n_439),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_446),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_467),
.C(n_470),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_489),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_505),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_471),
.C(n_480),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_501),
.C(n_502),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_495),
.A2(n_476),
.B(n_468),
.Y(n_500)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_500),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_469),
.C(n_472),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_485),
.B(n_478),
.C(n_475),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_488),
.A2(n_476),
.B(n_479),
.Y(n_504)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_504),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_497),
.B(n_436),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_481),
.A2(n_474),
.B1(n_441),
.B2(n_459),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_481),
.A2(n_462),
.B1(n_465),
.B2(n_463),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_487),
.B1(n_490),
.B2(n_441),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_511),
.A2(n_484),
.B1(n_487),
.B2(n_502),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_503),
.A2(n_491),
.B1(n_482),
.B2(n_496),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_517),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_508),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_518),
.B(n_519),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_465),
.Y(n_520)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_509),
.C(n_506),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_499),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_522),
.B(n_526),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_515),
.A2(n_507),
.B1(n_494),
.B2(n_511),
.Y(n_525)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_525),
.Y(n_531)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_516),
.A2(n_473),
.B(n_464),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_527),
.A2(n_517),
.B1(n_518),
.B2(n_512),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_528),
.A2(n_530),
.B(n_512),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_514),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_529),
.B(n_524),
.C(n_521),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_532),
.A2(n_533),
.B(n_455),
.Y(n_535)
);

AOI21xp33_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_531),
.B(n_524),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_535),
.B(n_528),
.Y(n_536)
);

NAND3xp33_ASAP7_75t_L g537 ( 
.A(n_536),
.B(n_413),
.C(n_509),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_519),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_459),
.C(n_434),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_488),
.Y(n_541)
);


endmodule