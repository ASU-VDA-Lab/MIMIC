module fake_jpeg_2107_n_382 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_8),
.B(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_45),
.Y(n_113)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_56),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_79),
.B(n_80),
.Y(n_90)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_18),
.B(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_29),
.B(n_12),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_60),
.B(n_65),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_19),
.B(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_70),
.Y(n_105)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_67),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_68),
.Y(n_124)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_73),
.Y(n_87)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_78),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_19),
.B(n_9),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_82),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_84),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_37),
.B1(n_42),
.B2(n_35),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_95),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_38),
.B1(n_36),
.B2(n_39),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_38),
.B1(n_36),
.B2(n_39),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_22),
.B1(n_40),
.B2(n_34),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_92),
.A2(n_110),
.B1(n_127),
.B2(n_129),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_51),
.B1(n_22),
.B2(n_34),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_51),
.A2(n_32),
.B1(n_40),
.B2(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_97),
.A2(n_114),
.B1(n_121),
.B2(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_45),
.A2(n_41),
.B1(n_31),
.B2(n_32),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_109),
.B1(n_116),
.B2(n_88),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g109 ( 
.A1(n_54),
.A2(n_31),
.B1(n_27),
.B2(n_15),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_23),
.B1(n_31),
.B2(n_41),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_72),
.A2(n_31),
.B1(n_27),
.B2(n_3),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_27),
.B1(n_1),
.B2(n_3),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_52),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_43),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_47),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_59),
.A2(n_7),
.B1(n_8),
.B2(n_82),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_132),
.B1(n_99),
.B2(n_118),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_62),
.A2(n_7),
.B1(n_68),
.B2(n_81),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_74),
.A2(n_48),
.B1(n_67),
.B2(n_46),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g175 ( 
.A1(n_134),
.A2(n_96),
.B1(n_133),
.B2(n_131),
.Y(n_175)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_135),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_136),
.B(n_137),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_105),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_61),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_138),
.B(n_139),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_126),
.C(n_90),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_139),
.C(n_145),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_141),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_173),
.B1(n_162),
.B2(n_150),
.Y(n_199)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_144),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_157),
.Y(n_181)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_147),
.B(n_149),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_104),
.A2(n_108),
.B1(n_116),
.B2(n_119),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_148),
.A2(n_149),
.B1(n_169),
.B2(n_167),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_134),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_162),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_103),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_154),
.Y(n_183)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_103),
.B(n_87),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_93),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_156),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_113),
.B(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_87),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_107),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_99),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_150),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_102),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_102),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_172),
.Y(n_216)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_131),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_175),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_96),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_177),
.Y(n_218)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_88),
.B(n_112),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_137),
.C(n_165),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_186),
.B(n_164),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_188),
.A2(n_192),
.B1(n_199),
.B2(n_151),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_157),
.B1(n_175),
.B2(n_142),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_191),
.A2(n_218),
.B1(n_209),
.B2(n_205),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_171),
.B1(n_176),
.B2(n_174),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_136),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_207),
.Y(n_230)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_144),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_196),
.B(n_210),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_180),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_160),
.Y(n_207)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_146),
.B(n_162),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_212),
.B(n_217),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_135),
.B(n_143),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_172),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_161),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_219),
.A2(n_244),
.B(n_246),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_222),
.C(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_226),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_181),
.B(n_186),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_227),
.Y(n_253)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_178),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_189),
.B1(n_195),
.B2(n_202),
.Y(n_260)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_232),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_141),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_234),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_181),
.B(n_141),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_184),
.B(n_141),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_235),
.B(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_185),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_182),
.B(n_166),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_165),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_239),
.B(n_251),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_242),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_196),
.B1(n_199),
.B2(n_192),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_245),
.B1(n_214),
.B2(n_201),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_200),
.B1(n_207),
.B2(n_212),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_195),
.B1(n_202),
.B2(n_208),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_183),
.B(n_197),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_206),
.A2(n_198),
.B(n_205),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_198),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_194),
.B(n_187),
.Y(n_249)
);

AOI221xp5_ASAP7_75t_L g267 ( 
.A1(n_249),
.A2(n_250),
.B1(n_193),
.B2(n_203),
.C(n_201),
.Y(n_267)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_254),
.B(n_261),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_193),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_262),
.C(n_270),
.Y(n_287)
);

INVxp67_ASAP7_75t_SL g283 ( 
.A(n_260),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_222),
.B(n_189),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_208),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_264),
.A2(n_271),
.B1(n_248),
.B2(n_227),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_219),
.A2(n_214),
.B(n_203),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_265),
.A2(n_269),
.B(n_278),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_267),
.A2(n_265),
.B1(n_263),
.B2(n_266),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_241),
.B(n_230),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_268),
.A2(n_247),
.B(n_221),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_193),
.B(n_214),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_220),
.B(n_201),
.C(n_244),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_243),
.A2(n_250),
.B1(n_230),
.B2(n_223),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_242),
.B(n_226),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_238),
.C(n_239),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_224),
.A2(n_236),
.B(n_232),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_284),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_233),
.B1(n_224),
.B2(n_245),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_293),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_273),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_235),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_286),
.B(n_290),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_257),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_240),
.Y(n_290)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_291),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_255),
.A2(n_228),
.B1(n_229),
.B2(n_225),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_292),
.A2(n_263),
.B1(n_264),
.B2(n_276),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_297),
.B(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_266),
.A2(n_237),
.B1(n_249),
.B2(n_251),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_299),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_256),
.A2(n_237),
.B(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_274),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_315),
.Y(n_325)
);

A2O1A1O1Ixp25_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_270),
.B(n_254),
.C(n_276),
.D(n_257),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_319),
.B(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_285),
.B(n_258),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_301),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_261),
.C(n_262),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_317),
.C(n_287),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_314),
.A2(n_283),
.B1(n_296),
.B2(n_277),
.Y(n_335)
);

OA21x2_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_272),
.B(n_252),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_271),
.C(n_275),
.Y(n_317)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_269),
.B(n_252),
.Y(n_319)
);

OAI322xp33_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_237),
.A3(n_260),
.B1(n_277),
.B2(n_288),
.C1(n_287),
.C2(n_300),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_297),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_337),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_303),
.A2(n_294),
.B(n_302),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_326),
.A2(n_322),
.B(n_307),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_L g348 ( 
.A1(n_327),
.A2(n_331),
.B(n_338),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_282),
.C(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_311),
.C(n_314),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_289),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_330),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_289),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_308),
.B(n_292),
.Y(n_331)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_332),
.B(n_334),
.Y(n_342)
);

INVx13_ASAP7_75t_L g333 ( 
.A(n_313),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_333),
.Y(n_347)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_306),
.B1(n_303),
.B2(n_316),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_320),
.A2(n_319),
.B1(n_306),
.B2(n_316),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_318),
.B1(n_304),
.B2(n_312),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_294),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_345),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_349),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_315),
.C(n_304),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_344),
.B(n_324),
.C(n_326),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_318),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_350),
.A2(n_351),
.B1(n_335),
.B2(n_330),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_331),
.A2(n_308),
.B1(n_321),
.B2(n_260),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_352),
.B(n_357),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_327),
.C(n_325),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_353),
.B(n_356),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_354),
.A2(n_358),
.B1(n_351),
.B2(n_341),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_349),
.B(n_332),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_336),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_323),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_325),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_361),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_342),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_338),
.B1(n_340),
.B2(n_346),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_362),
.B(n_367),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_260),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_360),
.B(n_348),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_339),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_329),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_350),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_345),
.B(n_355),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_366),
.B(n_359),
.C(n_353),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_373),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_371),
.A2(n_374),
.B1(n_369),
.B2(n_333),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g376 ( 
.A(n_372),
.B(n_365),
.C(n_364),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_376),
.B(n_362),
.C(n_373),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_334),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_378),
.B(n_379),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_380),
.B(n_375),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_321),
.Y(n_382)
);


endmodule