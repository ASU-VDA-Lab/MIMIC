module fake_jpeg_20094_n_74 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_22;
wire n_40;
wire n_73;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_67;
wire n_56;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;
wire n_70;
wire n_66;

BUFx10_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_5),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_24),
.A2(n_9),
.B1(n_18),
.B2(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_31),
.B1(n_33),
.B2(n_29),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_32),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_48),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_61),
.B1(n_57),
.B2(n_35),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_42),
.C(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_65),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_59),
.B1(n_53),
.B2(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_62),
.Y(n_68)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_52),
.B1(n_56),
.B2(n_54),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_69),
.C(n_30),
.Y(n_71)
);

OAI31xp33_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_32),
.A3(n_22),
.B(n_70),
.Y(n_72)
);

XNOR2x2_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_51),
.Y(n_74)
);


endmodule