module fake_jpeg_9121_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_65),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_42),
.B1(n_45),
.B2(n_40),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_67),
.B1(n_72),
.B2(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_68),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_51),
.B1(n_49),
.B2(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_9),
.B(n_11),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_75),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_39),
.B1(n_50),
.B2(n_5),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_25),
.B1(n_37),
.B2(n_7),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_44),
.B1(n_4),
.B2(n_3),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_4),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_8),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_89),
.A2(n_79),
.B1(n_83),
.B2(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_83),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_85),
.B1(n_84),
.B2(n_87),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_88),
.C(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_80),
.C(n_86),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_95),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_24),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_26),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_29),
.C(n_30),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_31),
.B(n_32),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_33),
.Y(n_102)
);


endmodule