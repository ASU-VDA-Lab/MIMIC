module fake_jpeg_27385_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_16),
.B(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_65),
.Y(n_76)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_44),
.B1(n_25),
.B2(n_28),
.Y(n_81)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx2_ASAP7_75t_SL g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_24),
.B1(n_32),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_62),
.A2(n_26),
.B1(n_19),
.B2(n_25),
.Y(n_108)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_24),
.B1(n_16),
.B2(n_31),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_29),
.B1(n_31),
.B2(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_35),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_39),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_82),
.Y(n_140)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_48),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_80),
.B(n_34),
.C(n_43),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_81),
.A2(n_93),
.B1(n_100),
.B2(n_108),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_46),
.B1(n_45),
.B2(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_84),
.B1(n_59),
.B2(n_54),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_46),
.B1(n_45),
.B2(n_41),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_21),
.B1(n_26),
.B2(n_28),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_35),
.Y(n_124)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_37),
.B1(n_47),
.B2(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_101),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_47),
.B1(n_19),
.B2(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_31),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_50),
.A2(n_19),
.B1(n_23),
.B2(n_22),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_110),
.B1(n_61),
.B2(n_53),
.Y(n_120)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_50),
.A2(n_28),
.B1(n_34),
.B2(n_22),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_60),
.Y(n_137)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_47),
.B1(n_22),
.B2(n_23),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_113),
.A2(n_34),
.B1(n_23),
.B2(n_25),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_43),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_49),
.C(n_75),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_115),
.A2(n_116),
.B1(n_121),
.B2(n_126),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_135),
.C(n_138),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_119),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_61),
.B1(n_49),
.B2(n_43),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_139),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_131),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_49),
.B1(n_30),
.B2(n_18),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_79),
.B(n_14),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_60),
.C(n_30),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_87),
.B(n_27),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_82),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_97),
.A2(n_30),
.B1(n_18),
.B2(n_27),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_144),
.A2(n_114),
.B1(n_108),
.B2(n_81),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_107),
.B1(n_94),
.B2(n_78),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_158),
.B1(n_142),
.B2(n_128),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_80),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_159),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_93),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_165),
.B(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_157),
.Y(n_181)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_80),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_76),
.Y(n_163)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_166),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_105),
.B(n_92),
.C(n_90),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_106),
.B1(n_104),
.B2(n_109),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_178),
.B1(n_126),
.B2(n_116),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_169),
.Y(n_210)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_86),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_114),
.B1(n_113),
.B2(n_100),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_172),
.A2(n_175),
.B1(n_176),
.B2(n_119),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_85),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_1),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_139),
.A2(n_105),
.B1(n_107),
.B2(n_89),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_127),
.A2(n_98),
.B1(n_112),
.B2(n_111),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_77),
.B1(n_99),
.B2(n_89),
.Y(n_176)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_77),
.B(n_91),
.C(n_102),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_102),
.B1(n_30),
.B2(n_3),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_188),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_131),
.B1(n_144),
.B2(n_121),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_182),
.A2(n_201),
.B(n_207),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_184),
.A2(n_187),
.B1(n_206),
.B2(n_157),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_168),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_117),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_186),
.B(n_195),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_151),
.A2(n_125),
.B1(n_142),
.B2(n_136),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_190),
.B1(n_196),
.B2(n_197),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_119),
.A3(n_128),
.B1(n_136),
.B2(n_145),
.C1(n_102),
.C2(n_141),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_141),
.B1(n_133),
.B2(n_118),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_118),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_158),
.A2(n_118),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_205),
.B1(n_156),
.B2(n_152),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_208),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_14),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_173),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_151),
.A2(n_14),
.B1(n_5),
.B2(n_6),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_153),
.A2(n_1),
.B(n_6),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_156),
.A2(n_6),
.B(n_7),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_148),
.B(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_212),
.B(n_227),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_214),
.B(n_208),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_187),
.C(n_146),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_225),
.C(n_214),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_217),
.A2(n_220),
.B1(n_234),
.B2(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_198),
.B1(n_180),
.B2(n_183),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_162),
.B1(n_159),
.B2(n_166),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_223),
.B1(n_193),
.B2(n_207),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_209),
.A2(n_170),
.B1(n_164),
.B2(n_154),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_192),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_226),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_146),
.C(n_147),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_183),
.A2(n_169),
.B(n_147),
.Y(n_228)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_228),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_150),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_176),
.B1(n_8),
.B2(n_9),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_188),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_7),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_8),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_243),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_227),
.B1(n_197),
.B2(n_200),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_191),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_245),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_256),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_235),
.B(n_189),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_253),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_235),
.B(n_225),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_228),
.C(n_230),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_258),
.C(n_259),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_215),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_182),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_218),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_201),
.C(n_203),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_201),
.C(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_222),
.B(n_237),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_267),
.A2(n_271),
.B(n_260),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_206),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_282),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_231),
.C(n_229),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_272),
.C(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_237),
.B(n_238),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_232),
.C(n_220),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_280),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_254),
.C(n_253),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_218),
.B1(n_226),
.B2(n_213),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_279),
.A2(n_13),
.B1(n_10),
.B2(n_11),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_257),
.B(n_213),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_193),
.C(n_205),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_255),
.C(n_240),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_211),
.Y(n_282)
);

AOI21x1_ASAP7_75t_SL g285 ( 
.A1(n_282),
.A2(n_250),
.B(n_252),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_274),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_296),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_247),
.C(n_246),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_295),
.C(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_255),
.C(n_261),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_266),
.B(n_236),
.C(n_234),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_8),
.C(n_9),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_275),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g299 ( 
.A1(n_286),
.A2(n_281),
.B(n_277),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_299),
.A2(n_301),
.B(n_284),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_311),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_269),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_303),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_280),
.B1(n_273),
.B2(n_274),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_9),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_297),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_273),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_10),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_11),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_312),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_310),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_316),
.Y(n_324)
);

INVx11_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_12),
.B1(n_13),
.B2(n_318),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_285),
.B(n_287),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_306),
.C(n_288),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_308),
.C(n_306),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_12),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_317),
.C(n_315),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_314),
.A2(n_287),
.B1(n_309),
.B2(n_13),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_319),
.B(n_11),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_312),
.B(n_316),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_324),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_327),
.C(n_321),
.Y(n_332)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_323),
.B(n_324),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_333),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_328),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_320),
.B(n_315),
.Y(n_339)
);


endmodule