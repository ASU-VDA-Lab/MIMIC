module fake_jpeg_24971_n_167 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_68),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_75),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_63),
.B1(n_61),
.B2(n_53),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_54),
.B1(n_58),
.B2(n_55),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_70),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_63),
.B1(n_47),
.B2(n_49),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_48),
.B1(n_72),
.B2(n_67),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_88),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_71),
.A3(n_49),
.B1(n_50),
.B2(n_59),
.Y(n_91)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_87),
.CI(n_18),
.CON(n_117),
.SN(n_117)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_98),
.B1(n_104),
.B2(n_107),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_100),
.Y(n_110)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_68),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_102),
.A2(n_87),
.B1(n_88),
.B2(n_52),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_64),
.B1(n_62),
.B2(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_68),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_48),
.B1(n_57),
.B2(n_52),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_102),
.B1(n_97),
.B2(n_90),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_0),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_20),
.B(n_43),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_115),
.A2(n_90),
.B(n_17),
.Y(n_120)
);

NOR2x1_ASAP7_75t_R g118 ( 
.A(n_117),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_121),
.Y(n_140)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_117),
.A2(n_93),
.B(n_106),
.C(n_27),
.D(n_30),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_120),
.B(n_123),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_125),
.B1(n_114),
.B2(n_115),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_2),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_126),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_15),
.B1(n_41),
.B2(n_40),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_3),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_3),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_127),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_135),
.B1(n_139),
.B2(n_137),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_112),
.B1(n_4),
.B2(n_5),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_14),
.C(n_38),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_42),
.C(n_36),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_11),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_141),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_22),
.B(n_37),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_148),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_146),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_152),
.B1(n_138),
.B2(n_136),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_132),
.A2(n_33),
.B(n_32),
.C(n_31),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_153),
.A2(n_145),
.B1(n_150),
.B2(n_143),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_156),
.C(n_155),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_143),
.B1(n_152),
.B2(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_144),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_134),
.C(n_142),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_147),
.B1(n_142),
.B2(n_29),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_165),
.B(n_7),
.Y(n_166)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_8),
.CON(n_167),
.SN(n_167)
);


endmodule