module real_aes_7039_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_109), .C(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g440 ( .A(n_0), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_1), .A2(n_145), .B(n_150), .C(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_2), .A2(n_140), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g458 ( .A(n_3), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_4), .B(n_164), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g719 ( .A1(n_5), .A2(n_15), .B1(n_720), .B2(n_721), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_5), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g475 ( .A1(n_6), .A2(n_140), .B(n_476), .Y(n_475) );
AND2x6_ASAP7_75t_L g145 ( .A(n_7), .B(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g174 ( .A(n_8), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_9), .B(n_43), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_9), .B(n_43), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_10), .A2(n_252), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_11), .B(n_155), .Y(n_191) );
INVx1_ASAP7_75t_L g480 ( .A(n_12), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_13), .B(n_154), .Y(n_528) );
INVx1_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g720 ( .A(n_15), .Y(n_720) );
INVx1_ASAP7_75t_L g540 ( .A(n_16), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g199 ( .A1(n_17), .A2(n_175), .B(n_200), .C(n_202), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_18), .B(n_164), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_19), .B(n_469), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_20), .B(n_140), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_21), .B(n_260), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_22), .A2(n_154), .B(n_156), .C(n_160), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_23), .B(n_164), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_24), .B(n_155), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_25), .A2(n_158), .B(n_202), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_26), .B(n_155), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_27), .Y(n_220) );
INVx1_ASAP7_75t_L g234 ( .A(n_28), .Y(n_234) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_29), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_30), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_31), .B(n_155), .Y(n_459) );
INVx1_ASAP7_75t_L g257 ( .A(n_32), .Y(n_257) );
INVx1_ASAP7_75t_L g493 ( .A(n_33), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_34), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g143 ( .A(n_35), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_36), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_37), .A2(n_154), .B(n_213), .C(n_215), .Y(n_212) );
INVxp67_ASAP7_75t_L g258 ( .A(n_38), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g211 ( .A(n_39), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g232 ( .A1(n_40), .A2(n_150), .B(n_233), .C(n_239), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_41), .A2(n_145), .B(n_150), .C(n_508), .Y(n_507) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_42), .A2(n_92), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_42), .Y(n_124) );
INVx1_ASAP7_75t_L g492 ( .A(n_44), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_45), .A2(n_172), .B(n_173), .C(n_176), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_46), .B(n_155), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_47), .A2(n_121), .B1(n_433), .B2(n_434), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_47), .Y(n_433) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_48), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_49), .Y(n_254) );
INVx1_ASAP7_75t_L g148 ( .A(n_50), .Y(n_148) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_51), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_52), .B(n_140), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_53), .A2(n_150), .B1(n_160), .B2(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_54), .A2(n_104), .B1(n_113), .B2(n_732), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_55), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_56), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g170 ( .A(n_57), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_58), .A2(n_172), .B(n_215), .C(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_59), .Y(n_521) );
INVx1_ASAP7_75t_L g477 ( .A(n_60), .Y(n_477) );
INVx1_ASAP7_75t_L g146 ( .A(n_61), .Y(n_146) );
INVx1_ASAP7_75t_L g137 ( .A(n_62), .Y(n_137) );
INVx1_ASAP7_75t_SL g214 ( .A(n_63), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_65), .B(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g223 ( .A(n_66), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_SL g468 ( .A1(n_67), .A2(n_215), .B(n_469), .C(n_470), .Y(n_468) );
INVxp67_ASAP7_75t_L g471 ( .A(n_68), .Y(n_471) );
INVx1_ASAP7_75t_L g112 ( .A(n_69), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_70), .A2(n_140), .B(n_169), .Y(n_168) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_71), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_72), .A2(n_140), .B(n_197), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_73), .Y(n_496) );
INVx1_ASAP7_75t_L g515 ( .A(n_74), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_75), .A2(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g198 ( .A(n_76), .Y(n_198) );
CKINVDCx16_ASAP7_75t_R g231 ( .A(n_77), .Y(n_231) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_78), .A2(n_446), .B1(n_717), .B2(n_723), .C1(n_727), .C2(n_728), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g516 ( .A1(n_79), .A2(n_145), .B(n_150), .C(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_80), .A2(n_140), .B(n_147), .Y(n_139) );
INVx1_ASAP7_75t_L g201 ( .A(n_81), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_82), .B(n_235), .Y(n_509) );
INVx2_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx1_ASAP7_75t_L g188 ( .A(n_84), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_85), .B(n_469), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_86), .A2(n_145), .B(n_150), .C(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g109 ( .A(n_87), .Y(n_109) );
OR2x2_ASAP7_75t_L g437 ( .A(n_87), .B(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g716 ( .A(n_87), .B(n_439), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_88), .A2(n_150), .B(n_222), .C(n_225), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_89), .A2(n_718), .B1(n_719), .B2(n_722), .Y(n_717) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_89), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_90), .B(n_167), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_91), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_92), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_93), .A2(n_145), .B(n_150), .C(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_94), .Y(n_532) );
INVx1_ASAP7_75t_L g467 ( .A(n_95), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_96), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_97), .B(n_235), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_98), .B(n_133), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_99), .B(n_133), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_100), .B(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g157 ( .A(n_101), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_102), .A2(n_140), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g732 ( .A(n_106), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g715 ( .A(n_109), .B(n_439), .Y(n_715) );
NOR2x2_ASAP7_75t_L g730 ( .A(n_109), .B(n_438), .Y(n_730) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_444), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g731 ( .A(n_116), .Y(n_731) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_435), .B(n_442), .Y(n_119) );
INVx1_ASAP7_75t_L g434 ( .A(n_121), .Y(n_434) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_431), .B2(n_432), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_122), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_125), .A2(n_715), .B1(n_724), .B2(n_725), .Y(n_723) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g432 ( .A(n_126), .Y(n_432) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_357), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_299), .C(n_329), .D(n_339), .Y(n_127) );
OAI211xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_204), .B(n_262), .C(n_289), .Y(n_128) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_129), .A2(n_304), .B1(n_385), .B2(n_386), .C1(n_387), .C2(n_388), .Y(n_384) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_179), .Y(n_129) );
AOI33xp33_ASAP7_75t_L g310 ( .A1(n_130), .A2(n_297), .A3(n_298), .B1(n_311), .B2(n_316), .B3(n_318), .Y(n_310) );
OAI211xp5_ASAP7_75t_SL g367 ( .A1(n_130), .A2(n_368), .B(n_370), .C(n_372), .Y(n_367) );
OR2x2_ASAP7_75t_L g383 ( .A(n_130), .B(n_369), .Y(n_383) );
INVx1_ASAP7_75t_L g416 ( .A(n_130), .Y(n_416) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_166), .Y(n_130) );
INVx2_ASAP7_75t_L g293 ( .A(n_131), .Y(n_293) );
AND2x2_ASAP7_75t_L g309 ( .A(n_131), .B(n_195), .Y(n_309) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_131), .Y(n_344) );
AND2x2_ASAP7_75t_L g373 ( .A(n_131), .B(n_166), .Y(n_373) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_139), .B(n_163), .Y(n_131) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_132), .A2(n_196), .B(n_203), .Y(n_195) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_132), .A2(n_209), .B(n_217), .Y(n_208) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx4_ASAP7_75t_L g165 ( .A(n_133), .Y(n_165) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_133), .A2(n_465), .B(n_472), .Y(n_464) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g250 ( .A(n_134), .Y(n_250) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_135), .B(n_136), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
BUFx2_ASAP7_75t_L g252 ( .A(n_140), .Y(n_252) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_141), .B(n_145), .Y(n_185) );
AND2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx1_ASAP7_75t_L g238 ( .A(n_142), .Y(n_238) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g151 ( .A(n_143), .Y(n_151) );
INVx1_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx1_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
INVx3_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx1_ASAP7_75t_L g469 ( .A(n_144), .Y(n_469) );
INVx4_ASAP7_75t_SL g162 ( .A(n_145), .Y(n_162) );
BUFx3_ASAP7_75t_L g239 ( .A(n_145), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_SL g147 ( .A1(n_148), .A2(n_149), .B(n_153), .C(n_162), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_SL g169 ( .A1(n_149), .A2(n_162), .B(n_170), .C(n_171), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g197 ( .A1(n_149), .A2(n_162), .B(n_198), .C(n_199), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_149), .A2(n_162), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_149), .A2(n_162), .B(n_254), .C(n_255), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_149), .A2(n_162), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_149), .A2(n_162), .B(n_477), .C(n_478), .Y(n_476) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_149), .A2(n_162), .B(n_537), .C(n_538), .Y(n_536) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x6_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
BUFx3_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_151), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_154), .B(n_214), .Y(n_213) );
INVx4_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g172 ( .A(n_155), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_158), .B(n_201), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_158), .A2(n_235), .B1(n_257), .B2(n_258), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_158), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g190 ( .A(n_159), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g491 ( .A1(n_159), .A2(n_190), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx2_ASAP7_75t_L g460 ( .A(n_160), .Y(n_460) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_162), .A2(n_185), .B1(n_490), .B2(n_494), .Y(n_489) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_164), .A2(n_475), .B(n_481), .Y(n_474) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_165), .B(n_194), .Y(n_193) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_219), .B(n_226), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_165), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_165), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g273 ( .A(n_166), .Y(n_273) );
BUFx3_ASAP7_75t_L g281 ( .A(n_166), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_166), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g292 ( .A(n_166), .B(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_166), .B(n_180), .Y(n_321) );
AND2x2_ASAP7_75t_L g390 ( .A(n_166), .B(n_324), .Y(n_390) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_178), .Y(n_166) );
INVx1_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
INVx2_ASAP7_75t_L g228 ( .A(n_167), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_L g230 ( .A1(n_167), .A2(n_185), .B(n_231), .C(n_232), .Y(n_230) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_167), .A2(n_535), .B(n_541), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
INVx5_ASAP7_75t_L g235 ( .A(n_175), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_175), .B(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_175), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g192 ( .A(n_176), .Y(n_192) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g202 ( .A(n_177), .Y(n_202) );
INVx2_ASAP7_75t_SL g284 ( .A(n_179), .Y(n_284) );
OR2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_195), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_180), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g326 ( .A(n_180), .Y(n_326) );
AND2x2_ASAP7_75t_L g337 ( .A(n_180), .B(n_293), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_180), .B(n_322), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_180), .B(n_324), .Y(n_369) );
AND2x2_ASAP7_75t_L g428 ( .A(n_180), .B(n_373), .Y(n_428) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g298 ( .A(n_181), .B(n_195), .Y(n_298) );
AND2x2_ASAP7_75t_L g308 ( .A(n_181), .B(n_309), .Y(n_308) );
BUFx3_ASAP7_75t_L g330 ( .A(n_181), .Y(n_330) );
AND3x2_ASAP7_75t_L g389 ( .A(n_181), .B(n_390), .C(n_391), .Y(n_389) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_193), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_182), .B(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_182), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_182), .B(n_532), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_185), .A2(n_220), .B(n_221), .Y(n_219) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_185), .A2(n_455), .B(n_456), .Y(n_454) );
OAI21xp5_ASAP7_75t_L g514 ( .A1(n_185), .A2(n_515), .B(n_516), .Y(n_514) );
O2A1O1Ixp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_191), .C(n_192), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_189), .A2(n_192), .B(n_223), .C(n_224), .Y(n_222) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_192), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_192), .A2(n_518), .B(n_519), .Y(n_517) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
INVx1_ASAP7_75t_SL g324 ( .A(n_195), .Y(n_324) );
NAND3xp33_ASAP7_75t_L g336 ( .A(n_195), .B(n_273), .C(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_242), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_205), .A2(n_308), .B(n_360), .C(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_207), .B(n_229), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_207), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_SL g376 ( .A(n_207), .Y(n_376) );
AND2x2_ASAP7_75t_L g397 ( .A(n_207), .B(n_244), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_207), .B(n_306), .Y(n_425) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AND2x2_ASAP7_75t_L g270 ( .A(n_208), .B(n_261), .Y(n_270) );
INVx2_ASAP7_75t_L g277 ( .A(n_208), .Y(n_277) );
AND2x2_ASAP7_75t_L g297 ( .A(n_208), .B(n_244), .Y(n_297) );
AND2x2_ASAP7_75t_L g347 ( .A(n_208), .B(n_229), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_208), .Y(n_351) );
INVx3_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_216), .Y(n_529) );
INVx2_ASAP7_75t_SL g261 ( .A(n_218), .Y(n_261) );
BUFx2_ASAP7_75t_L g287 ( .A(n_218), .Y(n_287) );
AND2x2_ASAP7_75t_L g414 ( .A(n_218), .B(n_229), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g260 ( .A(n_228), .Y(n_260) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_228), .A2(n_524), .B(n_531), .Y(n_523) );
INVx3_ASAP7_75t_SL g244 ( .A(n_229), .Y(n_244) );
AND2x2_ASAP7_75t_L g269 ( .A(n_229), .B(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g276 ( .A(n_229), .B(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g306 ( .A(n_229), .B(n_266), .Y(n_306) );
OR2x2_ASAP7_75t_L g315 ( .A(n_229), .B(n_261), .Y(n_315) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_229), .Y(n_333) );
AND2x2_ASAP7_75t_L g338 ( .A(n_229), .B(n_291), .Y(n_338) );
AND2x2_ASAP7_75t_L g366 ( .A(n_229), .B(n_246), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_229), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g404 ( .A(n_229), .B(n_245), .Y(n_404) );
OR2x6_ASAP7_75t_L g229 ( .A(n_230), .B(n_240), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .C(n_237), .Y(n_233) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_235), .A2(n_458), .B(n_459), .C(n_460), .Y(n_457) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_238), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x2_ASAP7_75t_L g328 ( .A(n_244), .B(n_277), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_244), .B(n_270), .Y(n_356) );
AND2x2_ASAP7_75t_L g374 ( .A(n_244), .B(n_291), .Y(n_374) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_261), .Y(n_245) );
AND2x2_ASAP7_75t_L g275 ( .A(n_246), .B(n_261), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_246), .B(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g313 ( .A(n_246), .Y(n_313) );
OR2x2_ASAP7_75t_L g361 ( .A(n_246), .B(n_281), .Y(n_361) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_251), .B(n_259), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_248), .A2(n_267), .B(n_268), .Y(n_266) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_248), .A2(n_514), .B(n_520), .Y(n_513) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AOI21xp5_ASAP7_75t_SL g505 ( .A1(n_249), .A2(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_250), .A2(n_454), .B(n_461), .Y(n_453) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_250), .A2(n_489), .B(n_495), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_250), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_259), .Y(n_268) );
AND2x2_ASAP7_75t_L g296 ( .A(n_261), .B(n_266), .Y(n_296) );
INVx1_ASAP7_75t_L g304 ( .A(n_261), .Y(n_304) );
AND2x2_ASAP7_75t_L g399 ( .A(n_261), .B(n_277), .Y(n_399) );
AOI222xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_271), .B1(n_274), .B2(n_278), .C1(n_282), .C2(n_285), .Y(n_262) );
INVx1_ASAP7_75t_L g394 ( .A(n_263), .Y(n_394) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_269), .Y(n_263) );
AND2x2_ASAP7_75t_L g290 ( .A(n_264), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g301 ( .A(n_264), .B(n_270), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_264), .B(n_292), .Y(n_317) );
OAI222xp33_ASAP7_75t_L g339 ( .A1(n_264), .A2(n_340), .B1(n_345), .B2(n_346), .C1(n_354), .C2(n_356), .Y(n_339) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g327 ( .A(n_266), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_266), .B(n_347), .Y(n_387) );
AND2x2_ASAP7_75t_L g398 ( .A(n_266), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g406 ( .A(n_269), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_271), .B(n_322), .Y(n_385) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_273), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g343 ( .A(n_273), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx3_ASAP7_75t_L g288 ( .A(n_276), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_276), .A2(n_379), .B(n_382), .C(n_384), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_276), .B(n_313), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_276), .B(n_296), .Y(n_418) );
AND2x2_ASAP7_75t_L g291 ( .A(n_277), .B(n_287), .Y(n_291) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g318 ( .A(n_280), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g307 ( .A(n_281), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g370 ( .A(n_281), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g409 ( .A(n_281), .B(n_309), .Y(n_409) );
INVx1_ASAP7_75t_L g421 ( .A(n_281), .Y(n_421) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_284), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g402 ( .A(n_287), .Y(n_402) );
A2O1A1Ixp33_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_292), .B(n_294), .C(n_298), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_290), .A2(n_320), .B1(n_335), .B2(n_338), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_291), .B(n_305), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_291), .B(n_313), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_292), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_SL g355 ( .A(n_292), .Y(n_355) );
AND2x2_ASAP7_75t_L g362 ( .A(n_292), .B(n_342), .Y(n_362) );
INVx2_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NOR4xp25_ASAP7_75t_L g300 ( .A(n_297), .B(n_301), .C(n_302), .D(n_305), .Y(n_300) );
INVx1_ASAP7_75t_SL g371 ( .A(n_298), .Y(n_371) );
AND2x2_ASAP7_75t_L g415 ( .A(n_298), .B(n_416), .Y(n_415) );
OAI211xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_307), .B(n_310), .C(n_319), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_306), .B(n_376), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_308), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_426) );
INVx1_ASAP7_75t_SL g381 ( .A(n_309), .Y(n_381) );
AND2x2_ASAP7_75t_L g420 ( .A(n_309), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_313), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_317), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_318), .B(n_343), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_325), .B(n_327), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g395 ( .A(n_322), .Y(n_395) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g423 ( .A(n_323), .Y(n_423) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
OAI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B(n_334), .Y(n_329) );
CKINVDCx16_ASAP7_75t_R g342 ( .A(n_330), .Y(n_342) );
OR2x2_ASAP7_75t_L g380 ( .A(n_330), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_333), .A2(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_337), .A2(n_364), .B1(n_367), .B2(n_374), .C(n_375), .Y(n_363) );
INVx1_ASAP7_75t_SL g407 ( .A(n_338), .Y(n_407) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OR2x2_ASAP7_75t_L g354 ( .A(n_342), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g391 ( .A(n_344), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_351), .B2(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_350), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR4xp25_ASAP7_75t_L g357 ( .A(n_358), .B(n_392), .C(n_405), .D(n_417), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g358 ( .A(n_359), .B(n_363), .C(n_378), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_361), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_368), .B(n_373), .Y(n_377) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI221xp5_ASAP7_75t_SL g405 ( .A1(n_380), .A2(n_406), .B1(n_407), .B2(n_408), .C(n_410), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_L g396 ( .A1(n_382), .A2(n_397), .B(n_398), .C(n_400), .Y(n_396) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_383), .A2(n_401), .B1(n_403), .B2(n_404), .Y(n_400) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B(n_395), .C(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g411 ( .A(n_404), .Y(n_411) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI221xp5_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_432), .A2(n_447), .B1(n_715), .B2(n_716), .Y(n_446) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g443 ( .A(n_437), .Y(n_443) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AOI21xp33_ASAP7_75t_SL g444 ( .A1(n_442), .A2(n_445), .B(n_731), .Y(n_444) );
INVx1_ASAP7_75t_L g724 ( .A(n_447), .Y(n_724) );
NAND2x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_631), .Y(n_447) );
NOR5xp2_ASAP7_75t_L g448 ( .A(n_449), .B(n_554), .C(n_586), .D(n_601), .E(n_618), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_482), .B(n_501), .C(n_542), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_463), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_451), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_451), .B(n_606), .Y(n_669) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_452), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_452), .B(n_498), .Y(n_555) );
AND2x2_ASAP7_75t_L g596 ( .A(n_452), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_452), .B(n_565), .Y(n_600) );
OR2x2_ASAP7_75t_L g637 ( .A(n_452), .B(n_488), .Y(n_637) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g487 ( .A(n_453), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g545 ( .A(n_453), .Y(n_545) );
OR2x2_ASAP7_75t_L g708 ( .A(n_453), .B(n_548), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_463), .A2(n_611), .B1(n_612), .B2(n_615), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_463), .B(n_545), .Y(n_694) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_473), .Y(n_463) );
AND2x2_ASAP7_75t_L g500 ( .A(n_464), .B(n_488), .Y(n_500) );
AND2x2_ASAP7_75t_L g547 ( .A(n_464), .B(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g552 ( .A(n_464), .Y(n_552) );
INVx3_ASAP7_75t_L g565 ( .A(n_464), .Y(n_565) );
OR2x2_ASAP7_75t_L g585 ( .A(n_464), .B(n_548), .Y(n_585) );
AND2x2_ASAP7_75t_L g604 ( .A(n_464), .B(n_474), .Y(n_604) );
BUFx2_ASAP7_75t_L g636 ( .A(n_464), .Y(n_636) );
AND2x4_ASAP7_75t_L g551 ( .A(n_473), .B(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g486 ( .A(n_474), .Y(n_486) );
INVx2_ASAP7_75t_L g499 ( .A(n_474), .Y(n_499) );
OR2x2_ASAP7_75t_L g567 ( .A(n_474), .B(n_548), .Y(n_567) );
AND2x2_ASAP7_75t_L g597 ( .A(n_474), .B(n_488), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_474), .B(n_545), .Y(n_614) );
AND2x2_ASAP7_75t_L g654 ( .A(n_474), .B(n_565), .Y(n_654) );
AND2x2_ASAP7_75t_SL g690 ( .A(n_474), .B(n_500), .Y(n_690) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_484), .B(n_497), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g668 ( .A(n_485), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g628 ( .A1(n_486), .A2(n_500), .B(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_486), .B(n_488), .Y(n_684) );
AND2x2_ASAP7_75t_L g620 ( .A(n_487), .B(n_621), .Y(n_620) );
INVx3_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_488), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_497), .B(n_545), .Y(n_713) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_498), .A2(n_656), .B1(n_657), .B2(n_662), .Y(n_655) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x2_ASAP7_75t_L g546 ( .A(n_499), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g584 ( .A(n_499), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g621 ( .A(n_499), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_500), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g675 ( .A(n_500), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_522), .Y(n_502) );
INVx4_ASAP7_75t_L g561 ( .A(n_503), .Y(n_561) );
AND2x2_ASAP7_75t_L g639 ( .A(n_503), .B(n_606), .Y(n_639) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_513), .Y(n_503) );
INVx3_ASAP7_75t_L g558 ( .A(n_504), .Y(n_558) );
AND2x2_ASAP7_75t_L g572 ( .A(n_504), .B(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g576 ( .A(n_504), .Y(n_576) );
INVx2_ASAP7_75t_L g590 ( .A(n_504), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_504), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g647 ( .A(n_504), .B(n_642), .Y(n_647) );
AND2x2_ASAP7_75t_L g712 ( .A(n_504), .B(n_682), .Y(n_712) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_511), .Y(n_504) );
AND2x2_ASAP7_75t_L g553 ( .A(n_513), .B(n_534), .Y(n_553) );
INVx2_ASAP7_75t_L g573 ( .A(n_513), .Y(n_573) );
INVx1_ASAP7_75t_L g578 ( .A(n_522), .Y(n_578) );
AND2x2_ASAP7_75t_L g624 ( .A(n_522), .B(n_572), .Y(n_624) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_533), .Y(n_522) );
INVx2_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_523), .B(n_573), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g606 ( .A(n_533), .B(n_563), .Y(n_606) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g559 ( .A(n_534), .Y(n_559) );
AND2x2_ASAP7_75t_L g642 ( .A(n_534), .B(n_573), .Y(n_642) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_549), .B(n_553), .Y(n_542) );
INVx1_ASAP7_75t_SL g587 ( .A(n_543), .Y(n_587) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_544), .B(n_551), .Y(n_644) );
INVx1_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g593 ( .A(n_545), .B(n_548), .Y(n_593) );
AND2x2_ASAP7_75t_L g622 ( .A(n_545), .B(n_566), .Y(n_622) );
OR2x2_ASAP7_75t_L g625 ( .A(n_545), .B(n_585), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_546), .A2(n_638), .B1(n_690), .B2(n_691), .C1(n_693), .C2(n_695), .Y(n_689) );
BUFx2_ASAP7_75t_L g603 ( .A(n_548), .Y(n_603) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g592 ( .A(n_551), .B(n_593), .Y(n_592) );
INVx3_ASAP7_75t_SL g609 ( .A(n_551), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_551), .B(n_603), .Y(n_663) );
AND2x2_ASAP7_75t_L g598 ( .A(n_553), .B(n_558), .Y(n_598) );
INVx1_ASAP7_75t_L g617 ( .A(n_553), .Y(n_617) );
OAI221xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_556), .B1(n_560), .B2(n_564), .C(n_568), .Y(n_554) );
OR2x2_ASAP7_75t_L g626 ( .A(n_556), .B(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
AND2x2_ASAP7_75t_L g611 ( .A(n_558), .B(n_581), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_558), .B(n_571), .Y(n_651) );
AND2x2_ASAP7_75t_L g656 ( .A(n_558), .B(n_606), .Y(n_656) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_558), .Y(n_666) );
NAND2x1_ASAP7_75t_SL g677 ( .A(n_558), .B(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g562 ( .A(n_559), .B(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g582 ( .A(n_559), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_559), .B(n_577), .Y(n_608) );
INVx1_ASAP7_75t_L g674 ( .A(n_559), .Y(n_674) );
INVx1_ASAP7_75t_L g649 ( .A(n_560), .Y(n_649) );
OR2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g661 ( .A(n_561), .Y(n_661) );
NOR2xp67_ASAP7_75t_L g673 ( .A(n_561), .B(n_674), .Y(n_673) );
INVx2_ASAP7_75t_L g678 ( .A(n_562), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_562), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g581 ( .A(n_563), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_563), .B(n_573), .Y(n_594) );
INVx1_ASAP7_75t_L g660 ( .A(n_563), .Y(n_660) );
INVx1_ASAP7_75t_L g681 ( .A(n_564), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OAI21xp5_ASAP7_75t_SL g568 ( .A1(n_569), .A2(n_574), .B(n_583), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g714 ( .A(n_570), .B(n_647), .Y(n_714) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g682 ( .A(n_571), .B(n_642), .Y(n_682) );
AOI32xp33_ASAP7_75t_L g595 ( .A1(n_572), .A2(n_578), .A3(n_596), .B1(n_598), .B2(n_599), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g697 ( .A1(n_572), .A2(n_604), .A3(n_687), .B1(n_698), .B2(n_699), .C1(n_700), .C2(n_702), .Y(n_697) );
INVx2_ASAP7_75t_L g577 ( .A(n_573), .Y(n_577) );
INVx1_ASAP7_75t_L g687 ( .A(n_573), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_575), .B(n_581), .Y(n_630) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_576), .B(n_642), .Y(n_692) );
INVx1_ASAP7_75t_L g579 ( .A(n_577), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_577), .B(n_606), .Y(n_696) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_585), .B(n_680), .Y(n_679) );
OAI221xp5_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_588), .B1(n_591), .B2(n_594), .C(n_595), .Y(n_586) );
OR2x2_ASAP7_75t_L g607 ( .A(n_588), .B(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g616 ( .A(n_588), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g641 ( .A(n_589), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g645 ( .A(n_599), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_605), .B1(n_607), .B2(n_609), .C(n_610), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_603), .A2(n_634), .B1(n_638), .B2(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_604), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_604), .Y(n_709) );
INVx1_ASAP7_75t_L g703 ( .A(n_606), .Y(n_703) );
INVx1_ASAP7_75t_SL g638 ( .A(n_607), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_609), .B(n_637), .Y(n_699) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_614), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g680 ( .A(n_614), .Y(n_680) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_623), .B1(n_625), .B2(n_626), .C(n_628), .Y(n_618) );
NOR2xp33_ASAP7_75t_SL g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_620), .A2(n_638), .B1(n_684), .B2(n_685), .Y(n_683) );
CKINVDCx14_ASAP7_75t_R g623 ( .A(n_624), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_625), .A2(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR3xp33_ASAP7_75t_SL g631 ( .A(n_632), .B(n_664), .C(n_688), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_633), .B(n_640), .C(n_648), .D(n_655), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g711 ( .A(n_636), .Y(n_711) );
INVx3_ASAP7_75t_SL g705 ( .A(n_637), .Y(n_705) );
OR2x2_ASAP7_75t_L g710 ( .A(n_637), .B(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_643), .B1(n_645), .B2(n_647), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_642), .B(n_660), .Y(n_701) );
INVxp67_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_650), .B(n_652), .Y(n_648) );
INVxp67_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_665), .A2(n_667), .B(n_670), .C(n_683), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g698 ( .A(n_669), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B1(n_676), .B2(n_679), .C1(n_681), .C2(n_682), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND4xp25_ASAP7_75t_SL g707 ( .A(n_680), .B(n_708), .C(n_709), .D(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND3xp33_ASAP7_75t_SL g688 ( .A(n_689), .B(n_697), .C(n_706), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_712), .B1(n_713), .B2(n_714), .Y(n_706) );
INVx1_ASAP7_75t_L g726 ( .A(n_716), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_717), .Y(n_727) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
endmodule