module real_jpeg_16452_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_553;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_632),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_0),
.B(n_633),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_1),
.A2(n_113),
.B1(n_313),
.B2(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_1),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_1),
.A2(n_374),
.B1(n_432),
.B2(n_436),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_1),
.A2(n_374),
.B1(n_547),
.B2(n_550),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_1),
.A2(n_374),
.B1(n_608),
.B2(n_609),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_47),
.B1(n_54),
.B2(n_56),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_2),
.A2(n_56),
.B1(n_68),
.B2(n_71),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_2),
.A2(n_56),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_2),
.A2(n_56),
.B1(n_293),
.B2(n_298),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_3),
.Y(n_230)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_3),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g364 ( 
.A(n_3),
.Y(n_364)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_5),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_5),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_119),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

AOI22x1_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_119),
.B1(n_252),
.B2(n_258),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_5),
.A2(n_119),
.B1(n_366),
.B2(n_368),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_6),
.B(n_353),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_6),
.A2(n_352),
.B(n_353),
.Y(n_418)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_6),
.Y(n_453)
);

OAI32xp33_ASAP7_75t_L g495 ( 
.A1(n_6),
.A2(n_150),
.A3(n_496),
.B1(n_501),
.B2(n_503),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_6),
.A2(n_415),
.B1(n_453),
.B2(n_537),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_6),
.B(n_158),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_6),
.A2(n_227),
.B1(n_607),
.B2(n_610),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_7),
.A2(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_7),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_7),
.A2(n_116),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_7),
.A2(n_116),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_7),
.A2(n_116),
.B1(n_298),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_8),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_8),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g569 ( 
.A(n_8),
.Y(n_569)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_8),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_9),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_9),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_9),
.A2(n_266),
.B1(n_339),
.B2(n_342),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_9),
.A2(n_266),
.B1(n_285),
.B2(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_9),
.A2(n_266),
.B1(n_507),
.B2(n_510),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_10),
.A2(n_376),
.B1(n_378),
.B2(n_379),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_10),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_10),
.A2(n_378),
.B1(n_411),
.B2(n_415),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_10),
.A2(n_378),
.B1(n_527),
.B2(n_530),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g590 ( 
.A1(n_10),
.A2(n_378),
.B1(n_591),
.B2(n_593),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_11),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g297 ( 
.A(n_11),
.Y(n_297)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_11),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_12),
.Y(n_633)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_13),
.A2(n_173),
.B1(n_176),
.B2(n_179),
.Y(n_172)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_13),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_13),
.A2(n_179),
.B1(n_316),
.B2(n_319),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_SL g388 ( 
.A1(n_13),
.A2(n_179),
.B1(n_389),
.B2(n_392),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_13),
.A2(n_179),
.B1(n_442),
.B2(n_447),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_14),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_62),
.B1(n_105),
.B2(n_108),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_62),
.B1(n_148),
.B2(n_152),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_14),
.A2(n_62),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_15),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_15),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_15),
.A2(n_310),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_15),
.A2(n_310),
.B1(n_485),
.B2(n_489),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_15),
.A2(n_310),
.B1(n_368),
.B2(n_554),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_17),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_17),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_17),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_17),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_17),
.Y(n_257)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_17),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_17),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g175 ( 
.A(n_19),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_19),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_162),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_160),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_24),
.B(n_63),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_24)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_25),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_25),
.A2(n_46),
.B1(n_57),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_25),
.A2(n_57),
.B1(n_112),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_25),
.A2(n_57),
.B1(n_172),
.B2(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_25),
.A2(n_57),
.B1(n_263),
.B2(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_25),
.A2(n_57),
.B1(n_373),
.B2(n_375),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_25),
.A2(n_57),
.B1(n_307),
.B2(n_375),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_25),
.A2(n_57),
.B1(n_373),
.B2(n_418),
.Y(n_417)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B(n_41),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AO22x2_ASAP7_75t_L g41 ( 
.A1(n_29),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_35),
.A2(n_187),
.B1(n_346),
.B2(n_351),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_36),
.Y(n_353)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_37),
.Y(n_265)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_111),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_42),
.Y(n_186)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_42),
.Y(n_435)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_43),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_44),
.Y(n_337)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_45),
.Y(n_349)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2x1_ASAP7_75t_R g452 ( 
.A(n_57),
.B(n_453),
.Y(n_452)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_60),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_155),
.C(n_157),
.Y(n_63)
);

FAx1_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_155),
.CI(n_157),
.CON(n_165),
.SN(n_165)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_110),
.C(n_122),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_65),
.A2(n_66),
.B1(n_122),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22x1_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_76),
.B1(n_104),
.B2(n_109),
.Y(n_66)
);

OAI22x1_ASAP7_75t_L g183 ( 
.A1(n_67),
.A2(n_76),
.B1(n_109),
.B2(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_73),
.Y(n_334)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_73),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_75),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_75),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_75),
.Y(n_343)
);

OAI22x1_ASAP7_75t_SL g314 ( 
.A1(n_76),
.A2(n_109),
.B1(n_214),
.B2(n_315),
.Y(n_314)
);

OAI22x1_ASAP7_75t_L g400 ( 
.A1(n_76),
.A2(n_109),
.B1(n_315),
.B2(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_76),
.A2(n_109),
.B1(n_410),
.B2(n_416),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_76),
.A2(n_109),
.B1(n_410),
.B2(n_431),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_76),
.A2(n_109),
.B1(n_431),
.B2(n_536),
.Y(n_535)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_77),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_77),
.A2(n_158),
.B1(n_213),
.B2(n_223),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_77),
.A2(n_158),
.B1(n_331),
.B2(n_338),
.Y(n_330)
);

OA21x2_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_93),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_83),
.Y(n_415)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_85),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_90),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_100),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_99),
.Y(n_261)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_107),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_107),
.Y(n_350)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_109),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_114),
.Y(n_309)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_115),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_122),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_122),
.B(n_182),
.C(n_183),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_183),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_137),
.B(n_147),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_123),
.A2(n_137),
.B1(n_147),
.B2(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_123),
.B(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_123),
.A2(n_137),
.B1(n_281),
.B2(n_388),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_123),
.A2(n_137),
.B1(n_484),
.B2(n_526),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_123),
.A2(n_137),
.B1(n_526),
.B2(n_546),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_123),
.A2(n_137),
.B1(n_546),
.B2(n_581),
.Y(n_580)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_124),
.A2(n_205),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_124),
.A2(n_250),
.B1(n_420),
.B2(n_423),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_124),
.A2(n_250),
.B1(n_420),
.B2(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_124),
.B(n_453),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.B1(n_131),
.B2(n_133),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_130),
.Y(n_242)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_130),
.Y(n_246)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_130),
.Y(n_367)
);

INVx5_ASAP7_75t_L g451 ( 
.A(n_130),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_130),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_130),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_131),
.Y(n_593)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_131),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_132),
.Y(n_302)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_137),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_137),
.B(n_281),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B1(n_142),
.B2(n_144),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_140),
.Y(n_393)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_145),
.Y(n_422)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_151),
.Y(n_211)
);

BUFx12f_ASAP7_75t_L g286 ( 
.A(n_151),
.Y(n_286)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_152),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_154),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_188),
.B(n_630),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_165),
.B(n_166),
.Y(n_631)
);

BUFx24_ASAP7_75t_SL g634 ( 
.A(n_165),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_171),
.C(n_180),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_171),
.B1(n_182),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_171),
.A2(n_182),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_175),
.Y(n_377)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_177),
.Y(n_380)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_325),
.B(n_627),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_269),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g627 ( 
.A1(n_192),
.A2(n_628),
.B(n_629),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_193),
.B(n_196),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.C(n_224),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_198),
.A2(n_201),
.B1(n_202),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_198),
.Y(n_324)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_202),
.A2(n_203),
.B(n_212),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_212),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_217),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_217),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_224),
.B(n_323),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_247),
.B(n_262),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_225),
.A2(n_226),
.B1(n_262),
.B2(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_225),
.A2(n_226),
.B1(n_249),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_239),
.Y(n_226)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_227),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_227),
.A2(n_355),
.B1(n_362),
.B2(n_365),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_227),
.A2(n_292),
.B1(n_365),
.B2(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_227),
.A2(n_234),
.B1(n_553),
.B2(n_557),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_227),
.A2(n_514),
.B1(n_590),
.B2(n_607),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

INVx6_ASAP7_75t_L g304 ( 
.A(n_228),
.Y(n_304)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_229),
.Y(n_515)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_230),
.Y(n_397)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_235),
.A2(n_290),
.B1(n_356),
.B2(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_237),
.Y(n_605)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_247),
.A2(n_248),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_249),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_256),
.Y(n_533)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_256),
.Y(n_583)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_257),
.Y(n_492)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_261),
.Y(n_391)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_262),
.Y(n_275)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_322),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_270),
.B(n_322),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_276),
.C(n_278),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_272),
.B(n_277),
.Y(n_470)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_278),
.B(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_306),
.C(n_314),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_279),
.B(n_464),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_287),
.B(n_289),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_280),
.B(n_287),
.Y(n_383)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_284),
.Y(n_529)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_286),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_289),
.B(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_303),
.B2(n_305),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_290),
.A2(n_441),
.B1(n_506),
.B2(n_512),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_290),
.A2(n_512),
.B1(n_589),
.B2(n_594),
.Y(n_588)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_296),
.Y(n_556)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_297),
.Y(n_370)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_300),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_302),
.Y(n_446)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_306),
.B(n_314),
.Y(n_464)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_473),
.B(n_622),
.Y(n_325)
);

NAND3xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_456),
.C(n_468),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_402),
.B(n_424),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_328),
.B(n_402),
.C(n_624),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_381),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_329),
.B(n_382),
.C(n_384),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_344),
.C(n_371),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_330),
.A2(n_371),
.B1(n_372),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_331),
.Y(n_416)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_343),
.Y(n_438)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_343),
.Y(n_500)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_343),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_354),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_345),
.B(n_354),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_357),
.Y(n_609)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_360),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_364),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_370),
.Y(n_592)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_398),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_394),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_386),
.A2(n_387),
.B1(n_394),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_388),
.Y(n_423)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_400),
.C(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.C(n_408),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_403),
.B(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_406),
.B(n_408),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_417),
.C(n_419),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_419),
.Y(n_427)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_417),
.B(n_427),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_454),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_425),
.B(n_454),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_428),
.C(n_429),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_426),
.B(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_428),
.B(n_429),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_439),
.C(n_452),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_430),
.B(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_439),
.A2(n_440),
.B1(n_452),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OAI32xp33_ASAP7_75t_L g566 ( 
.A1(n_448),
.A2(n_528),
.A3(n_567),
.B1(n_570),
.B2(n_572),
.Y(n_566)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_452),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_453),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_453),
.B(n_571),
.Y(n_570)
);

OAI21xp33_ASAP7_75t_SL g581 ( 
.A1(n_453),
.A2(n_570),
.B(n_582),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_453),
.B(n_603),
.Y(n_602)
);

A2O1A1O1Ixp25_ASAP7_75t_L g622 ( 
.A1(n_456),
.A2(n_468),
.B(n_623),
.C(n_625),
.D(n_626),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_467),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_457),
.B(n_467),
.Y(n_625)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.Y(n_457)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_463),
.B1(n_465),
.B2(n_466),
.Y(n_460)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_461),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_461),
.B(n_466),
.C(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_463),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_469),
.B(n_471),
.Y(n_626)
);

AOI21x1_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_516),
.B(n_621),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_477),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_475),
.B(n_477),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_482),
.C(n_493),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_478),
.A2(n_479),
.B1(n_519),
.B2(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_482),
.A2(n_493),
.B1(n_494),
.B2(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_482),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx5_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_504),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_495),
.A2(n_504),
.B1(n_505),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_495),
.Y(n_524)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_506),
.Y(n_557)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_541),
.B(n_620),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_SL g517 ( 
.A(n_518),
.B(n_522),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_518),
.B(n_522),
.Y(n_620)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.C(n_534),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_523),
.B(n_561),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_525),
.A2(n_534),
.B1(n_535),
.B2(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_525),
.Y(n_562)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

AOI21x1_ASAP7_75t_SL g541 ( 
.A1(n_542),
.A2(n_563),
.B(n_619),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_560),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_543),
.B(n_560),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_552),
.C(n_558),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_544),
.A2(n_545),
.B1(n_558),
.B2(n_559),
.Y(n_585)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_548),
.Y(n_551)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_552),
.B(n_585),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_553),
.Y(n_594)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

OAI21x1_ASAP7_75t_SL g563 ( 
.A1(n_564),
.A2(n_586),
.B(n_618),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_584),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_565),
.B(n_584),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_579),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_566),
.A2(n_579),
.B1(n_580),
.B2(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_566),
.Y(n_596)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_577),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx8_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_597),
.B(n_617),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_595),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_595),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_598),
.A2(n_613),
.B(n_616),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_599),
.B(n_606),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_602),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_614),
.B(n_615),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_614),
.B(n_615),
.Y(n_616)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);


endmodule