module fake_jpeg_27246_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_14),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_19),
.A2(n_3),
.B(n_4),
.Y(n_26)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_23),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_21),
.C(n_20),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_13),
.C(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_27),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_22),
.B1(n_12),
.B2(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_34),
.B1(n_22),
.B2(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_10),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_16),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.C(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_46),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_31),
.C(n_36),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_35),
.C(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_49),
.A2(n_41),
.B(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_51),
.A2(n_15),
.B1(n_11),
.B2(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_55),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_50),
.B1(n_48),
.B2(n_13),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_62),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_60),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_60),
.B(n_6),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_54),
.C(n_58),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_13),
.B(n_16),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_4),
.C(n_7),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.C(n_8),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_13),
.B(n_71),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_13),
.Y(n_73)
);


endmodule