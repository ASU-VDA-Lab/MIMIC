module fake_jpeg_19507_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_32),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_3),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_14),
.B(n_4),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_39),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_15),
.C(n_14),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_29),
.B1(n_31),
.B2(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_51),
.B1(n_54),
.B2(n_59),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_12),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_50),
.B(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_22),
.B1(n_17),
.B2(n_21),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_18),
.B(n_16),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_44),
.B(n_42),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_17),
.B1(n_21),
.B2(n_12),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_16),
.B(n_24),
.C(n_14),
.D(n_15),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_11),
.B1(n_0),
.B2(n_5),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_14),
.B(n_15),
.C(n_20),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_49),
.B1(n_41),
.B2(n_19),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_66),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_68),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_4),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_60),
.B(n_61),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_75),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_78),
.B(n_41),
.C(n_49),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_64),
.Y(n_79)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_73),
.C(n_75),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_69),
.B1(n_41),
.B2(n_20),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_87),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_79),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_95),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_80),
.C(n_76),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_94),
.A2(n_89),
.B(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_95),
.B(n_63),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_98),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_96),
.C(n_7),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_99),
.B1(n_7),
.B2(n_8),
.Y(n_102)
);


endmodule