module fake_netlist_6_2523_n_106 (n_7, n_6, n_12, n_4, n_2, n_15, n_16, n_3, n_5, n_1, n_14, n_13, n_0, n_9, n_11, n_8, n_17, n_10, n_106);

input n_7;
input n_6;
input n_12;
input n_4;
input n_2;
input n_15;
input n_16;
input n_3;
input n_5;
input n_1;
input n_14;
input n_13;
input n_0;
input n_9;
input n_11;
input n_8;
input n_17;
input n_10;

output n_106;

wire n_52;
wire n_91;
wire n_46;
wire n_18;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_19;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

AND2x4_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_1),
.Y(n_43)
);

NAND2x1p5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_23),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_31),
.B1(n_43),
.B2(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_48),
.B1(n_44),
.B2(n_51),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_48),
.B(n_38),
.C(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_44),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_29),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_42),
.B1(n_58),
.B2(n_54),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_58),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_54),
.B(n_30),
.C(n_26),
.Y(n_69)
);

AOI221xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_34),
.B1(n_27),
.B2(n_25),
.C(n_30),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_28),
.B1(n_44),
.B2(n_48),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_61),
.B1(n_48),
.B2(n_39),
.Y(n_72)
);

OAI222xp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_66),
.B1(n_67),
.B2(n_26),
.C1(n_41),
.C2(n_69),
.Y(n_73)
);

OAI211xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_67),
.B(n_66),
.C(n_41),
.Y(n_74)
);

OAI31xp33_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_32),
.A3(n_52),
.B(n_45),
.Y(n_75)
);

AOI221xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_52),
.B1(n_32),
.B2(n_50),
.C(n_53),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_74),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_46),
.C(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

OAI221xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_50),
.B1(n_57),
.B2(n_46),
.C(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_82),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_81),
.B1(n_73),
.B2(n_46),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

NAND4xp75_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_75),
.C(n_3),
.D(n_5),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_91),
.Y(n_93)
);

NAND2x1_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_86),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_84),
.B(n_87),
.Y(n_95)
);

AOI221xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_92),
.B1(n_89),
.B2(n_10),
.C(n_8),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_92),
.B(n_10),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_9),
.B1(n_49),
.B2(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_49),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_11),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_49),
.B(n_57),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_49),
.B(n_57),
.Y(n_106)
);


endmodule