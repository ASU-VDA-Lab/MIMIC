module fake_jpeg_12229_n_118 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_118);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.C(n_1),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_29),
.A2(n_40),
.B(n_48),
.C(n_34),
.Y(n_69)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_5),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_14),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_36),
.B(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2x1p5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_10),
.B(n_27),
.C(n_20),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_20),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_13),
.B1(n_15),
.B2(n_43),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_56),
.B1(n_70),
.B2(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_69),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_37),
.B1(n_35),
.B2(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_46),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_33),
.B(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_30),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_59),
.B1(n_71),
.B2(n_67),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_81),
.B(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_53),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_87),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_62),
.C(n_61),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_88),
.C(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_52),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_68),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_69),
.A2(n_56),
.B(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_57),
.C(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_59),
.B1(n_76),
.B2(n_71),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_105),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_102),
.B1(n_92),
.B2(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_78),
.B1(n_88),
.B2(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_107),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_73),
.C(n_94),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_89),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_112),
.C(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_114),
.A2(n_115),
.B1(n_97),
.B2(n_98),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_107),
.C(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_95),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_117),
.B(n_101),
.Y(n_118)
);


endmodule