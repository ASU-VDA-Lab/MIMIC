module fake_jpeg_1124_n_441 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_13),
.B(n_11),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx2_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_51),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_52),
.B(n_59),
.Y(n_105)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_53),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_28),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_56),
.B(n_66),
.Y(n_115)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_61),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_28),
.B(n_13),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_80),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_15),
.B(n_7),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_88),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_85),
.B(n_86),
.Y(n_151)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_7),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_18),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_92),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_94),
.Y(n_141)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_96),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_98),
.Y(n_133)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_29),
.B1(n_24),
.B2(n_40),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_98),
.B1(n_81),
.B2(n_87),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_53),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_113),
.A2(n_154),
.B1(n_99),
.B2(n_138),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_78),
.A2(n_31),
.B1(n_47),
.B2(n_26),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_118),
.A2(n_119),
.B1(n_126),
.B2(n_2),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_72),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_54),
.A2(n_43),
.B1(n_34),
.B2(n_47),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_125),
.A2(n_127),
.B1(n_153),
.B2(n_89),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_62),
.A2(n_47),
.B1(n_43),
.B2(n_20),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_49),
.A2(n_34),
.B1(n_45),
.B2(n_39),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_20),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_142),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_30),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_68),
.B(n_30),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_60),
.B(n_15),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_76),
.B(n_24),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_152),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_40),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_58),
.A2(n_39),
.B1(n_27),
.B2(n_48),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_94),
.A2(n_26),
.B1(n_48),
.B2(n_27),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_84),
.B(n_46),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_156),
.Y(n_205)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_158),
.A2(n_185),
.B(n_192),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_164),
.Y(n_203)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_160),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_161),
.A2(n_177),
.B1(n_181),
.B2(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_162),
.Y(n_231)
);

AO22x1_ASAP7_75t_SL g163 ( 
.A1(n_118),
.A2(n_96),
.B1(n_85),
.B2(n_82),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_170),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_172),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_167),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_73),
.B1(n_75),
.B2(n_69),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_187),
.B1(n_198),
.B2(n_130),
.Y(n_211)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_0),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_0),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_178),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_0),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_107),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_188),
.B1(n_189),
.B2(n_199),
.Y(n_208)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_115),
.A2(n_70),
.B1(n_85),
.B2(n_82),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_96),
.C(n_32),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_191),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_105),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_183),
.B(n_194),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_190),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_35),
.B1(n_32),
.B2(n_5),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_113),
.A2(n_35),
.B1(n_9),
.B2(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_107),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_115),
.B(n_2),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_108),
.B(n_8),
.C(n_9),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_10),
.B(n_12),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_112),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_196),
.Y(n_227)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_197),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_133),
.A2(n_136),
.B1(n_138),
.B2(n_99),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_107),
.A2(n_137),
.B1(n_150),
.B2(n_114),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_100),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_135),
.B1(n_130),
.B2(n_146),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_202),
.A2(n_224),
.B1(n_219),
.B2(n_217),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g204 ( 
.A(n_175),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_193),
.A2(n_173),
.B1(n_170),
.B2(n_171),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_210),
.A2(n_215),
.B1(n_229),
.B2(n_234),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_211),
.A2(n_167),
.B1(n_103),
.B2(n_137),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_117),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_214),
.B(n_221),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_173),
.A2(n_128),
.B1(n_117),
.B2(n_104),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_159),
.A2(n_130),
.B1(n_104),
.B2(n_146),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_219),
.A2(n_222),
.B1(n_235),
.B2(n_179),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_136),
.C(n_150),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_164),
.A2(n_120),
.B1(n_146),
.B2(n_144),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_178),
.B(n_166),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_228),
.B(n_226),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_163),
.A2(n_116),
.B1(n_144),
.B2(n_129),
.Y(n_229)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_100),
.B(n_101),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_230),
.A2(n_101),
.B(n_103),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_163),
.A2(n_120),
.B1(n_144),
.B2(n_129),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_182),
.A2(n_129),
.B1(n_120),
.B2(n_149),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

NOR3xp33_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_174),
.C(n_188),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_238),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_239),
.A2(n_245),
.B1(n_251),
.B2(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_194),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_162),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_242),
.B(n_243),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_195),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_172),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_248),
.B(n_250),
.Y(n_289)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_205),
.Y(n_249)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_228),
.B(n_191),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_212),
.A2(n_185),
.B1(n_200),
.B2(n_196),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g286 ( 
.A(n_253),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_203),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_232),
.C(n_241),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_185),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_185),
.B1(n_160),
.B2(n_157),
.Y(n_257)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_186),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_259),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_210),
.B1(n_208),
.B2(n_211),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_122),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_261),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_220),
.B(n_122),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_235),
.Y(n_276)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_263),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_SL g264 ( 
.A1(n_206),
.A2(n_169),
.B(n_101),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_266),
.A2(n_207),
.B(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_267),
.A2(n_227),
.B1(n_213),
.B2(n_237),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_208),
.B1(n_230),
.B2(n_218),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_258),
.A2(n_202),
.B1(n_206),
.B2(n_214),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_271),
.A2(n_287),
.B1(n_292),
.B2(n_295),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_232),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_274),
.B(n_296),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_266),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_247),
.B(n_221),
.Y(n_277)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_277),
.B(n_250),
.CI(n_248),
.CON(n_314),
.SN(n_314)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_282),
.A2(n_267),
.B1(n_249),
.B2(n_252),
.Y(n_322)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_258),
.A2(n_222),
.B1(n_234),
.B2(n_229),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_288),
.A2(n_244),
.B(n_265),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_242),
.A2(n_233),
.B1(n_227),
.B2(n_216),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_233),
.B1(n_197),
.B2(n_225),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_247),
.B(n_207),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_298),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_288),
.B(n_291),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_299),
.B(n_310),
.Y(n_339)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_300),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_269),
.A2(n_280),
.B1(n_289),
.B2(n_279),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_301),
.A2(n_309),
.B1(n_316),
.B2(n_312),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_280),
.A2(n_251),
.B1(n_256),
.B2(n_255),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_303),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_292),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_311),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_271),
.A2(n_256),
.B1(n_264),
.B2(n_239),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_269),
.A2(n_256),
.B1(n_238),
.B2(n_257),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_257),
.B1(n_259),
.B2(n_243),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_296),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_289),
.A2(n_257),
.B1(n_262),
.B2(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_261),
.B(n_257),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_312),
.A2(n_283),
.B(n_274),
.Y(n_336)
);

A2O1A1O1Ixp25_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_293),
.B(n_286),
.C(n_209),
.D(n_237),
.Y(n_344)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_315),
.B(n_318),
.Y(n_338)
);

OAI22x1_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_291),
.B1(n_276),
.B2(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_290),
.B(n_263),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_293),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_320),
.Y(n_340)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_321),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_322),
.A2(n_307),
.B1(n_302),
.B2(n_303),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_323),
.A2(n_327),
.B1(n_342),
.B2(n_345),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_325),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_301),
.A2(n_279),
.B1(n_290),
.B2(n_281),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_318),
.B(n_246),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_328),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_272),
.Y(n_329)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_343),
.C(n_344),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_317),
.B(n_270),
.Y(n_335)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_335),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_336),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_277),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_346),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_341),
.A2(n_322),
.B1(n_321),
.B2(n_249),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_302),
.A2(n_286),
.B1(n_278),
.B2(n_273),
.Y(n_342)
);

XOR2x2_ASAP7_75t_L g343 ( 
.A(n_314),
.B(n_293),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_309),
.B(n_223),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_316),
.B(n_167),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_299),
.B(n_286),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_347),
.B(n_336),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_308),
.C(n_316),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_364),
.C(n_366),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_306),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_297),
.Y(n_356)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_297),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_359),
.B(n_360),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_311),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_253),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_314),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_363),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_327),
.B(n_305),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_347),
.B(n_304),
.C(n_320),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_331),
.A2(n_319),
.B1(n_298),
.B2(n_300),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_367),
.A2(n_369),
.B1(n_253),
.B2(n_252),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_358),
.A2(n_331),
.B1(n_341),
.B2(n_346),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_372),
.A2(n_367),
.B1(n_384),
.B2(n_378),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_362),
.B(n_339),
.Y(n_373)
);

NAND3xp33_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_348),
.C(n_369),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_339),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_375),
.A2(n_378),
.B1(n_386),
.B2(n_366),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_323),
.C(n_342),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_385),
.C(n_165),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_361),
.A2(n_344),
.B1(n_330),
.B2(n_326),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_358),
.A2(n_325),
.B(n_209),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_380),
.A2(n_384),
.B(n_131),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_383),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_176),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_253),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_355),
.A2(n_359),
.B(n_364),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_156),
.C(n_180),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_354),
.Y(n_387)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_379),
.B(n_357),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_388),
.B(n_394),
.Y(n_402)
);

OAI221xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_351),
.B1(n_360),
.B2(n_348),
.C(n_363),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_409)
);

NAND2xp33_ASAP7_75t_SL g403 ( 
.A(n_391),
.B(n_392),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_353),
.B(n_349),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_371),
.B(n_365),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_372),
.A2(n_349),
.B1(n_253),
.B2(n_176),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_397),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_399),
.Y(n_401)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_400),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_370),
.C(n_385),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_406),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_370),
.C(n_396),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_392),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_380),
.C(n_383),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_109),
.C(n_139),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_374),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_411),
.B(n_112),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_412),
.A2(n_400),
.B1(n_381),
.B2(n_389),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_413),
.B(n_415),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_389),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_414),
.B(n_420),
.Y(n_427)
);

AOI322xp5_ASAP7_75t_L g417 ( 
.A1(n_405),
.A2(n_403),
.A3(n_402),
.B1(n_409),
.B2(n_406),
.C1(n_410),
.C2(n_407),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_417),
.A2(n_418),
.B(n_422),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_401),
.A2(n_140),
.B(n_131),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_404),
.B(n_139),
.C(n_121),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_421),
.Y(n_429)
);

AOI21xp33_ASAP7_75t_L g422 ( 
.A1(n_401),
.A2(n_140),
.B(n_121),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_416),
.A2(n_140),
.B(n_121),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_423),
.A2(n_428),
.B(n_3),
.Y(n_433)
);

AOI31xp67_ASAP7_75t_L g424 ( 
.A1(n_419),
.A2(n_140),
.A3(n_10),
.B(n_12),
.Y(n_424)
);

O2A1O1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_424),
.A2(n_3),
.B(n_5),
.C(n_429),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_419),
.B(n_12),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_426),
.A2(n_418),
.B(n_121),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_430),
.B(n_431),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_426),
.A2(n_5),
.B(n_2),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_433),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_425),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_434),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_436),
.A2(n_427),
.B(n_3),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_438),
.A2(n_439),
.B(n_435),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_437),
.A2(n_3),
.B(n_5),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);


endmodule