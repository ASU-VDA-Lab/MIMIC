module fake_jpeg_15198_n_88 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_88);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_88;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_20),
.Y(n_25)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_22),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_22),
.A2(n_18),
.B1(n_13),
.B2(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_26),
.A2(n_31),
.B1(n_20),
.B2(n_19),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_9),
.B(n_17),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_15),
.B1(n_10),
.B2(n_12),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_22),
.A2(n_11),
.B1(n_16),
.B2(n_17),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_34),
.B1(n_32),
.B2(n_35),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_20),
.B1(n_19),
.B2(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_38),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_24),
.Y(n_36)
);

AOI31xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_26),
.A3(n_23),
.B(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_41),
.B1(n_25),
.B2(n_40),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_42),
.B1(n_36),
.B2(n_33),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_55),
.B1(n_44),
.B2(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_54),
.B(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_39),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_23),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_50),
.C(n_49),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_62),
.A2(n_57),
.B1(n_52),
.B2(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_61),
.C(n_65),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_57),
.B(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_68),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_73),
.C(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_68),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_14),
.A3(n_27),
.B1(n_30),
.B2(n_7),
.C1(n_4),
.C2(n_6),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_77),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_69),
.B(n_10),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_30),
.C(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_80),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_75),
.A2(n_4),
.B(n_8),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_27),
.C(n_6),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_0),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_1),
.B(n_2),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_81),
.C(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_86),
.B(n_3),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_84),
.Y(n_88)
);


endmodule