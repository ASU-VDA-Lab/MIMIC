module real_jpeg_4922_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_1),
.Y(n_87)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_3),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_4),
.B(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_5),
.Y(n_89)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_8),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_8),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_63),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_12),
.A2(n_40),
.B(n_62),
.Y(n_11)
);

OAI21xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_24),
.B(n_39),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_20),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_16),
.Y(n_14)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_35),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B(n_34),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_51),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_45),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_45),
.B(n_49),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_60),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_57),
.Y(n_61)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_61),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_96),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_83),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_90),
.B1(n_91),
.B2(n_95),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_86),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);


endmodule