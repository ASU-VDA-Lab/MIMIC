module fake_jpeg_25526_n_275 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_38),
.Y(n_44)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_54),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_46),
.B(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_36),
.B(n_26),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_17),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_15),
.C(n_28),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_58),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_79),
.B1(n_66),
.B2(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_62),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_23),
.B1(n_16),
.B2(n_26),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_65),
.B1(n_78),
.B2(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_49),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_23),
.B1(n_16),
.B2(n_21),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_35),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_18),
.B(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_18),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_17),
.C(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_23),
.B1(n_21),
.B2(n_30),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_62),
.A2(n_27),
.B(n_17),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_106),
.B(n_22),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_91),
.B(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_45),
.B1(n_50),
.B2(n_32),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_104),
.B1(n_107),
.B2(n_64),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_100),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_38),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_72),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_24),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_57),
.A2(n_66),
.B1(n_55),
.B2(n_76),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_80),
.B1(n_70),
.B2(n_64),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_35),
.C(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_10),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_32),
.B1(n_47),
.B2(n_20),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_27),
.B(n_22),
.C(n_19),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_47),
.B1(n_20),
.B2(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_77),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_74),
.C(n_67),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_96),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_71),
.B(n_0),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_126),
.B(n_98),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_106),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_120),
.Y(n_135)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_37),
.B(n_47),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_130),
.B(n_90),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_123),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx10_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_131),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_37),
.B1(n_48),
.B2(n_43),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_101),
.A2(n_38),
.B(n_19),
.Y(n_126)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_73),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_129),
.B1(n_94),
.B2(n_84),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_97),
.A2(n_22),
.B(n_19),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_100),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_146),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_141),
.B(n_142),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_91),
.B1(n_107),
.B2(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_84),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_153),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_132),
.B(n_126),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_145),
.B(n_155),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_86),
.B(n_96),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_150),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_157),
.B1(n_122),
.B2(n_52),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_111),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_93),
.B1(n_56),
.B2(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_160),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_105),
.B(n_93),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_89),
.B(n_73),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_131),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_29),
.B(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_158),
.B(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_120),
.B1(n_123),
.B2(n_121),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_176),
.B1(n_162),
.B2(n_152),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_119),
.B1(n_127),
.B2(n_122),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_174),
.A2(n_189),
.B1(n_149),
.B2(n_158),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_48),
.C(n_28),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_185),
.C(n_186),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_29),
.B(n_28),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_182),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_20),
.B1(n_29),
.B2(n_3),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_137),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_134),
.B(n_146),
.C(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_48),
.C(n_20),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_137),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_159),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_185),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_136),
.C(n_156),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_175),
.C(n_166),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_196),
.A2(n_172),
.B1(n_174),
.B2(n_187),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_175),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_205),
.B1(n_178),
.B2(n_165),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_155),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_204),
.Y(n_211)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_147),
.C(n_152),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_159),
.B1(n_138),
.B2(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_208),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_138),
.Y(n_209)
);

AO21x1_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_193),
.B(n_198),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_212),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_199),
.C(n_203),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_195),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_172),
.B(n_184),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_216),
.A2(n_202),
.B(n_204),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_183),
.B1(n_182),
.B2(n_171),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_166),
.C(n_177),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_222),
.B(n_190),
.C(n_212),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_173),
.B1(n_189),
.B2(n_7),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_196),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_217),
.C(n_211),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_230),
.B(n_233),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_231),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_191),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_194),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_238),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_173),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_213),
.B1(n_218),
.B2(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_245),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_247),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_235),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_210),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_248),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_220),
.B1(n_223),
.B2(n_211),
.C(n_8),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_4),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_4),
.C(n_5),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_255),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_231),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_257),
.C(n_249),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_261),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_254),
.A2(n_241),
.B(n_250),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_255),
.B(n_12),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_243),
.Y(n_261)
);

AOI32xp33_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_244),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_264),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_5),
.C(n_9),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_262),
.C(n_261),
.Y(n_268)
);

AOI321xp33_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_267),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_270),
.B(n_11),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_271),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_13),
.Y(n_275)
);


endmodule