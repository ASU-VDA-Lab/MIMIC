module real_jpeg_31090_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_0),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_0),
.Y(n_246)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_1),
.Y(n_320)
);

NAND2x1_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_2),
.B(n_162),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_2),
.B(n_349),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_2),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_2),
.B(n_429),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_2),
.B(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_3),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_3),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g312 ( 
.A(n_3),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_3),
.B(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_3),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_3),
.B(n_408),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_4),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_4),
.B(n_131),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_4),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_39),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_4),
.B(n_272),
.Y(n_271)
);

AND2x4_ASAP7_75t_SL g316 ( 
.A(n_4),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_4),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_5),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_5),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_5),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_5),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_6),
.B(n_245),
.Y(n_328)
);

NAND2x1p5_ASAP7_75t_L g391 ( 
.A(n_6),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_6),
.B(n_446),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_6),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_7),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_8),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_8),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_9),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_10),
.Y(n_125)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_10),
.Y(n_163)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_11),
.Y(n_80)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_11),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_12),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_12),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_12),
.B(n_39),
.Y(n_165)
);

AND2x4_ASAP7_75t_SL g283 ( 
.A(n_12),
.B(n_284),
.Y(n_283)
);

AND2x4_ASAP7_75t_SL g345 ( 
.A(n_12),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_12),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_12),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_13),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_13),
.B(n_49),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_13),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_13),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_13),
.B(n_34),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_13),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_14),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_14),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_14),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_14),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_14),
.B(n_49),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_14),
.B(n_330),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_540),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_15),
.B(n_541),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_16),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_16),
.B(n_268),
.Y(n_267)
);

NAND2x1_ASAP7_75t_L g321 ( 
.A(n_16),
.B(n_88),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_16),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_16),
.B(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_16),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_17),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_18),
.Y(n_347)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_18),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_19),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_19),
.B(n_327),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_19),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_19),
.B(n_433),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_19),
.B(n_92),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_485),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_362),
.B(n_482),
.Y(n_23)
);

AOI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_258),
.B(n_360),
.Y(n_24)
);

OAI21x1_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_169),
.B(n_256),
.Y(n_25)
);

NOR3xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_148),
.C(n_151),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_28),
.B(n_149),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_83),
.Y(n_28)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_29),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_29),
.B(n_358),
.C(n_359),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_53),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_30),
.B(n_54),
.C(n_65),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.C(n_47),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_31),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_155)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_36),
.Y(n_195)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_40),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_168)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_46),
.Y(n_530)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

OA21x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_60),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_59),
.Y(n_273)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_64),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_64),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_SL g337 ( 
.A(n_64),
.B(n_292),
.C(n_303),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_72),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_67),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_71),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_73),
.B(n_81),
.C(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_75),
.Y(n_219)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_76),
.Y(n_179)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_80),
.Y(n_270)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_84),
.B(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_127),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_85),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_101),
.C(n_115),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_87),
.B(n_91),
.C(n_96),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_89),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_95),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_95),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_95),
.Y(n_431)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_99),
.Y(n_216)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_99),
.Y(n_373)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_100),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_100),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_115),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_110),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_102),
.B(n_105),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_114),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_120),
.B1(n_121),
.B2(n_126),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_125),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_127),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_143),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_128),
.B(n_144),
.C(n_147),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_130),
.B(n_136),
.C(n_141),
.Y(n_302)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_141),
.B2(n_142),
.Y(n_134)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_144),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_151),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_166),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_152),
.B(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_154),
.B(n_167),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.C(n_159),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_156),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_161),
.B1(n_164),
.B2(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_251),
.B(n_255),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_210),
.B(n_250),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_198),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_172),
.B(n_198),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_191),
.C(n_197),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_173),
.A2(n_174),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_180),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_204),
.C(n_205),
.Y(n_203)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_185),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_192),
.B1(n_197),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_196),
.Y(n_213)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_195),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_197),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_202),
.B2(n_209),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_206),
.C(n_209),
.Y(n_252)
);

XOR2x1_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI21x1_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_224),
.B(n_249),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_SL g249 ( 
.A(n_212),
.B(n_220),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.C(n_217),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_232),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_233),
.B(n_248),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_226),
.B(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_230),
.Y(n_240)
);

BUFx4f_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_230),
.B(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_241),
.B(n_247),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_305),
.B(n_354),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_259),
.B(n_305),
.C(n_361),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_288),
.C(n_290),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_260),
.B(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_261),
.B(n_263),
.C(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_276),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g339 ( 
.A1(n_264),
.A2(n_271),
.B(n_275),
.C(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_267),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_267),
.B(n_274),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx3_ASAP7_75t_SL g404 ( 
.A(n_273),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_276),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_SL g455 ( 
.A(n_277),
.B(n_282),
.C(n_286),
.Y(n_455)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_283),
.C(n_287),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_287),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_289),
.B(n_291),
.Y(n_356)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_301),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_293),
.B(n_297),
.C(n_300),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_306),
.B(n_477),
.C(n_478),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_336),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_309),
.Y(n_478)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_322),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_321),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_311),
.B(n_321),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_312),
.Y(n_399)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_315),
.Y(n_378)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_316),
.Y(n_398)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_320),
.Y(n_515)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_321),
.B(n_398),
.C(n_399),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_321),
.B(n_398),
.C(n_399),
.Y(n_462)
);

XNOR2x1_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_323),
.Y(n_458)
);

AO22x1_ASAP7_75t_L g452 ( 
.A1(n_324),
.A2(n_453),
.B1(n_454),
.B2(n_458),
.Y(n_452)
);

OA22x2_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_329),
.B1(n_334),
.B2(n_335),
.Y(n_324)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_325),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_325),
.B(n_335),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_328),
.A2(n_385),
.B1(n_391),
.B2(n_394),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_328),
.B(n_388),
.C(n_391),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_328),
.B(n_388),
.C(n_391),
.Y(n_534)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_329),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_329),
.B(n_384),
.C(n_385),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_329),
.B(n_334),
.Y(n_456)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_336),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_R g470 ( 
.A(n_337),
.B(n_471),
.C(n_472),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_337),
.B(n_471),
.C(n_472),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_339),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_341),
.Y(n_472)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_342),
.B(n_345),
.C(n_465),
.Y(n_464)
);

OAI22x1_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_348),
.B2(n_353),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_348),
.Y(n_465)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_357),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_475),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_363),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_466),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_364),
.B(n_466),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_450),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_415),
.B1(n_448),
.B2(n_449),
.Y(n_365)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_395),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_367),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_383),
.C(n_386),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_369),
.B(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_374),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_379),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_379),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_379),
.B2(n_380),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_386),
.B(n_468),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_390),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_391),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_391),
.A2(n_394),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_394),
.B(n_437),
.C(n_444),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_405),
.B1(n_413),
.B2(n_414),
.Y(n_395)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_396),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.C(n_403),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_401),
.B1(n_403),
.B2(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_403),
.B(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_403),
.Y(n_461)
);

MAJx2_ASAP7_75t_L g533 ( 
.A(n_403),
.B(n_534),
.C(n_535),
.Y(n_533)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_405),
.Y(n_414)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

XOR2x1_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_412),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_407),
.Y(n_535)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_415),
.Y(n_491)
);

XOR2x1_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_435),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_421),
.Y(n_416)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_417),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_419),
.B(n_420),
.Y(n_417)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_421),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_427),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_423),
.B(n_502),
.C(n_503),
.Y(n_501)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_432),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_428),
.Y(n_502)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_432),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_436),
.B(n_518),
.C(n_519),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_436),
.B(n_518),
.C(n_519),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_443),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_444),
.A2(n_445),
.B1(n_506),
.B2(n_510),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_449),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_450),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_459),
.C(n_463),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_474),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.C(n_457),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_459),
.B(n_464),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_462),
.Y(n_459)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.C(n_473),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_479),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_479),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_537),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_492),
.Y(n_487)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_488),
.B(n_492),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.C(n_491),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.C(n_496),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_516),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_504),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_505),
.B(n_511),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_506),
.Y(n_510)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_520),
.B1(n_521),
.B2(n_536),
.Y(n_516)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_523),
.B1(n_532),
.B2(n_533),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

XOR2x1_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);

XNOR2x1_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_531),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);


endmodule