module fake_aes_11962_n_622 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_622);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_622;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_61), .Y(n_78) );
HB1xp67_ASAP7_75t_L g79 ( .A(n_72), .Y(n_79) );
BUFx5_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_67), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_17), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_58), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_12), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_10), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_36), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_25), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_45), .Y(n_89) );
INVx1_ASAP7_75t_SL g90 ( .A(n_74), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_41), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_73), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_27), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_53), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_24), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_65), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_29), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_11), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_37), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_16), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_9), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_64), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_55), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_60), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_52), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_63), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_11), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_69), .B(n_22), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_47), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_42), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_16), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_80), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_82), .A2(n_0), .B1(n_2), .B2(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_80), .Y(n_119) );
INVx4_ASAP7_75t_L g120 ( .A(n_115), .Y(n_120) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_83), .B(n_34), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_115), .B(n_0), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_80), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_79), .B(n_2), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_107), .B(n_3), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_84), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_104), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_101), .Y(n_130) );
CKINVDCx8_ASAP7_75t_R g131 ( .A(n_83), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_80), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_80), .Y(n_134) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_78), .A2(n_39), .B(n_76), .Y(n_135) );
INVxp33_ASAP7_75t_SL g136 ( .A(n_88), .Y(n_136) );
BUFx8_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
AND2x2_ASAP7_75t_SL g138 ( .A(n_78), .B(n_35), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_100), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_85), .B(n_4), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g141 ( .A1(n_102), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
OA21x2_ASAP7_75t_L g144 ( .A1(n_86), .A2(n_43), .B(n_75), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_107), .B(n_7), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_88), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_85), .B(n_8), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_87), .Y(n_148) );
OR2x2_ASAP7_75t_L g149 ( .A(n_120), .B(n_116), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_117), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_123), .B(n_108), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_137), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_120), .B(n_91), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
NAND3xp33_ASAP7_75t_L g156 ( .A(n_137), .B(n_93), .C(n_111), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_120), .B(n_103), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_122), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_123), .A2(n_116), .B1(n_102), .B2(n_103), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_146), .B(n_92), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_123), .A2(n_108), .B1(n_87), .B2(n_89), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_122), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_120), .B(n_94), .Y(n_164) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_138), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_146), .B(n_95), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_146), .B(n_92), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_137), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_140), .B(n_147), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_133), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_124), .Y(n_171) );
XNOR2xp5_ASAP7_75t_L g172 ( .A(n_118), .B(n_9), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_140), .A2(n_89), .B1(n_114), .B2(n_112), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_138), .A2(n_96), .B1(n_97), .B2(n_114), .Y(n_174) );
INVxp67_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_146), .B(n_136), .Y(n_176) );
OAI22xp33_ASAP7_75t_L g177 ( .A1(n_118), .A2(n_96), .B1(n_97), .B2(n_109), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_124), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_122), .Y(n_179) );
INVx5_ASAP7_75t_L g180 ( .A(n_122), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_122), .Y(n_181) );
AOI22xp5_ASAP7_75t_L g182 ( .A1(n_138), .A2(n_81), .B1(n_110), .B2(n_99), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_133), .B(n_106), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_127), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_139), .B(n_106), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_SL g187 ( .A1(n_176), .A2(n_126), .B(n_121), .C(n_148), .Y(n_187) );
INVxp67_ASAP7_75t_L g188 ( .A(n_175), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_154), .B(n_131), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_165), .A2(n_137), .B1(n_140), .B2(n_147), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_153), .B(n_131), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_174), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g193 ( .A1(n_172), .A2(n_129), .B1(n_141), .B2(n_125), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_167), .B(n_148), .Y(n_194) );
AND2x6_ASAP7_75t_SL g195 ( .A(n_186), .B(n_147), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_167), .B(n_143), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_165), .A2(n_147), .B1(n_140), .B2(n_143), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_157), .B(n_145), .Y(n_200) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_165), .A2(n_129), .B1(n_141), .B2(n_144), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_154), .Y(n_202) );
NAND2x1_ASAP7_75t_L g203 ( .A(n_169), .B(n_144), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_157), .B(n_119), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_174), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_170), .B(n_119), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_158), .Y(n_208) );
NOR3xp33_ASAP7_75t_L g209 ( .A(n_177), .B(n_90), .C(n_98), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_169), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_169), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_169), .Y(n_213) );
NOR2xp67_ASAP7_75t_L g214 ( .A(n_182), .B(n_10), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_153), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_182), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_170), .B(n_132), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_168), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_169), .A2(n_132), .B1(n_127), .B2(n_134), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g220 ( .A1(n_151), .A2(n_144), .B1(n_135), .B2(n_142), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_169), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_170), .B(n_134), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_168), .B(n_105), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_164), .B(n_142), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_151), .A2(n_142), .B1(n_130), .B2(n_113), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_169), .A2(n_142), .B1(n_130), .B2(n_135), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_149), .B(n_144), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_151), .A2(n_142), .B1(n_130), .B2(n_135), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_149), .B(n_142), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_152), .Y(n_231) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_152), .B(n_135), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_186), .B(n_130), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_162), .B(n_130), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_215), .B(n_160), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_214), .B(n_156), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_207), .A2(n_184), .B(n_166), .Y(n_238) );
O2A1O1Ixp5_ASAP7_75t_L g239 ( .A1(n_203), .A2(n_185), .B(n_161), .C(n_171), .Y(n_239) );
AOI21x1_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_185), .B(n_161), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_188), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_228), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_233), .A2(n_151), .B1(n_173), .B2(n_172), .Y(n_243) );
NOR2xp67_ASAP7_75t_L g244 ( .A(n_216), .B(n_12), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_199), .A2(n_151), .B1(n_150), .B2(n_171), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_189), .B(n_151), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_228), .Y(n_247) );
AOI21x1_ASAP7_75t_L g248 ( .A1(n_227), .A2(n_178), .B(n_150), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_192), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_189), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_202), .B(n_151), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_201), .A2(n_178), .B1(n_180), .B2(n_181), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_217), .A2(n_183), .B(n_181), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_222), .A2(n_183), .B(n_163), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_202), .A2(n_180), .B1(n_179), .B2(n_15), .Y(n_255) );
O2A1O1Ixp5_ASAP7_75t_L g256 ( .A1(n_235), .A2(n_180), .B(n_179), .C(n_48), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_218), .B(n_180), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_193), .A2(n_179), .B1(n_180), .B2(n_15), .C(n_17), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_218), .B(n_180), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
OR2x6_ASAP7_75t_SL g261 ( .A(n_206), .B(n_13), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_SL g262 ( .A1(n_226), .A2(n_179), .B(n_49), .C(n_50), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_206), .B(n_13), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_215), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_194), .A2(n_179), .B(n_51), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_231), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_196), .A2(n_14), .B(n_18), .C(n_20), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_227), .A2(n_46), .B(n_71), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_216), .B(n_14), .C(n_18), .Y(n_270) );
NOR2xp33_ASAP7_75t_R g271 ( .A(n_192), .B(n_21), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_215), .B(n_26), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_209), .A2(n_77), .B(n_31), .C(n_32), .Y(n_273) );
INVx4_ASAP7_75t_L g274 ( .A(n_195), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_231), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g276 ( .A1(n_230), .A2(n_187), .B(n_200), .C(n_190), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_229), .A2(n_200), .B1(n_220), .B2(n_219), .Y(n_277) );
AO32x1_ASAP7_75t_L g278 ( .A1(n_232), .A2(n_28), .A3(n_33), .B1(n_40), .B2(n_44), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_200), .B(n_54), .Y(n_279) );
O2A1O1Ixp33_ASAP7_75t_L g280 ( .A1(n_191), .A2(n_70), .B(n_57), .C(n_59), .Y(n_280) );
O2A1O1Ixp33_ASAP7_75t_L g281 ( .A1(n_223), .A2(n_56), .B(n_62), .C(n_66), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_276), .A2(n_210), .B(n_213), .C(n_212), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
AO31x2_ASAP7_75t_L g284 ( .A1(n_277), .A2(n_224), .A3(n_221), .B(n_198), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_243), .A2(n_221), .B1(n_225), .B2(n_232), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_246), .B(n_232), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_238), .A2(n_245), .B(n_253), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_258), .A2(n_197), .B1(n_198), .B2(n_204), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_252), .A2(n_197), .B(n_204), .C(n_208), .Y(n_289) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_239), .A2(n_208), .B(n_211), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_240), .A2(n_211), .B(n_68), .Y(n_291) );
CKINVDCx11_ASAP7_75t_R g292 ( .A(n_261), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_277), .A2(n_252), .A3(n_269), .B(n_268), .Y(n_293) );
AO32x2_ASAP7_75t_L g294 ( .A1(n_245), .A2(n_274), .A3(n_278), .B1(n_258), .B2(n_248), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_263), .B(n_250), .Y(n_295) );
A2O1A1Ixp33_ASAP7_75t_L g296 ( .A1(n_279), .A2(n_273), .B(n_244), .C(n_275), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_254), .A2(n_279), .B(n_257), .Y(n_297) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_264), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_250), .A2(n_260), .B1(n_251), .B2(n_255), .Y(n_299) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_256), .A2(n_265), .B(n_242), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_241), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_270), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_237), .A2(n_266), .B1(n_247), .B2(n_264), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_264), .Y(n_304) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_237), .A2(n_280), .B(n_272), .C(n_236), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_237), .B(n_249), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_236), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_271), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_259), .Y(n_309) );
NOR2xp67_ASAP7_75t_SL g310 ( .A(n_278), .B(n_281), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_262), .A2(n_240), .B(n_239), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_278), .A2(n_203), .B(n_218), .Y(n_312) );
AO31x2_ASAP7_75t_L g313 ( .A1(n_277), .A2(n_252), .A3(n_269), .B(n_268), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_165), .B(n_238), .C(n_190), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_296), .B(n_314), .C(n_303), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_287), .A2(n_312), .B(n_300), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_283), .B(n_295), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_300), .A2(n_297), .B(n_305), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_302), .A2(n_292), .B1(n_301), .B2(n_306), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_311), .A2(n_289), .B(n_290), .Y(n_320) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_291), .A2(n_290), .B(n_303), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g323 ( .A1(n_308), .A2(n_285), .B1(n_299), .B2(n_288), .C(n_282), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_298), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_286), .A2(n_309), .B(n_288), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_310), .A2(n_298), .B1(n_304), .B2(n_294), .C(n_284), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_304), .A2(n_293), .B(n_313), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_284), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_293), .A2(n_313), .B(n_294), .Y(n_332) );
OA21x2_ASAP7_75t_L g333 ( .A1(n_293), .A2(n_313), .B(n_294), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_287), .A2(n_296), .B(n_312), .Y(n_334) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_314), .A2(n_276), .B(n_277), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_192), .B1(n_249), .B2(n_193), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_307), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_287), .A2(n_296), .B(n_312), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_302), .A2(n_192), .B1(n_165), .B2(n_193), .Y(n_340) );
AO21x2_ASAP7_75t_L g341 ( .A1(n_312), .A2(n_287), .B(n_300), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_287), .A2(n_296), .B(n_312), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_333), .B(n_331), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_322), .Y(n_344) );
AO21x2_ASAP7_75t_L g345 ( .A1(n_316), .A2(n_342), .B(n_339), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_329), .B(n_315), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_331), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g349 ( .A1(n_323), .A2(n_335), .B1(n_317), .B2(n_337), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_337), .Y(n_350) );
OR2x6_ASAP7_75t_L g351 ( .A(n_325), .B(n_338), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_333), .B(n_338), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_341), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_341), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_324), .B(n_330), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_327), .B(n_326), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_333), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_332), .B(n_341), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_324), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_321), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_336), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_318), .A2(n_334), .B(n_320), .Y(n_365) );
AO21x2_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_316), .B(n_334), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_319), .B(n_333), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_324), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_325), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_333), .B(n_331), .Y(n_370) );
AO21x1_ASAP7_75t_SL g371 ( .A1(n_331), .A2(n_335), .B(n_330), .Y(n_371) );
INVx3_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
AO22x1_ASAP7_75t_L g373 ( .A1(n_367), .A2(n_364), .B1(n_363), .B2(n_344), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_343), .B(n_370), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_343), .B(n_370), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_347), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_369), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_369), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_370), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_367), .B(n_363), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_364), .A2(n_349), .B1(n_367), .B2(n_366), .Y(n_385) );
OAI221xp5_ASAP7_75t_SL g386 ( .A1(n_364), .A2(n_349), .B1(n_350), .B2(n_346), .C(n_357), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_352), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_359), .B(n_352), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_357), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_359), .B(n_358), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_358), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_366), .B(n_346), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_351), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_366), .B(n_346), .Y(n_396) );
BUFx2_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
NOR2x1_ASAP7_75t_SL g398 ( .A(n_351), .B(n_371), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_344), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_366), .B(n_345), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_351), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_364), .A2(n_366), .B1(n_350), .B2(n_346), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_345), .B(n_354), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_354), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_345), .B(n_346), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_354), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_345), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_355), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_355), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_348), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_406), .Y(n_411) );
NAND2xp33_ASAP7_75t_R g412 ( .A(n_374), .B(n_372), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_399), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_383), .B(n_345), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_374), .B(n_346), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_399), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_387), .B(n_346), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_399), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_387), .B(n_365), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_383), .B(n_348), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_376), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_376), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_387), .B(n_365), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_377), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_388), .B(n_365), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_374), .B(n_371), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_375), .B(n_371), .Y(n_428) );
NOR2xp67_ASAP7_75t_L g429 ( .A(n_407), .B(n_360), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_375), .B(n_361), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_383), .B(n_360), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_391), .B(n_356), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_388), .B(n_361), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_391), .B(n_356), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_375), .B(n_361), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_407), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_398), .B(n_362), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_388), .B(n_362), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_392), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_391), .B(n_356), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_382), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_380), .B(n_356), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_390), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_380), .B(n_368), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_382), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_389), .B(n_356), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_384), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_389), .B(n_368), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_389), .B(n_368), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_400), .B(n_368), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_400), .B(n_368), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_384), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_408), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_400), .B(n_372), .Y(n_456) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_407), .B(n_372), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_410), .B(n_372), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_443), .B(n_385), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_419), .B(n_402), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_419), .B(n_402), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_419), .B(n_403), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_443), .B(n_385), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_411), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_421), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_421), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_445), .B(n_386), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_429), .B(n_397), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_443), .B(n_403), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_420), .B(n_403), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_423), .B(n_393), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_420), .B(n_422), .Y(n_472) );
XOR2xp5_ASAP7_75t_L g473 ( .A(n_432), .B(n_373), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_429), .B(n_397), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_422), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_424), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_423), .B(n_396), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_424), .B(n_390), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_423), .B(n_425), .Y(n_479) );
INVxp33_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_425), .B(n_393), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_413), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_414), .B(n_405), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_416), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_426), .B(n_373), .Y(n_485) );
NOR2x1_ASAP7_75t_L g486 ( .A(n_457), .B(n_372), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_426), .B(n_407), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_437), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_442), .B(n_404), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_442), .B(n_404), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_425), .B(n_396), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_416), .B(n_418), .Y(n_492) );
NOR2xp67_ASAP7_75t_L g493 ( .A(n_444), .B(n_405), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_446), .B(n_409), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_446), .B(n_409), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_418), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_414), .B(n_405), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_448), .B(n_408), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_438), .B(n_378), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_427), .B(n_398), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_417), .B(n_393), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_417), .B(n_393), .Y(n_502) );
INVx2_ASAP7_75t_SL g503 ( .A(n_438), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_417), .B(n_415), .Y(n_504) );
OAI211xp5_ASAP7_75t_SL g505 ( .A1(n_436), .A2(n_401), .B(n_395), .C(n_394), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_437), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_453), .B(n_379), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_453), .B(n_379), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_415), .B(n_393), .Y(n_509) );
INVx1_ASAP7_75t_SL g510 ( .A(n_500), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_479), .B(n_428), .Y(n_511) );
NOR2x1_ASAP7_75t_L g512 ( .A(n_500), .B(n_457), .Y(n_512) );
NOR2xp67_ASAP7_75t_SL g513 ( .A(n_503), .B(n_412), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_484), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_479), .B(n_427), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_504), .B(n_428), .Y(n_516) );
OR2x6_ASAP7_75t_L g517 ( .A(n_468), .B(n_444), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_473), .A2(n_386), .B1(n_441), .B2(n_434), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_462), .B(n_454), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_476), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_473), .A2(n_434), .B1(n_441), .B2(n_432), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_462), .B(n_454), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_476), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_488), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_467), .A2(n_440), .B1(n_396), .B2(n_452), .C(n_451), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_504), .B(n_456), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_488), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_460), .B(n_433), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_500), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_484), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_509), .B(n_456), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_465), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_460), .B(n_433), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_469), .B(n_433), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_461), .B(n_439), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_466), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_461), .A2(n_451), .B1(n_456), .B2(n_452), .C1(n_447), .C2(n_396), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_459), .B(n_439), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_480), .B(n_463), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_470), .B(n_439), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_475), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_472), .B(n_430), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_483), .B(n_430), .Y(n_545) );
INVx3_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_480), .A2(n_458), .B(n_436), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_483), .B(n_435), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_497), .B(n_435), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_482), .B(n_458), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_478), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_509), .B(n_451), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_517), .A2(n_512), .B(n_525), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_520), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_523), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_541), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_551), .B(n_497), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_524), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_527), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_529), .B(n_492), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_532), .Y(n_562) );
OAI211xp5_ASAP7_75t_L g563 ( .A1(n_525), .A2(n_503), .B(n_493), .C(n_485), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_552), .B(n_487), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_545), .B(n_491), .Y(n_566) );
AND2x2_ASAP7_75t_SL g567 ( .A(n_529), .B(n_438), .Y(n_567) );
AOI211x1_ASAP7_75t_SL g568 ( .A1(n_521), .A2(n_505), .B(n_499), .C(n_498), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_542), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_544), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_529), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_548), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_549), .Y(n_573) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_518), .A2(n_496), .B(n_436), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_510), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_539), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_540), .B(n_481), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g578 ( .A1(n_539), .A2(n_481), .B(n_471), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_538), .B(n_477), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_517), .A2(n_492), .B1(n_468), .B2(n_474), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_554), .A2(n_517), .B1(n_546), .B2(n_530), .Y(n_581) );
OAI222xp33_ASAP7_75t_L g582 ( .A1(n_576), .A2(n_513), .B1(n_530), .B2(n_514), .C1(n_522), .C2(n_519), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_580), .B(n_546), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_574), .A2(n_537), .B1(n_396), .B2(n_550), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_572), .B(n_550), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_564), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_563), .A2(n_471), .B1(n_477), .B2(n_491), .Y(n_587) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_574), .A2(n_514), .B(n_547), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_564), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_558), .B(n_516), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_578), .A2(n_501), .B1(n_502), .B2(n_511), .Y(n_591) );
OAI222xp33_ASAP7_75t_L g592 ( .A1(n_561), .A2(n_575), .B1(n_571), .B2(n_558), .C1(n_573), .C2(n_579), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g593 ( .A1(n_568), .A2(n_546), .B(n_496), .C(n_533), .Y(n_593) );
NAND2x1_ASAP7_75t_SL g594 ( .A(n_562), .B(n_515), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_567), .A2(n_502), .B1(n_501), .B2(n_543), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_565), .A2(n_452), .B1(n_436), .B2(n_438), .Y(n_596) );
OAI211xp5_ASAP7_75t_L g597 ( .A1(n_583), .A2(n_570), .B(n_569), .C(n_579), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g598 ( .A1(n_581), .A2(n_555), .B(n_560), .Y(n_598) );
AOI21xp5_ASAP7_75t_L g599 ( .A1(n_581), .A2(n_556), .B(n_559), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_586), .Y(n_600) );
OAI211xp5_ASAP7_75t_SL g601 ( .A1(n_584), .A2(n_535), .B(n_528), .C(n_577), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_588), .A2(n_557), .B1(n_531), .B2(n_553), .Y(n_602) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_592), .A2(n_468), .B(n_474), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_L g604 ( .A1(n_582), .A2(n_566), .B(n_474), .C(n_534), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_593), .B(n_486), .C(n_541), .Y(n_605) );
NAND5xp2_ASAP7_75t_L g606 ( .A(n_604), .B(n_587), .C(n_595), .D(n_596), .E(n_591), .Y(n_606) );
NAND5xp2_ASAP7_75t_L g607 ( .A(n_605), .B(n_590), .C(n_589), .D(n_585), .E(n_594), .Y(n_607) );
AOI211x1_ASAP7_75t_L g608 ( .A1(n_597), .A2(n_526), .B(n_489), .C(n_490), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_600), .Y(n_609) );
OAI211xp5_ASAP7_75t_SL g610 ( .A1(n_602), .A2(n_603), .B(n_599), .C(n_598), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_609), .Y(n_611) );
NOR4xp25_ASAP7_75t_L g612 ( .A(n_610), .B(n_601), .C(n_440), .D(n_495), .Y(n_612) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_606), .B(n_431), .C(n_450), .Y(n_613) );
INVxp67_ASAP7_75t_L g614 ( .A(n_611), .Y(n_614) );
OR2x6_ASAP7_75t_L g615 ( .A(n_613), .B(n_608), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_615), .A2(n_607), .B1(n_612), .B2(n_431), .Y(n_616) );
OAI22xp5_ASAP7_75t_SL g617 ( .A1(n_614), .A2(n_381), .B1(n_395), .B2(n_401), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_617), .Y(n_618) );
AOI221xp5_ASAP7_75t_SL g619 ( .A1(n_618), .A2(n_616), .B1(n_455), .B2(n_508), .C(n_507), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_619), .A2(n_449), .B1(n_447), .B2(n_455), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_620), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g622 ( .A1(n_621), .A2(n_449), .B1(n_447), .B2(n_381), .Y(n_622) );
endmodule