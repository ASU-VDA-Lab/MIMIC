module fake_jpeg_7229_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_25),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_58),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_61),
.Y(n_81)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_2),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_4),
.Y(n_73)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_71),
.Y(n_103)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_35),
.B1(n_50),
.B2(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_73),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_49),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_34),
.C(n_49),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_52),
.B1(n_48),
.B2(n_34),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_88),
.B(n_75),
.C(n_84),
.Y(n_91)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_87),
.B1(n_89),
.B2(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_5),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_47),
.B(n_8),
.C(n_12),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_97),
.C(n_101),
.Y(n_108)
);

NOR2xp67_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_13),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_106),
.B1(n_101),
.B2(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_108),
.B(n_94),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_112),
.A2(n_104),
.B1(n_81),
.B2(n_67),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_73),
.B(n_102),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_114),
.A2(n_92),
.B1(n_98),
.B2(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_116),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_95),
.B1(n_99),
.B2(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_107),
.C(n_100),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_14),
.B(n_15),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_17),
.B(n_18),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_19),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_23),
.Y(n_124)
);


endmodule