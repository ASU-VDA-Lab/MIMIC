module fake_netlist_1_12508_n_14 (n_3, n_1, n_2, n_0, n_14);
input n_3;
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
NAND2x1_ASAP7_75t_L g4 ( .A(n_3), .B(n_0), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
NAND2xp33_ASAP7_75t_L g6 ( .A(n_2), .B(n_1), .Y(n_6) );
AND2x4_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
HB1xp67_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_8), .B(n_4), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_6), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_10), .B(n_7), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_9), .B(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_13), .B(n_12), .Y(n_14) );
endmodule