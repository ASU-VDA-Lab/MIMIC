module fake_jpeg_26639_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_23),
.B1(n_14),
.B2(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_44),
.B1(n_45),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_24),
.B1(n_23),
.B2(n_13),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_24),
.B1(n_23),
.B2(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_25),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_55),
.Y(n_72)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_45),
.B1(n_63),
.B2(n_58),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_58),
.Y(n_67)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_40),
.B1(n_37),
.B2(n_27),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_30),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_27),
.B1(n_43),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_73),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_38),
.B1(n_43),
.B2(n_27),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_45),
.B1(n_43),
.B2(n_33),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_60),
.B(n_46),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_80),
.B(n_32),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_47),
.C(n_48),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_68),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_34),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_34),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_61),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_61),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_44),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_32),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_80),
.B(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_95),
.B(n_101),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_71),
.B(n_15),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_74),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_34),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_80),
.B1(n_79),
.B2(n_66),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_98),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_123),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_68),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_104),
.A2(n_105),
.B(n_92),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_77),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_115),
.C(n_102),
.Y(n_132)
);

NAND2x1_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_75),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_111),
.B(n_118),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_77),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_66),
.B1(n_65),
.B2(n_73),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_119),
.B1(n_37),
.B2(n_49),
.Y(n_146)
);

OAI21x1_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_73),
.B(n_67),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_67),
.B1(n_80),
.B2(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_96),
.B1(n_89),
.B2(n_102),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_127),
.A2(n_144),
.B(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_133),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_32),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_102),
.B1(n_90),
.B2(n_93),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_141),
.B1(n_143),
.B2(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_15),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_150),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_138),
.A2(n_111),
.B(n_105),
.Y(n_151)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_92),
.B1(n_89),
.B2(n_99),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_92),
.B1(n_100),
.B2(n_99),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_146),
.B1(n_76),
.B2(n_49),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_99),
.B1(n_100),
.B2(n_81),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_107),
.A2(n_64),
.A3(n_44),
.B1(n_70),
.B2(n_33),
.Y(n_144)
);

INVx5_ASAP7_75t_SL g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_148),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_86),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_78),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_86),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_SL g187 ( 
.A(n_151),
.B(n_152),
.C(n_154),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_106),
.B(n_115),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_135),
.B1(n_128),
.B2(n_133),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_120),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_161),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_76),
.B1(n_57),
.B2(n_64),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_164),
.B1(n_168),
.B2(n_171),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_165),
.B1(n_176),
.B2(n_34),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_57),
.B1(n_53),
.B2(n_52),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_52),
.B1(n_53),
.B2(n_97),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_17),
.B1(n_37),
.B2(n_40),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_127),
.A2(n_97),
.B(n_17),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_39),
.B1(n_35),
.B2(n_28),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_6),
.B(n_10),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_6),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_166),
.B(n_140),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_180),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_125),
.B1(n_145),
.B2(n_139),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_179),
.A2(n_183),
.B1(n_193),
.B2(n_194),
.Y(n_202)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_170),
.B(n_126),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_182),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_169),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_143),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_130),
.Y(n_188)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_62),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_168),
.B1(n_175),
.B2(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_54),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_155),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_16),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_16),
.B1(n_13),
.B2(n_19),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_16),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_169),
.B(n_13),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_197),
.B1(n_165),
.B2(n_180),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_214),
.B1(n_39),
.B2(n_21),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_158),
.C(n_161),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_205),
.C(n_217),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_203),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_152),
.C(n_167),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_210),
.B1(n_213),
.B2(n_215),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_173),
.B1(n_172),
.B2(n_163),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_159),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_19),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_159),
.B1(n_35),
.B2(n_39),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_39),
.B1(n_35),
.B2(n_31),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_185),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_191),
.C(n_188),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_202),
.A2(n_183),
.B1(n_187),
.B2(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_219),
.A2(n_223),
.B1(n_209),
.B2(n_214),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_209),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_39),
.B(n_1),
.C(n_2),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_215),
.B(n_213),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_34),
.B1(n_39),
.B2(n_31),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_21),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

OAI22x1_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_9),
.B1(n_11),
.B2(n_10),
.Y(n_226)
);

OAI321xp33_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_218),
.A3(n_206),
.B1(n_200),
.B2(n_3),
.C(n_4),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_19),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_21),
.Y(n_228)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_31),
.C(n_29),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_234),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_8),
.B(n_11),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_204),
.B(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_31),
.C(n_29),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_239),
.B(n_240),
.Y(n_256)
);

AO221x1_ASAP7_75t_L g240 ( 
.A1(n_226),
.A2(n_219),
.B1(n_221),
.B2(n_234),
.C(n_222),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_21),
.B1(n_12),
.B2(n_8),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_245),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_221),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_239),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_12),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_230),
.B1(n_221),
.B2(n_229),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_5),
.B1(n_7),
.B2(n_11),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_229),
.C(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_252),
.C(n_255),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_6),
.B1(n_10),
.B2(n_8),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_29),
.C(n_28),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_29),
.C(n_28),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_28),
.C(n_21),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.C(n_0),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_12),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_238),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_262),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_243),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_6),
.B(n_10),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_266),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_265),
.A2(n_5),
.B1(n_7),
.B2(n_2),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_269),
.C(n_258),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_5),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_275),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_253),
.C(n_259),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.C(n_0),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_5),
.C(n_7),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_272),
.A2(n_260),
.B(n_263),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_279),
.C(n_276),
.Y(n_281)
);

AOI21x1_ASAP7_75t_SL g280 ( 
.A1(n_278),
.A2(n_273),
.B(n_270),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.C(n_0),
.Y(n_282)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_0),
.C(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_2),
.C(n_0),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_284),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_1),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_1),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_287),
.Y(n_288)
);


endmodule