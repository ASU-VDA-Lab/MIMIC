module fake_ariane_1126_n_6109 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_322, n_251, n_506, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_6109);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_506;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_6109;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_5712;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_625;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_4567;
wire n_786;
wire n_5833;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_2382;
wire n_1213;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_5586;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5984;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_619;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3891;
wire n_3372;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_5179;
wire n_2435;
wire n_5680;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_5549;
wire n_1087;
wire n_632;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_2632;
wire n_5557;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_670;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_5773;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_5858;
wire n_5985;
wire n_604;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_688;
wire n_636;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_986;
wire n_1104;
wire n_887;
wire n_2125;
wire n_1156;
wire n_5123;
wire n_4974;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_3931;
wire n_2190;
wire n_1523;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_5889;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5904;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_1044;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_608;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_811;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_642;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_5921;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_4825;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_5679;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_3595;
wire n_2068;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4164;
wire n_4126;
wire n_5030;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_1056;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_5743;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_875;
wire n_6022;
wire n_2828;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_5705;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_5763;
wire n_3633;
wire n_857;
wire n_6061;
wire n_1235;
wire n_4001;
wire n_2584;
wire n_1462;
wire n_5701;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_6013;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_5478;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_2324;
wire n_840;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_2740;
wire n_1991;
wire n_614;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_5844;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_5938;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_4574;
wire n_896;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_774;
wire n_5548;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3895;
wire n_3707;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_3058;
wire n_946;
wire n_757;
wire n_2047;
wire n_5355;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_5915;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_6046;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_1808;
wire n_6091;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_675;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_610;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_645;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_1276;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_1528;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_612;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2685;
wire n_2061;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_4498;
wire n_772;
wire n_1245;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_3429;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_652;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_5981;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_5735;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_5935;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_5488;
wire n_1105;
wire n_5727;
wire n_3599;
wire n_5988;
wire n_5646;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_5832;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_5470;
wire n_1092;
wire n_4374;
wire n_3205;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_982;
wire n_915;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_4977;
wire n_2492;
wire n_3425;
wire n_2939;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_595;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_2264;
wire n_1950;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_5606;
wire n_2310;
wire n_5911;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_918;
wire n_1968;
wire n_5645;
wire n_639;
wire n_5020;
wire n_673;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6107;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_5631;
wire n_3481;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_5608;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_1204;
wire n_2428;
wire n_994;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_607;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_5887;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_684;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_939;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_4761;
wire n_2052;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_5932;
wire n_1299;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_2797;
wire n_5823;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_1069;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_603;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_850;
wire n_4299;
wire n_5625;
wire n_2407;
wire n_690;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_5570;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_5978;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_665;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_672;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_5290;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_5847;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_5718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5546;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_5544;
wire n_5660;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_5610;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_5808;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_5710;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_2220;
wire n_6108;
wire n_6100;
wire n_4433;
wire n_2829;
wire n_5862;
wire n_1914;
wire n_2253;
wire n_5886;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_5630;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_6057;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_3968;
wire n_1365;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_5793;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_627;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3492;
wire n_3044;
wire n_3737;
wire n_5657;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_618;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_643;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_897;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_1659;
wire n_3955;
wire n_885;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_5903;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_5446;
wire n_4561;
wire n_3291;
wire n_597;
wire n_1541;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_3289;
wire n_1955;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_5962;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_613;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_6007;
wire n_621;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_5692;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_5952;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_1077;
wire n_5980;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_5790;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_648;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_654;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_5859;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4609;
wire n_4361;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_723;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1982;
wire n_641;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_954;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_599;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_4014;
wire n_3547;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_782;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_5900;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_5851;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_634;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_5656;
wire n_1988;
wire n_5678;
wire n_5865;
wire n_6050;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_2155;
wire n_615;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_5659;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_598;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_6028;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_5943;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_5857;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2932;
wire n_2027;
wire n_600;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3922;
wire n_3039;
wire n_2195;
wire n_5455;
wire n_1467;
wire n_5209;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_3996;
wire n_3761;
wire n_2031;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_657;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_5972;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_624;
wire n_5577;
wire n_876;
wire n_5872;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_602;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_3694;
wire n_771;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_605;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6039;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_5868;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_5986;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4409;
wire n_4191;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_601;
wire n_628;
wire n_5863;
wire n_3790;
wire n_907;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5774;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_609;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_5925;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_5813;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_5714;
wire n_2169;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_6092;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_5924;
wire n_1845;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_5782;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_596;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_937;
wire n_1631;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_487),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_368),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_288),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_90),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_334),
.Y(n_599)
);

BUFx5_ASAP7_75t_L g600 ( 
.A(n_25),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_456),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_316),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_459),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_404),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_147),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_23),
.Y(n_606)
);

CKINVDCx14_ASAP7_75t_R g607 ( 
.A(n_343),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_81),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_585),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_118),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_328),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_410),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_569),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_229),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_357),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_361),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_428),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_489),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_532),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_80),
.Y(n_620)
);

INVx1_ASAP7_75t_SL g621 ( 
.A(n_133),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_341),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_131),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_497),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_254),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_589),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_222),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_65),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_127),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_175),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_477),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_570),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_392),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_508),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_19),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_137),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_384),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_452),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_565),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_78),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_399),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_131),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_110),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_163),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_453),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_126),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_125),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_433),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_480),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_319),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_227),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_146),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_587),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_477),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_378),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_6),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_500),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_54),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_414),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_476),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_176),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_445),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_86),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_170),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_179),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_380),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_230),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_230),
.Y(n_669)
);

BUFx10_ASAP7_75t_L g670 ( 
.A(n_324),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_57),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_358),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_246),
.Y(n_673)
);

INVxp33_ASAP7_75t_L g674 ( 
.A(n_263),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_510),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_539),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_102),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_160),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_311),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_367),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_370),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_356),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_472),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_150),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_475),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_490),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_47),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_385),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_285),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_360),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_408),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_80),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_269),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_329),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_299),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_470),
.Y(n_696)
);

CKINVDCx14_ASAP7_75t_R g697 ( 
.A(n_237),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_454),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_14),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_125),
.Y(n_700)
);

BUFx10_ASAP7_75t_L g701 ( 
.A(n_491),
.Y(n_701)
);

BUFx10_ASAP7_75t_L g702 ( 
.A(n_21),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_306),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_172),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_418),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_507),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_436),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_272),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_344),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_400),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_35),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_343),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_498),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_203),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_272),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_474),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_219),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_425),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_126),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_437),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_392),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_492),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_524),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_35),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_312),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_424),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_123),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_493),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_519),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_386),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_387),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_529),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_247),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_304),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_239),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_525),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_14),
.Y(n_737)
);

BUFx5_ASAP7_75t_L g738 ( 
.A(n_518),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_246),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_393),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_577),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_561),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_576),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_451),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_464),
.Y(n_745)
);

CKINVDCx14_ASAP7_75t_R g746 ( 
.A(n_404),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_360),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_283),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_113),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_344),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_308),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_453),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_460),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_201),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_320),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_232),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_132),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_155),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_515),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_348),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_209),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_167),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_581),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_455),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_409),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_484),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_6),
.Y(n_767)
);

BUFx5_ASAP7_75t_L g768 ( 
.A(n_522),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_135),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_319),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_301),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_248),
.Y(n_772)
);

BUFx8_ASAP7_75t_SL g773 ( 
.A(n_72),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_314),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_447),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_419),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_64),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_288),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_435),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_489),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_591),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_250),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_221),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_491),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_511),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_385),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_395),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_27),
.Y(n_788)
);

CKINVDCx20_ASAP7_75t_R g789 ( 
.A(n_262),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_25),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_496),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_201),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_593),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_16),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_95),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_169),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_358),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_145),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_427),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_442),
.Y(n_800)
);

INVx1_ASAP7_75t_SL g801 ( 
.A(n_53),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_434),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_17),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_48),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_171),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_380),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_253),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_420),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_487),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_419),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_37),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_407),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_458),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_18),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_560),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_506),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_528),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_405),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_53),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_92),
.Y(n_820)
);

INVx1_ASAP7_75t_SL g821 ( 
.A(n_554),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_73),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_432),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_457),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_428),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_539),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_328),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_144),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_64),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_237),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_422),
.Y(n_831)
);

BUFx5_ASAP7_75t_L g832 ( 
.A(n_519),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_347),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_335),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_45),
.Y(n_835)
);

CKINVDCx16_ASAP7_75t_R g836 ( 
.A(n_42),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_350),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_366),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_522),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_194),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_381),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_327),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_97),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_120),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_171),
.Y(n_845)
);

CKINVDCx14_ASAP7_75t_R g846 ( 
.A(n_383),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_10),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_259),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_336),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_367),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_463),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_104),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_238),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_254),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_531),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_372),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_342),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_362),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_115),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_441),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_484),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_421),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_543),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_102),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_167),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_488),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_194),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_411),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_190),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_359),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_156),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_115),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_215),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_439),
.Y(n_874)
);

BUFx5_ASAP7_75t_L g875 ( 
.A(n_546),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_264),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_334),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_188),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_273),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_306),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_530),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_77),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_527),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_513),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_216),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_322),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_104),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_100),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_45),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_399),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_119),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_238),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_521),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_350),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_242),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_279),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_185),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_83),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_431),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_43),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_277),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_155),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_594),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_108),
.Y(n_904)
);

BUFx5_ASAP7_75t_L g905 ( 
.A(n_70),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_542),
.Y(n_906)
);

CKINVDCx14_ASAP7_75t_R g907 ( 
.A(n_365),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_26),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_242),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_100),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_245),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_427),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_175),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_450),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_431),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_181),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_346),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_509),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_172),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_530),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_19),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_299),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_65),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_231),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_512),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_78),
.Y(n_926)
);

BUFx10_ASAP7_75t_L g927 ( 
.A(n_579),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_270),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_315),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_443),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_377),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_499),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_87),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_202),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_566),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_182),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_555),
.Y(n_937)
);

BUFx2_ASAP7_75t_L g938 ( 
.A(n_454),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_475),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_217),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_398),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_526),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_29),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_227),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_289),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_40),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_515),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_203),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_204),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_543),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_473),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_412),
.Y(n_952)
);

BUFx8_ASAP7_75t_SL g953 ( 
.A(n_216),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_553),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_403),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_386),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_405),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_336),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_516),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_121),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_408),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_31),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_28),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_363),
.Y(n_964)
);

BUFx10_ASAP7_75t_L g965 ( 
.A(n_218),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_410),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_48),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_463),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_320),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_110),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_307),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_0),
.Y(n_972)
);

CKINVDCx16_ASAP7_75t_R g973 ( 
.A(n_574),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_406),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_137),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_327),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_42),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_311),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_82),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_483),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_424),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_403),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_495),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_136),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_429),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_468),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_50),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_582),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_345),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_314),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_389),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_448),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_390),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_187),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_547),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_535),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_553),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_573),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_270),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_277),
.Y(n_1000)
);

CKINVDCx20_ASAP7_75t_R g1001 ( 
.A(n_473),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_369),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_586),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_146),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_178),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_377),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_538),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_234),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_141),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_302),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_537),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_293),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_129),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_333),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_212),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_106),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_401),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_560),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_469),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_490),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_391),
.Y(n_1021)
);

INVxp33_ASAP7_75t_L g1022 ( 
.A(n_286),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_524),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_393),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_400),
.Y(n_1025)
);

CKINVDCx16_ASAP7_75t_R g1026 ( 
.A(n_373),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_240),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_375),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_378),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_388),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_351),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_429),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_422),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_345),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_359),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_355),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_544),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_113),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_73),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_411),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_470),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_302),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_442),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_267),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_412),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_223),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_517),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_2),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_523),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_274),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_449),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_41),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_467),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_494),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_205),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_186),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_109),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_371),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_296),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_588),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_547),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_23),
.Y(n_1062)
);

CKINVDCx20_ASAP7_75t_R g1063 ( 
.A(n_364),
.Y(n_1063)
);

BUFx5_ASAP7_75t_L g1064 ( 
.A(n_262),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_471),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_55),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_538),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_518),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_513),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_458),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_251),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_459),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_220),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_291),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_281),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_558),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_116),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_402),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_364),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_558),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_536),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_245),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_9),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_34),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_91),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_269),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_374),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_520),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_43),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_105),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_580),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_28),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_471),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_12),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_260),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_517),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_382),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_47),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_50),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_235),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_435),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_413),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_169),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_217),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_81),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_532),
.Y(n_1106)
);

CKINVDCx16_ASAP7_75t_R g1107 ( 
.A(n_373),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_501),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_341),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_527),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_239),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_361),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_409),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_214),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_526),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_292),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_476),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_74),
.Y(n_1118)
);

CKINVDCx20_ASAP7_75t_R g1119 ( 
.A(n_280),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_291),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_263),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_40),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_351),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_551),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_124),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_315),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_788),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_788),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_607),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1064),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_697),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_788),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_746),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_788),
.Y(n_1134)
);

BUFx2_ASAP7_75t_SL g1135 ( 
.A(n_927),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_846),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1064),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_907),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_850),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_973),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_850),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_850),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_973),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_773),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_953),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_741),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_850),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1123),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1123),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_741),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_927),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1123),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_639),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_639),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_1064),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_927),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_639),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1064),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_781),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_728),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_728),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_927),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_747),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_724),
.B(n_0),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_747),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_728),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_776),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_787),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_776),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_836),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_595),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_787),
.Y(n_1172)
);

BUFx10_ASAP7_75t_L g1173 ( 
.A(n_612),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_836),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_612),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_787),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_868),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_830),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_868),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_830),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_877),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_877),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1026),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1026),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_830),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1082),
.Y(n_1186)
);

CKINVDCx16_ASAP7_75t_R g1187 ( 
.A(n_1082),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1107),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1107),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_918),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1116),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_918),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_596),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1124),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1125),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1064),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_918),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_781),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1056),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_1056),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_1056),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1093),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1122),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_724),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1126),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1064),
.Y(n_1206)
);

NOR2xp67_ASAP7_75t_L g1207 ( 
.A(n_666),
.B(n_1),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_599),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_614),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_603),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1064),
.Y(n_1211)
);

CKINVDCx16_ASAP7_75t_R g1212 ( 
.A(n_627),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1064),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1093),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1109),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1109),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1109),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_598),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_604),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_606),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_608),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_666),
.B(n_2),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_640),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1064),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_598),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_598),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_610),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_781),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_700),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_613),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1064),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_600),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_613),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_617),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_610),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_622),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_623),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_817),
.B(n_861),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_610),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_624),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_684),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_684),
.Y(n_1242)
);

NOR2xp67_ASAP7_75t_L g1243 ( 
.A(n_682),
.B(n_3),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_684),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_720),
.Y(n_1245)
);

BUFx2_ASAP7_75t_SL g1246 ( 
.A(n_903),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_699),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_612),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_699),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_699),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_725),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_625),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_725),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_629),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_725),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_631),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_636),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_600),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_642),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_643),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_612),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_729),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_729),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_729),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_739),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_600),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_644),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_739),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_647),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_682),
.B(n_3),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_721),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_739),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_793),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_750),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_627),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_600),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_648),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_650),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_651),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_653),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_655),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_722),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_750),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_627),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_656),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_791),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_791),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_736),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_791),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_817),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_657),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_660),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_661),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_670),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_861),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_662),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_834),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_834),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_663),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_834),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_866),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_866),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_866),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_664),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_886),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_665),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_886),
.Y(n_1307)
);

CKINVDCx16_ASAP7_75t_R g1308 ( 
.A(n_670),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_938),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_886),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_612),
.Y(n_1311)
);

BUFx5_ASAP7_75t_L g1312 ( 
.A(n_793),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_913),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_938),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_913),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_789),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_913),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_794),
.Y(n_1318)
);

CKINVDCx16_ASAP7_75t_R g1319 ( 
.A(n_670),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_928),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_928),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_667),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_668),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_669),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_799),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_928),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_932),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_677),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_678),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_932),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_932),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_970),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_679),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_970),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_942),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_970),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_681),
.Y(n_1337)
);

INVx2_ASAP7_75t_SL g1338 ( 
.A(n_670),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1014),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_600),
.Y(n_1340)
);

CKINVDCx16_ASAP7_75t_R g1341 ( 
.A(n_701),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_600),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1014),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_SL g1344 ( 
.A(n_903),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_683),
.Y(n_1345)
);

CKINVDCx20_ASAP7_75t_R g1346 ( 
.A(n_812),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1014),
.Y(n_1347)
);

CKINVDCx20_ASAP7_75t_R g1348 ( 
.A(n_859),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1021),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_667),
.Y(n_1350)
);

CKINVDCx16_ASAP7_75t_R g1351 ( 
.A(n_701),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_685),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1021),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_686),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_600),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1021),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_687),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_942),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1040),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_600),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_691),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1040),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_692),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1040),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_667),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_694),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_865),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1081),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1114),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1114),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1114),
.Y(n_1371)
);

BUFx5_ASAP7_75t_L g1372 ( 
.A(n_597),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1081),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_738),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_874),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_904),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_695),
.Y(n_1377)
);

CKINVDCx20_ASAP7_75t_R g1378 ( 
.A(n_934),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1121),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1121),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_597),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_696),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_698),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_601),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_703),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_601),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_602),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_955),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_738),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_602),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_605),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_605),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_611),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_611),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_706),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_738),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_708),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_738),
.Y(n_1398)
);

CKINVDCx16_ASAP7_75t_R g1399 ( 
.A(n_701),
.Y(n_1399)
);

INVx2_ASAP7_75t_SL g1400 ( 
.A(n_701),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_710),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_738),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_615),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_738),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1097),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_738),
.B(n_4),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_667),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_712),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_713),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_615),
.B(n_4),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_968),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_715),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_716),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_717),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_738),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_718),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_616),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_719),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_616),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_726),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_727),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_975),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1001),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1010),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1032),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_730),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1046),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_731),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1058),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_618),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_768),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_768),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_618),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_768),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_733),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1027),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_619),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_734),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_619),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_737),
.Y(n_1440)
);

CKINVDCx16_ASAP7_75t_R g1441 ( 
.A(n_702),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_620),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_740),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_620),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_768),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_744),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_676),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_628),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_628),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_632),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_632),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_634),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_634),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_768),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_768),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_745),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1063),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1070),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_748),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_635),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_749),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_635),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_637),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1027),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_637),
.B(n_5),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_638),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_751),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_752),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_638),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_641),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_641),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_753),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_757),
.Y(n_1473)
);

BUFx2_ASAP7_75t_SL g1474 ( 
.A(n_768),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_760),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_645),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_761),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_762),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_711),
.B(n_5),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_645),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_764),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_646),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_646),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1071),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_767),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_770),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_652),
.Y(n_1487)
);

CKINVDCx16_ASAP7_75t_R g1488 ( 
.A(n_702),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_1073),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_771),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_711),
.B(n_7),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_652),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_768),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_658),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_777),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_780),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_783),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_784),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_658),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_659),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_785),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1087),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_1098),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_786),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_659),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_671),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1110),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1119),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_790),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_676),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_671),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_676),
.Y(n_1512)
);

CKINVDCx16_ASAP7_75t_R g1513 ( 
.A(n_702),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_621),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_795),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_796),
.Y(n_1516)
);

CKINVDCx20_ASAP7_75t_R g1517 ( 
.A(n_702),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_672),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_797),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_798),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_672),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_965),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_800),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_802),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_673),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_768),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_965),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_673),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_803),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_675),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_804),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_965),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_805),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_965),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_807),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_649),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_808),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_675),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_680),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_680),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_832),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_813),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_832),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_814),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_816),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_832),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_818),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_819),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_824),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_688),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_688),
.Y(n_1551)
);

BUFx2_ASAP7_75t_L g1552 ( 
.A(n_835),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_690),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_690),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_704),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_649),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_704),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_837),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_705),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_705),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_839),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_707),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_841),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_707),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_709),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_832),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_843),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_709),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_847),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_732),
.Y(n_1570)
);

INVxp67_ASAP7_75t_SL g1571 ( 
.A(n_1159),
.Y(n_1571)
);

INVxp33_ASAP7_75t_L g1572 ( 
.A(n_1290),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1171),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1203),
.Y(n_1574)
);

INVxp67_ASAP7_75t_L g1575 ( 
.A(n_1514),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1135),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1127),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1128),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1132),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1134),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1187),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1139),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1209),
.Y(n_1583)
);

CKINVDCx16_ASAP7_75t_R g1584 ( 
.A(n_1212),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1159),
.Y(n_1585)
);

BUFx2_ASAP7_75t_L g1586 ( 
.A(n_1163),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1144),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1144),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1223),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1145),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1141),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1198),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1142),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1147),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1148),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1149),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1140),
.Y(n_1597)
);

CKINVDCx16_ASAP7_75t_R g1598 ( 
.A(n_1275),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1152),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1153),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1154),
.Y(n_1601)
);

INVxp33_ASAP7_75t_L g1602 ( 
.A(n_1314),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1140),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1175),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1160),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1198),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1161),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1166),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1193),
.Y(n_1609)
);

BUFx2_ASAP7_75t_L g1610 ( 
.A(n_1163),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1435),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1168),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1172),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1176),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1229),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1178),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1175),
.Y(n_1617)
);

INVxp33_ASAP7_75t_SL g1618 ( 
.A(n_1143),
.Y(n_1618)
);

INVxp67_ASAP7_75t_SL g1619 ( 
.A(n_1228),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1143),
.Y(n_1620)
);

BUFx2_ASAP7_75t_SL g1621 ( 
.A(n_1517),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1180),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1252),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1175),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_1254),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_1256),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1185),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1190),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1192),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1173),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1197),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1199),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1202),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1257),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1214),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1215),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1175),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1216),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1217),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1407),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1259),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1260),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1245),
.Y(n_1643)
);

CKINVDCx20_ASAP7_75t_R g1644 ( 
.A(n_1271),
.Y(n_1644)
);

INVxp33_ASAP7_75t_SL g1645 ( 
.A(n_1129),
.Y(n_1645)
);

CKINVDCx14_ASAP7_75t_R g1646 ( 
.A(n_1129),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1447),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1379),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1288),
.Y(n_1649)
);

INVxp33_ASAP7_75t_SL g1650 ( 
.A(n_1131),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1380),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_1316),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1381),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1384),
.Y(n_1654)
);

CKINVDCx20_ASAP7_75t_R g1655 ( 
.A(n_1318),
.Y(n_1655)
);

INVxp67_ASAP7_75t_SL g1656 ( 
.A(n_1436),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1386),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1387),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1145),
.Y(n_1659)
);

INVxp33_ASAP7_75t_L g1660 ( 
.A(n_1335),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_1464),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1165),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1390),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1391),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1392),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1393),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1394),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1403),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1417),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1346),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1419),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1282),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1430),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1165),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1433),
.Y(n_1675)
);

CKINVDCx20_ASAP7_75t_R g1676 ( 
.A(n_1348),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1437),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1175),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1261),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1267),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1439),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1442),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1367),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1444),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1448),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1449),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1325),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1167),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1450),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1451),
.Y(n_1690)
);

CKINVDCx16_ASAP7_75t_R g1691 ( 
.A(n_1294),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1167),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1452),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1261),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1453),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1460),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1462),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1463),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1466),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1429),
.Y(n_1700)
);

HB1xp67_ASAP7_75t_L g1701 ( 
.A(n_1169),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1469),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1470),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1471),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1476),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1261),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1480),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1484),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1261),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1489),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1482),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1483),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1487),
.Y(n_1713)
);

CKINVDCx16_ASAP7_75t_R g1714 ( 
.A(n_1308),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1375),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1376),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1378),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1492),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1299),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1494),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1499),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1261),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1500),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1505),
.Y(n_1724)
);

CKINVDCx14_ASAP7_75t_R g1725 ( 
.A(n_1131),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1133),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1304),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1306),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1311),
.Y(n_1729)
);

CKINVDCx16_ASAP7_75t_R g1730 ( 
.A(n_1319),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1506),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1511),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1518),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1521),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1525),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1438),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1528),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1530),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1538),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1323),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1539),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1540),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1324),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1311),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_SL g1745 ( 
.A(n_1284),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1328),
.Y(n_1746)
);

CKINVDCx14_ASAP7_75t_R g1747 ( 
.A(n_1133),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1329),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1550),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1551),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_1388),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1553),
.Y(n_1752)
);

INVxp33_ASAP7_75t_L g1753 ( 
.A(n_1524),
.Y(n_1753)
);

CKINVDCx20_ASAP7_75t_R g1754 ( 
.A(n_1411),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1333),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1554),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1552),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1555),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1337),
.Y(n_1759)
);

CKINVDCx16_ASAP7_75t_R g1760 ( 
.A(n_1341),
.Y(n_1760)
);

CKINVDCx16_ASAP7_75t_R g1761 ( 
.A(n_1351),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1311),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1557),
.Y(n_1763)
);

CKINVDCx16_ASAP7_75t_R g1764 ( 
.A(n_1399),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1559),
.Y(n_1765)
);

INVxp67_ASAP7_75t_L g1766 ( 
.A(n_1536),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1560),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1345),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1422),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1169),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1352),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1170),
.Y(n_1772)
);

INVxp67_ASAP7_75t_SL g1773 ( 
.A(n_1404),
.Y(n_1773)
);

CKINVDCx16_ASAP7_75t_R g1774 ( 
.A(n_1441),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1556),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1170),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1311),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1562),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1564),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1311),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1565),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1354),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1568),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1570),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1357),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1361),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_1423),
.Y(n_1787)
);

INVxp33_ASAP7_75t_SL g1788 ( 
.A(n_1136),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1157),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1151),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1157),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1200),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1424),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1200),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1201),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1151),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1156),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1201),
.Y(n_1798)
);

CKINVDCx20_ASAP7_75t_R g1799 ( 
.A(n_1425),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1406),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1218),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1225),
.Y(n_1802)
);

INVxp33_ASAP7_75t_SL g1803 ( 
.A(n_1136),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1156),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1226),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1227),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1427),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1235),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1246),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1239),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1241),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1242),
.Y(n_1812)
);

INVxp33_ASAP7_75t_SL g1813 ( 
.A(n_1138),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1457),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1244),
.Y(n_1815)
);

INVxp33_ASAP7_75t_SL g1816 ( 
.A(n_1138),
.Y(n_1816)
);

CKINVDCx20_ASAP7_75t_R g1817 ( 
.A(n_1458),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1247),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1204),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1249),
.Y(n_1820)
);

INVxp67_ASAP7_75t_SL g1821 ( 
.A(n_1415),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1250),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1502),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1174),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1251),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1522),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1253),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1322),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1255),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_1503),
.Y(n_1830)
);

INVxp67_ASAP7_75t_SL g1831 ( 
.A(n_1431),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1295),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1162),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1262),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1322),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1263),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1264),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1162),
.Y(n_1838)
);

CKINVDCx16_ASAP7_75t_R g1839 ( 
.A(n_1488),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1265),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1268),
.Y(n_1841)
);

BUFx6f_ASAP7_75t_L g1842 ( 
.A(n_1322),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1507),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1272),
.Y(n_1844)
);

BUFx3_ASAP7_75t_L g1845 ( 
.A(n_1431),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1274),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1527),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1191),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1283),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1191),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1286),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1194),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1287),
.Y(n_1853)
);

BUFx5_ASAP7_75t_L g1854 ( 
.A(n_1546),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1289),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1297),
.Y(n_1856)
);

CKINVDCx16_ASAP7_75t_R g1857 ( 
.A(n_1513),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1298),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1300),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1301),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1173),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1194),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1322),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1195),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1195),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_1508),
.Y(n_1866)
);

CKINVDCx20_ASAP7_75t_R g1867 ( 
.A(n_1532),
.Y(n_1867)
);

INVxp33_ASAP7_75t_L g1868 ( 
.A(n_1238),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1205),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1205),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1302),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1303),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1305),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1230),
.Y(n_1874)
);

INVxp33_ASAP7_75t_L g1875 ( 
.A(n_1309),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1307),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1208),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1177),
.Y(n_1878)
);

CKINVDCx20_ASAP7_75t_R g1879 ( 
.A(n_1534),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1310),
.Y(n_1880)
);

INVxp67_ASAP7_75t_SL g1881 ( 
.A(n_1230),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1313),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1179),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1233),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1173),
.Y(n_1885)
);

CKINVDCx20_ASAP7_75t_R g1886 ( 
.A(n_1179),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1315),
.Y(n_1887)
);

INVxp33_ASAP7_75t_SL g1888 ( 
.A(n_1210),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1317),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1322),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1320),
.Y(n_1891)
);

CKINVDCx20_ASAP7_75t_R g1892 ( 
.A(n_1181),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_1210),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1321),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1326),
.Y(n_1895)
);

BUFx2_ASAP7_75t_SL g1896 ( 
.A(n_1284),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1219),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1327),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1330),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1331),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1248),
.Y(n_1901)
);

CKINVDCx20_ASAP7_75t_R g1902 ( 
.A(n_1181),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1332),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1334),
.Y(n_1904)
);

HB1xp67_ASAP7_75t_L g1905 ( 
.A(n_1182),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1248),
.Y(n_1906)
);

CKINVDCx14_ASAP7_75t_R g1907 ( 
.A(n_1182),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1219),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1350),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1336),
.Y(n_1910)
);

CKINVDCx20_ASAP7_75t_R g1911 ( 
.A(n_1183),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1350),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1339),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1343),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1220),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1347),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1358),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1220),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1349),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1353),
.Y(n_1920)
);

CKINVDCx20_ASAP7_75t_R g1921 ( 
.A(n_1183),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1356),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1221),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1184),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1184),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1359),
.Y(n_1926)
);

HB1xp67_ASAP7_75t_L g1927 ( 
.A(n_1186),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_1186),
.Y(n_1928)
);

CKINVDCx16_ASAP7_75t_R g1929 ( 
.A(n_1344),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1577),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1604),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1604),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1578),
.Y(n_1933)
);

CKINVDCx6p67_ASAP7_75t_R g1934 ( 
.A(n_1584),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1575),
.Y(n_1935)
);

OAI21x1_ASAP7_75t_L g1936 ( 
.A1(n_1800),
.A2(n_1258),
.B(n_1232),
.Y(n_1936)
);

BUFx8_ASAP7_75t_SL g1937 ( 
.A(n_1573),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1819),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1790),
.A2(n_1150),
.B1(n_1146),
.B2(n_1164),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1845),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1617),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1874),
.B(n_1233),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1617),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1881),
.B(n_1338),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1845),
.Y(n_1945)
);

BUFx3_ASAP7_75t_L g1946 ( 
.A(n_1854),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1579),
.Y(n_1947)
);

CKINVDCx6p67_ASAP7_75t_R g1948 ( 
.A(n_1598),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1624),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_SL g1950 ( 
.A1(n_1867),
.A2(n_1150),
.B1(n_1146),
.B2(n_1188),
.Y(n_1950)
);

BUFx8_ASAP7_75t_SL g1951 ( 
.A(n_1573),
.Y(n_1951)
);

AND2x6_ASAP7_75t_L g1952 ( 
.A(n_1580),
.B(n_1273),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1623),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1582),
.Y(n_1954)
);

AND2x6_ASAP7_75t_L g1955 ( 
.A(n_1591),
.B(n_1273),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1884),
.B(n_1338),
.Y(n_1956)
);

BUFx8_ASAP7_75t_L g1957 ( 
.A(n_1586),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1896),
.A2(n_829),
.B1(n_1022),
.B2(n_674),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1624),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1637),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1679),
.Y(n_1961)
);

BUFx8_ASAP7_75t_L g1962 ( 
.A(n_1610),
.Y(n_1962)
);

BUFx6f_ASAP7_75t_L g1963 ( 
.A(n_1679),
.Y(n_1963)
);

BUFx12f_ASAP7_75t_L g1964 ( 
.A(n_1587),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1609),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_SL g1966 ( 
.A(n_1929),
.B(n_1188),
.Y(n_1966)
);

OAI21x1_ASAP7_75t_L g1967 ( 
.A1(n_1637),
.A2(n_1258),
.B(n_1232),
.Y(n_1967)
);

AND2x4_ASAP7_75t_L g1968 ( 
.A(n_1571),
.B(n_1400),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1640),
.B(n_1585),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1593),
.B(n_1400),
.Y(n_1970)
);

BUFx8_ASAP7_75t_L g1971 ( 
.A(n_1674),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1594),
.Y(n_1972)
);

BUFx6f_ASAP7_75t_L g1973 ( 
.A(n_1679),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1678),
.Y(n_1974)
);

OAI22x1_ASAP7_75t_SL g1975 ( 
.A1(n_1867),
.A2(n_1189),
.B1(n_1234),
.B2(n_1221),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1842),
.Y(n_1976)
);

BUFx2_ASAP7_75t_L g1977 ( 
.A(n_1832),
.Y(n_1977)
);

INVx6_ASAP7_75t_L g1978 ( 
.A(n_1861),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1581),
.Y(n_1979)
);

BUFx8_ASAP7_75t_L g1980 ( 
.A(n_1692),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1678),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1592),
.B(n_1474),
.Y(n_1982)
);

INVx3_ASAP7_75t_L g1983 ( 
.A(n_1842),
.Y(n_1983)
);

INVx2_ASAP7_75t_SL g1984 ( 
.A(n_1719),
.Y(n_1984)
);

NOR2x1_ASAP7_75t_L g1985 ( 
.A(n_1789),
.B(n_1207),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1801),
.Y(n_1986)
);

BUFx12f_ASAP7_75t_L g1987 ( 
.A(n_1588),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1606),
.B(n_1312),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1694),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1802),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1805),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1806),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1706),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1706),
.A2(n_1276),
.B(n_1266),
.Y(n_1994)
);

OAI21x1_ASAP7_75t_L g1995 ( 
.A1(n_1709),
.A2(n_1276),
.B(n_1266),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1727),
.Y(n_1996)
);

BUFx6f_ASAP7_75t_L g1997 ( 
.A(n_1842),
.Y(n_1997)
);

HB1xp67_ASAP7_75t_L g1998 ( 
.A(n_1917),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1842),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1868),
.B(n_1362),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1709),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_L g2002 ( 
.A(n_1722),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1611),
.Y(n_2003)
);

OAI22x1_ASAP7_75t_R g2004 ( 
.A1(n_1883),
.A2(n_1189),
.B1(n_1236),
.B2(n_1234),
.Y(n_2004)
);

INVx2_ASAP7_75t_SL g2005 ( 
.A(n_1623),
.Y(n_2005)
);

BUFx12f_ASAP7_75t_L g2006 ( 
.A(n_1590),
.Y(n_2006)
);

BUFx6f_ASAP7_75t_L g2007 ( 
.A(n_1729),
.Y(n_2007)
);

BUFx12f_ASAP7_75t_L g2008 ( 
.A(n_1659),
.Y(n_2008)
);

OAI21x1_ASAP7_75t_L g2009 ( 
.A1(n_1744),
.A2(n_1342),
.B(n_1340),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1625),
.Y(n_2010)
);

BUFx12f_ASAP7_75t_L g2011 ( 
.A(n_1625),
.Y(n_2011)
);

BUFx12f_ASAP7_75t_L g2012 ( 
.A(n_1626),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1772),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1808),
.Y(n_2014)
);

BUFx8_ASAP7_75t_SL g2015 ( 
.A(n_1574),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1810),
.Y(n_2016)
);

CKINVDCx6p67_ASAP7_75t_R g2017 ( 
.A(n_1691),
.Y(n_2017)
);

OA21x2_ASAP7_75t_L g2018 ( 
.A1(n_1762),
.A2(n_1342),
.B(n_1340),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1811),
.Y(n_2019)
);

BUFx8_ASAP7_75t_SL g2020 ( 
.A(n_1574),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1648),
.B(n_1364),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1812),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1777),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1576),
.B(n_1236),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1777),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1815),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1619),
.B(n_1312),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1818),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1809),
.B(n_1237),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1780),
.Y(n_2030)
);

INVx5_ASAP7_75t_L g2031 ( 
.A(n_1630),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1736),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1790),
.A2(n_1243),
.B1(n_1270),
.B2(n_1222),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1651),
.B(n_1653),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1780),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1647),
.B(n_1312),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1654),
.B(n_1369),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1828),
.Y(n_2038)
);

OA21x2_ASAP7_75t_L g2039 ( 
.A1(n_1828),
.A2(n_1360),
.B(n_1355),
.Y(n_2039)
);

INVx3_ASAP7_75t_L g2040 ( 
.A(n_1835),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1835),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1630),
.B(n_1656),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1791),
.B(n_1373),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1863),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1630),
.Y(n_2045)
);

BUFx6f_ASAP7_75t_L g2046 ( 
.A(n_1863),
.Y(n_2046)
);

AND2x4_ASAP7_75t_L g2047 ( 
.A(n_1792),
.B(n_1410),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1890),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1820),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1890),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1657),
.B(n_1370),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1909),
.Y(n_2052)
);

INVx3_ASAP7_75t_L g2053 ( 
.A(n_1909),
.Y(n_2053)
);

AND2x6_ASAP7_75t_L g2054 ( 
.A(n_1595),
.B(n_732),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1912),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1912),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1822),
.Y(n_2057)
);

BUFx12f_ASAP7_75t_L g2058 ( 
.A(n_1626),
.Y(n_2058)
);

INVx3_ASAP7_75t_L g2059 ( 
.A(n_1854),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1885),
.Y(n_2060)
);

NOR2x1_ASAP7_75t_L g2061 ( 
.A(n_1794),
.B(n_1479),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_1757),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1596),
.A2(n_1360),
.B(n_1355),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1825),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1827),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1661),
.B(n_1312),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1829),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1834),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1796),
.B(n_1237),
.Y(n_2069)
);

BUFx6f_ASAP7_75t_L g2070 ( 
.A(n_1836),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1837),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1658),
.B(n_1371),
.Y(n_2072)
);

AND2x6_ASAP7_75t_L g2073 ( 
.A(n_1599),
.B(n_735),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1840),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1663),
.B(n_1240),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1634),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1841),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1844),
.Y(n_2078)
);

AOI22xp5_ASAP7_75t_L g2079 ( 
.A1(n_1796),
.A2(n_1491),
.B1(n_621),
.B2(n_689),
.Y(n_2079)
);

OAI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1797),
.A2(n_1368),
.B1(n_919),
.B2(n_1054),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1846),
.Y(n_2081)
);

AND2x4_ASAP7_75t_L g2082 ( 
.A(n_1795),
.B(n_1465),
.Y(n_2082)
);

BUFx6f_ASAP7_75t_L g2083 ( 
.A(n_1849),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_1851),
.Y(n_2084)
);

BUFx12f_ASAP7_75t_L g2085 ( 
.A(n_1634),
.Y(n_2085)
);

OAI22x1_ASAP7_75t_R g2086 ( 
.A1(n_1883),
.A2(n_1892),
.B1(n_1902),
.B2(n_1886),
.Y(n_2086)
);

INVx3_ASAP7_75t_L g2087 ( 
.A(n_1901),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_1745),
.B(n_1240),
.Y(n_2088)
);

INVxp67_ASAP7_75t_L g2089 ( 
.A(n_1672),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1853),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1797),
.A2(n_689),
.B1(n_723),
.B2(n_630),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1855),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_1798),
.B(n_792),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_1687),
.Y(n_2094)
);

OAI22x1_ASAP7_75t_L g2095 ( 
.A1(n_1766),
.A2(n_1405),
.B1(n_723),
.B2(n_778),
.Y(n_2095)
);

BUFx6f_ASAP7_75t_L g2096 ( 
.A(n_1856),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_1901),
.Y(n_2097)
);

BUFx3_ASAP7_75t_L g2098 ( 
.A(n_1906),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1858),
.Y(n_2099)
);

CKINVDCx5p33_ASAP7_75t_R g2100 ( 
.A(n_1641),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1600),
.B(n_792),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1859),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1860),
.Y(n_2103)
);

CKINVDCx16_ASAP7_75t_R g2104 ( 
.A(n_1714),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1871),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_SL g2106 ( 
.A1(n_1879),
.A2(n_778),
.B1(n_801),
.B2(n_630),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1804),
.A2(n_714),
.B1(n_1054),
.B2(n_919),
.Y(n_2107)
);

BUFx6f_ASAP7_75t_L g2108 ( 
.A(n_1872),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1873),
.Y(n_2109)
);

BUFx6f_ASAP7_75t_L g2110 ( 
.A(n_1876),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1880),
.Y(n_2111)
);

BUFx6f_ASAP7_75t_L g2112 ( 
.A(n_1882),
.Y(n_2112)
);

OA21x2_ASAP7_75t_L g2113 ( 
.A1(n_1887),
.A2(n_1389),
.B(n_1374),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1889),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1891),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1894),
.Y(n_2116)
);

OAI22x1_ASAP7_75t_R g2117 ( 
.A1(n_1886),
.A2(n_1277),
.B1(n_1278),
.B2(n_1269),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1895),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_1898),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_1899),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1900),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1664),
.B(n_1269),
.Y(n_2122)
);

AND2x6_ASAP7_75t_L g2123 ( 
.A(n_1601),
.B(n_735),
.Y(n_2123)
);

CKINVDCx20_ASAP7_75t_R g2124 ( 
.A(n_1583),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1903),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1904),
.Y(n_2126)
);

BUFx6f_ASAP7_75t_L g2127 ( 
.A(n_1910),
.Y(n_2127)
);

AO22x1_ASAP7_75t_L g2128 ( 
.A1(n_1753),
.A2(n_821),
.B1(n_879),
.B2(n_801),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1913),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1914),
.Y(n_2130)
);

BUFx6f_ASAP7_75t_L g2131 ( 
.A(n_1916),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1919),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_1605),
.A2(n_1389),
.B(n_1374),
.Y(n_2133)
);

AND2x4_ASAP7_75t_L g2134 ( 
.A(n_1607),
.B(n_845),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_1920),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1922),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_1926),
.Y(n_2137)
);

AND2x6_ASAP7_75t_L g2138 ( 
.A(n_1608),
.B(n_754),
.Y(n_2138)
);

INVx2_ASAP7_75t_SL g2139 ( 
.A(n_1641),
.Y(n_2139)
);

INVxp33_ASAP7_75t_SL g2140 ( 
.A(n_1642),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1612),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_1745),
.Y(n_2142)
);

AND2x4_ASAP7_75t_L g2143 ( 
.A(n_1613),
.B(n_845),
.Y(n_2143)
);

CKINVDCx8_ASAP7_75t_R g2144 ( 
.A(n_1621),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1614),
.Y(n_2145)
);

CKINVDCx11_ASAP7_75t_R g2146 ( 
.A(n_1892),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1616),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1622),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_1627),
.B(n_852),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_1628),
.Y(n_2150)
);

AND2x4_ASAP7_75t_L g2151 ( 
.A(n_1629),
.B(n_852),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_1631),
.B(n_922),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1632),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1633),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1635),
.B(n_922),
.Y(n_2155)
);

INVx3_ASAP7_75t_L g2156 ( 
.A(n_1636),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1638),
.Y(n_2157)
);

CKINVDCx5p33_ASAP7_75t_R g2158 ( 
.A(n_1642),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1639),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_1665),
.B(n_945),
.Y(n_2160)
);

OA21x2_ASAP7_75t_L g2161 ( 
.A1(n_1666),
.A2(n_1398),
.B(n_1396),
.Y(n_2161)
);

BUFx3_ASAP7_75t_L g2162 ( 
.A(n_1667),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1668),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1669),
.Y(n_2164)
);

BUFx6f_ASAP7_75t_L g2165 ( 
.A(n_1671),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1673),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1675),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1677),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1681),
.Y(n_2169)
);

CKINVDCx20_ASAP7_75t_R g2170 ( 
.A(n_1583),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_1682),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1684),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1685),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1686),
.Y(n_2174)
);

INVx6_ASAP7_75t_L g2175 ( 
.A(n_1773),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1689),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1690),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_1693),
.B(n_1277),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1695),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1696),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_1697),
.B(n_945),
.Y(n_2181)
);

AOI22x1_ASAP7_75t_SL g2182 ( 
.A1(n_1879),
.A2(n_879),
.B1(n_971),
.B2(n_966),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_1698),
.Y(n_2183)
);

INVx3_ASAP7_75t_L g2184 ( 
.A(n_1699),
.Y(n_2184)
);

CKINVDCx5p33_ASAP7_75t_R g2185 ( 
.A(n_1680),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1702),
.Y(n_2186)
);

XOR2xp5_ASAP7_75t_L g2187 ( 
.A(n_1589),
.B(n_1561),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1703),
.Y(n_2188)
);

INVx3_ASAP7_75t_L g2189 ( 
.A(n_1704),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_1680),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_1705),
.A2(n_1398),
.B(n_1396),
.Y(n_2191)
);

HB1xp67_ASAP7_75t_L g2192 ( 
.A(n_1700),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1707),
.Y(n_2193)
);

AND2x2_ASAP7_75t_SL g2194 ( 
.A(n_1730),
.B(n_693),
.Y(n_2194)
);

AND2x4_ASAP7_75t_L g2195 ( 
.A(n_1711),
.B(n_983),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1712),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1713),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1718),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1821),
.B(n_1372),
.Y(n_2199)
);

INVx3_ASAP7_75t_L g2200 ( 
.A(n_1720),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1721),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1723),
.Y(n_2202)
);

OAI22x1_ASAP7_75t_L g2203 ( 
.A1(n_1775),
.A2(n_821),
.B1(n_971),
.B2(n_966),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1724),
.B(n_983),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_1731),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1732),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1733),
.B(n_1002),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1734),
.B(n_1278),
.Y(n_2208)
);

OAI21x1_ASAP7_75t_L g2209 ( 
.A1(n_1735),
.A2(n_1432),
.B(n_1402),
.Y(n_2209)
);

BUFx6f_ASAP7_75t_L g2210 ( 
.A(n_1737),
.Y(n_2210)
);

INVx4_ASAP7_75t_L g2211 ( 
.A(n_1745),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_1738),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1739),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_1741),
.Y(n_2214)
);

OR2x2_ASAP7_75t_L g2215 ( 
.A(n_1875),
.B(n_1279),
.Y(n_2215)
);

INVx3_ASAP7_75t_L g2216 ( 
.A(n_1742),
.Y(n_2216)
);

BUFx8_ASAP7_75t_L g2217 ( 
.A(n_1776),
.Y(n_2217)
);

OAI21x1_ASAP7_75t_L g2218 ( 
.A1(n_1749),
.A2(n_1432),
.B(n_1402),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_1750),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_SL g2220 ( 
.A1(n_1589),
.A2(n_1377),
.B1(n_1408),
.B2(n_1293),
.Y(n_2220)
);

NOR2x1_ASAP7_75t_L g2221 ( 
.A(n_1752),
.B(n_754),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1831),
.B(n_1372),
.Y(n_2222)
);

OAI22x1_ASAP7_75t_R g2223 ( 
.A1(n_1902),
.A2(n_1280),
.B1(n_1281),
.B2(n_1279),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1756),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_1758),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1763),
.Y(n_2226)
);

BUFx6f_ASAP7_75t_L g2227 ( 
.A(n_1765),
.Y(n_2227)
);

NOR2xp33_ASAP7_75t_SL g2228 ( 
.A(n_1726),
.B(n_1280),
.Y(n_2228)
);

BUFx3_ASAP7_75t_L g2229 ( 
.A(n_1767),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1778),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1779),
.B(n_1372),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1781),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1783),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1784),
.A2(n_1445),
.B(n_1434),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1728),
.Y(n_2235)
);

BUFx3_ASAP7_75t_L g2236 ( 
.A(n_1728),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1804),
.B(n_1372),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_SL g2238 ( 
.A(n_1833),
.B(n_1281),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1740),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1740),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1743),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1743),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_1746),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_1746),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1748),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1748),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1755),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1755),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1759),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_1833),
.A2(n_714),
.B1(n_1111),
.B2(n_1039),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1759),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_1768),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1768),
.Y(n_2253)
);

BUFx6f_ASAP7_75t_L g2254 ( 
.A(n_1771),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_1572),
.B(n_1285),
.Y(n_2255)
);

INVx2_ASAP7_75t_L g2256 ( 
.A(n_1771),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1782),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1782),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_1602),
.B(n_1285),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_1662),
.B(n_1002),
.Y(n_2260)
);

NAND2xp33_ASAP7_75t_L g2261 ( 
.A(n_1838),
.B(n_832),
.Y(n_2261)
);

XNOR2x2_ASAP7_75t_L g2262 ( 
.A(n_1826),
.B(n_1012),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_1785),
.Y(n_2263)
);

BUFx2_ASAP7_75t_L g2264 ( 
.A(n_1911),
.Y(n_2264)
);

BUFx8_ASAP7_75t_SL g2265 ( 
.A(n_1615),
.Y(n_2265)
);

AOI22xp5_ASAP7_75t_L g2266 ( 
.A1(n_1838),
.A2(n_1041),
.B1(n_1120),
.B2(n_1012),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1785),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_1786),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_1660),
.B(n_1291),
.Y(n_2269)
);

OAI22x1_ASAP7_75t_SL g2270 ( 
.A1(n_1911),
.A2(n_1292),
.B1(n_1293),
.B2(n_1291),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1877),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1688),
.Y(n_2272)
);

CKINVDCx5p33_ASAP7_75t_R g2273 ( 
.A(n_1807),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1701),
.Y(n_2274)
);

OAI21x1_ASAP7_75t_L g2275 ( 
.A1(n_1770),
.A2(n_1445),
.B(n_1434),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1897),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1848),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1824),
.Y(n_2278)
);

BUFx6f_ASAP7_75t_L g2279 ( 
.A(n_1848),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1888),
.B(n_1372),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1850),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_1708),
.Y(n_2282)
);

BUFx12f_ASAP7_75t_L g2283 ( 
.A(n_1710),
.Y(n_2283)
);

BUFx8_ASAP7_75t_SL g2284 ( 
.A(n_1615),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1878),
.Y(n_2285)
);

INVx5_ASAP7_75t_L g2286 ( 
.A(n_1760),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1905),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1924),
.Y(n_2288)
);

BUFx2_ASAP7_75t_L g2289 ( 
.A(n_1921),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1850),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_1852),
.Y(n_2291)
);

INVx4_ASAP7_75t_L g2292 ( 
.A(n_1852),
.Y(n_2292)
);

BUFx12f_ASAP7_75t_L g2293 ( 
.A(n_1862),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_1907),
.A2(n_1618),
.B1(n_1597),
.B2(n_1603),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_1862),
.Y(n_2295)
);

OA21x2_ASAP7_75t_L g2296 ( 
.A1(n_1864),
.A2(n_1455),
.B(n_1454),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_1646),
.B(n_1725),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1925),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1864),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1865),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1869),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1927),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_1869),
.B(n_1099),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1870),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_1870),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_1921),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1893),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_1928),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1893),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_1908),
.Y(n_2310)
);

CKINVDCx16_ASAP7_75t_R g2311 ( 
.A(n_1761),
.Y(n_2311)
);

BUFx3_ASAP7_75t_L g2312 ( 
.A(n_1908),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1915),
.Y(n_2313)
);

BUFx6f_ASAP7_75t_L g2314 ( 
.A(n_1915),
.Y(n_2314)
);

OA21x2_ASAP7_75t_L g2315 ( 
.A1(n_1918),
.A2(n_1455),
.B(n_1454),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1814),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_1747),
.B(n_1292),
.Y(n_2317)
);

INVx5_ASAP7_75t_L g2318 ( 
.A(n_1764),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_1918),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1923),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_1923),
.B(n_1296),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1597),
.Y(n_2322)
);

BUFx12f_ASAP7_75t_L g2323 ( 
.A(n_1603),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1620),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1888),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_1928),
.B(n_1099),
.Y(n_2326)
);

AND2x4_ASAP7_75t_L g2327 ( 
.A(n_1847),
.B(n_755),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1774),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_1839),
.B(n_1296),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1857),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_1823),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1942),
.B(n_2042),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2141),
.Y(n_2333)
);

AND2x6_ASAP7_75t_L g2334 ( 
.A(n_2297),
.B(n_755),
.Y(n_2334)
);

INVxp67_ASAP7_75t_SL g2335 ( 
.A(n_1965),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2141),
.Y(n_2336)
);

CKINVDCx5p33_ASAP7_75t_R g2337 ( 
.A(n_1953),
.Y(n_2337)
);

NAND2xp33_ASAP7_75t_SL g2338 ( 
.A(n_2242),
.B(n_1363),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_1953),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2154),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_1945),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_2010),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2154),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2159),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1942),
.B(n_1956),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2159),
.Y(n_2346)
);

HB1xp67_ASAP7_75t_L g2347 ( 
.A(n_1935),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2163),
.Y(n_2348)
);

CKINVDCx20_ASAP7_75t_R g2349 ( 
.A(n_2124),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2163),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_1935),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2297),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2172),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2191),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_1940),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_2010),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2215),
.B(n_1618),
.Y(n_2357)
);

CKINVDCx5p33_ASAP7_75t_R g2358 ( 
.A(n_2076),
.Y(n_2358)
);

OA21x2_ASAP7_75t_L g2359 ( 
.A1(n_1936),
.A2(n_1526),
.B(n_1493),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_1938),
.B(n_1843),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_L g2361 ( 
.A(n_2215),
.B(n_1645),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_2076),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2172),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2173),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2191),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1956),
.B(n_1363),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2209),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2255),
.B(n_2259),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2173),
.Y(n_2369)
);

INVx3_ASAP7_75t_L g2370 ( 
.A(n_1945),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2100),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_1940),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2174),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2174),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2218),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2286),
.B(n_756),
.Y(n_2376)
);

HB1xp67_ASAP7_75t_L g2377 ( 
.A(n_1938),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_R g2378 ( 
.A(n_2158),
.B(n_1866),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2158),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2286),
.B(n_756),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2255),
.B(n_1366),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2176),
.Y(n_2382)
);

CKINVDCx5p33_ASAP7_75t_R g2383 ( 
.A(n_2185),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2176),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2197),
.Y(n_2385)
);

CKINVDCx20_ASAP7_75t_R g2386 ( 
.A(n_2170),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2197),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2218),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2201),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_1940),
.Y(n_2390)
);

XOR2xp5_ASAP7_75t_L g2391 ( 
.A(n_2187),
.B(n_2185),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2234),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2201),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2226),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2226),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_2251),
.Y(n_2396)
);

NOR2xp33_ASAP7_75t_R g2397 ( 
.A(n_2251),
.B(n_1866),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2286),
.Y(n_2398)
);

BUFx10_ASAP7_75t_L g2399 ( 
.A(n_2088),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2234),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2230),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2230),
.Y(n_2402)
);

CKINVDCx20_ASAP7_75t_R g2403 ( 
.A(n_1937),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1994),
.Y(n_2404)
);

BUFx3_ASAP7_75t_L g2405 ( 
.A(n_2286),
.Y(n_2405)
);

CKINVDCx20_ASAP7_75t_R g2406 ( 
.A(n_1951),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_2268),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_1994),
.Y(n_2408)
);

INVx3_ASAP7_75t_L g2409 ( 
.A(n_1945),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1930),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2268),
.Y(n_2411)
);

CKINVDCx5p33_ASAP7_75t_R g2412 ( 
.A(n_2015),
.Y(n_2412)
);

BUFx6f_ASAP7_75t_L g2413 ( 
.A(n_1940),
.Y(n_2413)
);

BUFx8_ASAP7_75t_L g2414 ( 
.A(n_2264),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1956),
.B(n_1366),
.Y(n_2415)
);

CKINVDCx5p33_ASAP7_75t_R g2416 ( 
.A(n_2020),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_1994),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2286),
.B(n_758),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2265),
.Y(n_2419)
);

CKINVDCx20_ASAP7_75t_R g2420 ( 
.A(n_2284),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1956),
.B(n_1377),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_R g2422 ( 
.A(n_2273),
.B(n_1751),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2286),
.B(n_758),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1930),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_1933),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_2011),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_2011),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_1945),
.Y(n_2428)
);

CKINVDCx20_ASAP7_75t_R g2429 ( 
.A(n_2187),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_1994),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_1940),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2018),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_2318),
.B(n_759),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1933),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_1947),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2184),
.B(n_2189),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2259),
.B(n_1382),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2018),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1947),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2140),
.Y(n_2440)
);

CKINVDCx20_ASAP7_75t_R g2441 ( 
.A(n_2086),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2018),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2018),
.Y(n_2443)
);

AND2x4_ASAP7_75t_L g2444 ( 
.A(n_2318),
.B(n_759),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_2012),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1954),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2184),
.B(n_1382),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_SL g2448 ( 
.A(n_2279),
.B(n_1650),
.Y(n_2448)
);

BUFx8_ASAP7_75t_L g2449 ( 
.A(n_2264),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_1963),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2039),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_1954),
.Y(n_2452)
);

XNOR2x2_ASAP7_75t_L g2453 ( 
.A(n_2262),
.B(n_1039),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2269),
.B(n_1383),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2039),
.Y(n_2455)
);

OAI21x1_ASAP7_75t_L g2456 ( 
.A1(n_1967),
.A2(n_1137),
.B(n_1130),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2269),
.B(n_1383),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2039),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_1972),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_1977),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2089),
.B(n_1650),
.Y(n_2461)
);

BUFx2_ASAP7_75t_L g2462 ( 
.A(n_1977),
.Y(n_2462)
);

CKINVDCx20_ASAP7_75t_R g2463 ( 
.A(n_2086),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_1979),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_2012),
.Y(n_2465)
);

CKINVDCx5p33_ASAP7_75t_R g2466 ( 
.A(n_2058),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_1972),
.Y(n_2467)
);

HB1xp67_ASAP7_75t_L g2468 ( 
.A(n_1979),
.Y(n_2468)
);

CKINVDCx20_ASAP7_75t_R g2469 ( 
.A(n_2146),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2184),
.B(n_1385),
.Y(n_2470)
);

HB1xp67_ASAP7_75t_L g2471 ( 
.A(n_2013),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_1967),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1986),
.Y(n_2473)
);

INVx3_ASAP7_75t_L g2474 ( 
.A(n_2161),
.Y(n_2474)
);

CKINVDCx5p33_ASAP7_75t_R g2475 ( 
.A(n_2085),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_1986),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2085),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_1995),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_1964),
.Y(n_2479)
);

INVxp33_ASAP7_75t_L g2480 ( 
.A(n_2117),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_1963),
.Y(n_2481)
);

BUFx8_ASAP7_75t_L g2482 ( 
.A(n_2289),
.Y(n_2482)
);

NOR2xp33_ASAP7_75t_R g2483 ( 
.A(n_2273),
.B(n_2316),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_1964),
.Y(n_2484)
);

BUFx8_ASAP7_75t_L g2485 ( 
.A(n_2289),
.Y(n_2485)
);

AND2x4_ASAP7_75t_L g2486 ( 
.A(n_2318),
.B(n_765),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1990),
.Y(n_2487)
);

AND3x2_ASAP7_75t_L g2488 ( 
.A(n_2228),
.B(n_1111),
.C(n_1643),
.Y(n_2488)
);

BUFx6f_ASAP7_75t_L g2489 ( 
.A(n_1963),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_1995),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_2279),
.B(n_1788),
.Y(n_2491)
);

BUFx2_ASAP7_75t_L g2492 ( 
.A(n_2013),
.Y(n_2492)
);

BUFx6f_ASAP7_75t_L g2493 ( 
.A(n_1963),
.Y(n_2493)
);

BUFx2_ASAP7_75t_L g2494 ( 
.A(n_2316),
.Y(n_2494)
);

BUFx6f_ASAP7_75t_L g2495 ( 
.A(n_1963),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_1990),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_1991),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2321),
.B(n_1395),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2009),
.Y(n_2499)
);

CKINVDCx5p33_ASAP7_75t_R g2500 ( 
.A(n_1987),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2063),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2321),
.B(n_1397),
.Y(n_2502)
);

BUFx12f_ASAP7_75t_L g2503 ( 
.A(n_1957),
.Y(n_2503)
);

CKINVDCx20_ASAP7_75t_R g2504 ( 
.A(n_2104),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_1991),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2094),
.B(n_1397),
.Y(n_2506)
);

CKINVDCx20_ASAP7_75t_R g2507 ( 
.A(n_2104),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1992),
.Y(n_2508)
);

INVxp67_ASAP7_75t_L g2509 ( 
.A(n_2192),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_1987),
.Y(n_2510)
);

CKINVDCx5p33_ASAP7_75t_R g2511 ( 
.A(n_2006),
.Y(n_2511)
);

BUFx3_ASAP7_75t_L g2512 ( 
.A(n_2318),
.Y(n_2512)
);

HB1xp67_ASAP7_75t_L g2513 ( 
.A(n_1998),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2063),
.Y(n_2514)
);

CKINVDCx16_ASAP7_75t_R g2515 ( 
.A(n_2311),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_2006),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_1992),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2133),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2014),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2008),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2014),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2016),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2161),
.Y(n_2523)
);

CKINVDCx20_ASAP7_75t_R g2524 ( 
.A(n_2311),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_SL g2525 ( 
.A1(n_2106),
.A2(n_1644),
.B1(n_1649),
.B2(n_1643),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2008),
.Y(n_2526)
);

OAI21x1_ASAP7_75t_L g2527 ( 
.A1(n_1936),
.A2(n_2133),
.B(n_2059),
.Y(n_2527)
);

NOR2xp67_ASAP7_75t_L g2528 ( 
.A(n_2318),
.B(n_1401),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_2293),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2318),
.B(n_765),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2161),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2016),
.Y(n_2532)
);

CKINVDCx16_ASAP7_75t_R g2533 ( 
.A(n_2117),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2019),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2277),
.B(n_1803),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2019),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2022),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_2293),
.Y(n_2538)
);

BUFx10_ASAP7_75t_L g2539 ( 
.A(n_2029),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2113),
.Y(n_2540)
);

HB1xp67_ASAP7_75t_L g2541 ( 
.A(n_2003),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2113),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2283),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2022),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2283),
.Y(n_2545)
);

BUFx3_ASAP7_75t_L g2546 ( 
.A(n_2236),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2026),
.Y(n_2547)
);

AND2x6_ASAP7_75t_L g2548 ( 
.A(n_1946),
.B(n_766),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_2323),
.Y(n_2549)
);

AND2x4_ASAP7_75t_L g2550 ( 
.A(n_2236),
.B(n_766),
.Y(n_2550)
);

AND3x1_ASAP7_75t_L g2551 ( 
.A(n_1939),
.B(n_772),
.C(n_769),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2026),
.Y(n_2552)
);

CKINVDCx5p33_ASAP7_75t_R g2553 ( 
.A(n_2323),
.Y(n_2553)
);

OAI22xp5_ASAP7_75t_SL g2554 ( 
.A1(n_2106),
.A2(n_1649),
.B1(n_1652),
.B2(n_1644),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_1934),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_1934),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_2032),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_1948),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_1948),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2028),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2028),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2113),
.Y(n_2562)
);

BUFx2_ASAP7_75t_L g2563 ( 
.A(n_2312),
.Y(n_2563)
);

CKINVDCx20_ASAP7_75t_R g2564 ( 
.A(n_2223),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2049),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_2161),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2200),
.B(n_1408),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2277),
.B(n_1813),
.Y(n_2568)
);

CKINVDCx20_ASAP7_75t_R g2569 ( 
.A(n_2223),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2049),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2057),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2057),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2017),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_1973),
.Y(n_2574)
);

BUFx2_ASAP7_75t_L g2575 ( 
.A(n_2312),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2071),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2113),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_1973),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2236),
.Y(n_2579)
);

NAND2xp5_ASAP7_75t_L g2580 ( 
.A(n_2200),
.B(n_1409),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2071),
.Y(n_2581)
);

AND2x2_ASAP7_75t_L g2582 ( 
.A(n_2282),
.B(n_1409),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2074),
.Y(n_2583)
);

BUFx6f_ASAP7_75t_L g2584 ( 
.A(n_1973),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2074),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2092),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2092),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2099),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_R g2589 ( 
.A(n_1984),
.B(n_1787),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_1931),
.Y(n_2590)
);

HB1xp67_ASAP7_75t_L g2591 ( 
.A(n_2062),
.Y(n_2591)
);

INVxp67_ASAP7_75t_L g2592 ( 
.A(n_2306),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2099),
.Y(n_2593)
);

CKINVDCx5p33_ASAP7_75t_R g2594 ( 
.A(n_2244),
.Y(n_2594)
);

BUFx6f_ASAP7_75t_L g2595 ( 
.A(n_1973),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2244),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2102),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_2244),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_1931),
.Y(n_2599)
);

BUFx2_ASAP7_75t_L g2600 ( 
.A(n_2312),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_1932),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2306),
.Y(n_2602)
);

CKINVDCx5p33_ASAP7_75t_R g2603 ( 
.A(n_1957),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_1957),
.Y(n_2604)
);

INVx1_ASAP7_75t_SL g2605 ( 
.A(n_2308),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2200),
.B(n_1412),
.Y(n_2606)
);

CKINVDCx5p33_ASAP7_75t_R g2607 ( 
.A(n_1957),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2001),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2102),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_1932),
.Y(n_2610)
);

BUFx6f_ASAP7_75t_L g2611 ( 
.A(n_1973),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2317),
.B(n_1412),
.Y(n_2612)
);

NOR2xp67_ASAP7_75t_L g2613 ( 
.A(n_1984),
.B(n_1413),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2105),
.Y(n_2614)
);

INVx3_ASAP7_75t_L g2615 ( 
.A(n_2001),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2279),
.B(n_1816),
.Y(n_2616)
);

BUFx2_ASAP7_75t_L g2617 ( 
.A(n_2308),
.Y(n_2617)
);

CKINVDCx5p33_ASAP7_75t_R g2618 ( 
.A(n_1962),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2105),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_1962),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2317),
.B(n_1413),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_1962),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2111),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_1941),
.Y(n_2624)
);

AND2x2_ASAP7_75t_L g2625 ( 
.A(n_2000),
.B(n_1414),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_1962),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_1996),
.Y(n_2627)
);

CKINVDCx20_ASAP7_75t_R g2628 ( 
.A(n_2004),
.Y(n_2628)
);

CKINVDCx5p33_ASAP7_75t_R g2629 ( 
.A(n_1996),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2111),
.Y(n_2630)
);

CKINVDCx20_ASAP7_75t_R g2631 ( 
.A(n_2004),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2115),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2115),
.Y(n_2633)
);

CKINVDCx6p67_ASAP7_75t_R g2634 ( 
.A(n_2194),
.Y(n_2634)
);

CKINVDCx5p33_ASAP7_75t_R g2635 ( 
.A(n_1971),
.Y(n_2635)
);

CKINVDCx5p33_ASAP7_75t_R g2636 ( 
.A(n_1971),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2000),
.B(n_1414),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_1971),
.Y(n_2638)
);

INVx4_ASAP7_75t_L g2639 ( 
.A(n_2175),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2279),
.B(n_1816),
.Y(n_2640)
);

CKINVDCx20_ASAP7_75t_R g2641 ( 
.A(n_1950),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2005),
.B(n_1416),
.Y(n_2642)
);

CKINVDCx20_ASAP7_75t_R g2643 ( 
.A(n_1950),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2200),
.B(n_1416),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2121),
.Y(n_2645)
);

BUFx2_ASAP7_75t_L g2646 ( 
.A(n_1971),
.Y(n_2646)
);

BUFx3_ASAP7_75t_L g2647 ( 
.A(n_1978),
.Y(n_2647)
);

CKINVDCx20_ASAP7_75t_R g2648 ( 
.A(n_1980),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2281),
.B(n_1418),
.Y(n_2649)
);

OA21x2_ASAP7_75t_L g2650 ( 
.A1(n_2275),
.A2(n_1526),
.B(n_1493),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_1980),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2121),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_1980),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2129),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_1980),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2001),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_2001),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2242),
.B(n_769),
.Y(n_2658)
);

CKINVDCx5p33_ASAP7_75t_R g2659 ( 
.A(n_2217),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2216),
.B(n_2224),
.Y(n_2660)
);

AND2x4_ASAP7_75t_L g2661 ( 
.A(n_2242),
.B(n_772),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_1941),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2129),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2034),
.Y(n_2664)
);

CKINVDCx20_ASAP7_75t_R g2665 ( 
.A(n_2217),
.Y(n_2665)
);

CKINVDCx5p33_ASAP7_75t_R g2666 ( 
.A(n_2217),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2216),
.B(n_1418),
.Y(n_2667)
);

AND3x2_ASAP7_75t_L g2668 ( 
.A(n_1966),
.B(n_1655),
.C(n_1652),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2034),
.Y(n_2669)
);

INVx3_ASAP7_75t_L g2670 ( 
.A(n_2001),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_1943),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_1997),
.Y(n_2672)
);

NOR2xp67_ASAP7_75t_L g2673 ( 
.A(n_2292),
.B(n_1420),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2145),
.Y(n_2674)
);

CKINVDCx5p33_ASAP7_75t_R g2675 ( 
.A(n_2217),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2145),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2147),
.Y(n_2677)
);

INVxp67_ASAP7_75t_L g2678 ( 
.A(n_2005),
.Y(n_2678)
);

HB1xp67_ASAP7_75t_L g2679 ( 
.A(n_2331),
.Y(n_2679)
);

INVx3_ASAP7_75t_L g2680 ( 
.A(n_2002),
.Y(n_2680)
);

HB1xp67_ASAP7_75t_L g2681 ( 
.A(n_2331),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_1943),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2148),
.Y(n_2683)
);

BUFx2_ASAP7_75t_L g2684 ( 
.A(n_2194),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2150),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_2294),
.Y(n_2686)
);

NOR2xp33_ASAP7_75t_R g2687 ( 
.A(n_2144),
.B(n_1715),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2144),
.Y(n_2688)
);

CKINVDCx5p33_ASAP7_75t_R g2689 ( 
.A(n_2242),
.Y(n_2689)
);

BUFx3_ASAP7_75t_L g2690 ( 
.A(n_1978),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2150),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2153),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2153),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2021),
.Y(n_2694)
);

CKINVDCx16_ASAP7_75t_R g2695 ( 
.A(n_2329),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2021),
.Y(n_2696)
);

NOR2xp33_ASAP7_75t_L g2697 ( 
.A(n_2281),
.B(n_1420),
.Y(n_2697)
);

CKINVDCx5p33_ASAP7_75t_R g2698 ( 
.A(n_2242),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2139),
.B(n_1421),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2037),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2254),
.Y(n_2701)
);

AND2x2_ASAP7_75t_L g2702 ( 
.A(n_2139),
.B(n_1421),
.Y(n_2702)
);

INVx3_ASAP7_75t_L g2703 ( 
.A(n_2002),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2216),
.B(n_1426),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2037),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_2254),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2051),
.Y(n_2707)
);

CKINVDCx20_ASAP7_75t_R g2708 ( 
.A(n_2220),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2051),
.Y(n_2709)
);

CKINVDCx5p33_ASAP7_75t_R g2710 ( 
.A(n_2254),
.Y(n_2710)
);

CKINVDCx16_ASAP7_75t_R g2711 ( 
.A(n_2329),
.Y(n_2711)
);

NOR2xp33_ASAP7_75t_R g2712 ( 
.A(n_2190),
.B(n_1717),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_2254),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2216),
.B(n_1426),
.Y(n_2714)
);

NOR2xp33_ASAP7_75t_L g2715 ( 
.A(n_2290),
.B(n_1428),
.Y(n_2715)
);

INVxp33_ASAP7_75t_L g2716 ( 
.A(n_2220),
.Y(n_2716)
);

HB1xp67_ASAP7_75t_L g2717 ( 
.A(n_2331),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2072),
.Y(n_2718)
);

BUFx6f_ASAP7_75t_L g2719 ( 
.A(n_1997),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2190),
.B(n_1428),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_SL g2721 ( 
.A(n_2279),
.B(n_1456),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2254),
.Y(n_2722)
);

CKINVDCx5p33_ASAP7_75t_R g2723 ( 
.A(n_2270),
.Y(n_2723)
);

CKINVDCx20_ASAP7_75t_R g2724 ( 
.A(n_1939),
.Y(n_2724)
);

INVxp67_ASAP7_75t_L g2725 ( 
.A(n_2295),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_1949),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2002),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2072),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2270),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_L g2730 ( 
.A(n_2224),
.B(n_1440),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2166),
.Y(n_2731)
);

CKINVDCx5p33_ASAP7_75t_R g2732 ( 
.A(n_2295),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_1949),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_1959),
.Y(n_2734)
);

AND2x6_ASAP7_75t_L g2735 ( 
.A(n_1946),
.B(n_774),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2327),
.B(n_1440),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2224),
.B(n_1443),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_1959),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_1960),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2331),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2166),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2325),
.B(n_1443),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_1960),
.Y(n_2743)
);

AND2x4_ASAP7_75t_L g2744 ( 
.A(n_2252),
.B(n_774),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2167),
.Y(n_2745)
);

BUFx3_ASAP7_75t_L g2746 ( 
.A(n_1978),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_2295),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_1974),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2295),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2167),
.Y(n_2750)
);

CKINVDCx20_ASAP7_75t_R g2751 ( 
.A(n_2295),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2314),
.Y(n_2752)
);

INVx3_ASAP7_75t_L g2753 ( 
.A(n_2002),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2224),
.B(n_1446),
.Y(n_2754)
);

INVx1_ASAP7_75t_SL g2755 ( 
.A(n_2328),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2168),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_1978),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2314),
.Y(n_2758)
);

NAND2xp33_ASAP7_75t_R g2759 ( 
.A(n_2243),
.B(n_1446),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2327),
.B(n_2075),
.Y(n_2760)
);

AND2x4_ASAP7_75t_L g2761 ( 
.A(n_2252),
.B(n_775),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_2314),
.Y(n_2762)
);

INVx3_ASAP7_75t_L g2763 ( 
.A(n_2002),
.Y(n_2763)
);

AOI22xp33_ASAP7_75t_L g2764 ( 
.A1(n_2760),
.A2(n_2194),
.B1(n_2079),
.B2(n_2327),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2404),
.Y(n_2765)
);

NOR2xp33_ASAP7_75t_L g2766 ( 
.A(n_2357),
.B(n_2325),
.Y(n_2766)
);

BUFx3_ASAP7_75t_L g2767 ( 
.A(n_2398),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2333),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2404),
.Y(n_2769)
);

NAND3xp33_ASAP7_75t_L g2770 ( 
.A(n_2649),
.B(n_2715),
.C(n_2697),
.Y(n_2770)
);

NAND3xp33_ASAP7_75t_L g2771 ( 
.A(n_2535),
.B(n_2319),
.C(n_2314),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2351),
.B(n_2328),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2462),
.B(n_2330),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2336),
.Y(n_2774)
);

BUFx3_ASAP7_75t_L g2775 ( 
.A(n_2398),
.Y(n_2775)
);

AO21x2_ASAP7_75t_L g2776 ( 
.A1(n_2540),
.A2(n_2275),
.B(n_2237),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_SL g2777 ( 
.A(n_2689),
.B(n_2314),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2340),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_SL g2779 ( 
.A(n_2689),
.B(n_2319),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2343),
.Y(n_2780)
);

INVx2_ASAP7_75t_L g2781 ( 
.A(n_2408),
.Y(n_2781)
);

BUFx2_ASAP7_75t_L g2782 ( 
.A(n_2492),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2344),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2346),
.Y(n_2784)
);

INVx3_ASAP7_75t_L g2785 ( 
.A(n_2639),
.Y(n_2785)
);

OAI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2345),
.A2(n_2280),
.B1(n_2252),
.B2(n_2300),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2590),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_SL g2788 ( 
.A(n_2698),
.B(n_2319),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2590),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2599),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2368),
.B(n_2252),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2599),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2332),
.B(n_2300),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2601),
.Y(n_2794)
);

INVx5_ASAP7_75t_L g2795 ( 
.A(n_2548),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2348),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_SL g2797 ( 
.A(n_2698),
.B(n_2319),
.Y(n_2797)
);

INVx2_ASAP7_75t_SL g2798 ( 
.A(n_2639),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2350),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2744),
.B(n_2300),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2601),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_2610),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2353),
.Y(n_2803)
);

AND2x6_ASAP7_75t_L g2804 ( 
.A(n_2405),
.B(n_2320),
.Y(n_2804)
);

BUFx2_ASAP7_75t_L g2805 ( 
.A(n_2471),
.Y(n_2805)
);

INVxp33_ASAP7_75t_L g2806 ( 
.A(n_2422),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2664),
.B(n_2305),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_SL g2808 ( 
.A(n_2701),
.B(n_2320),
.Y(n_2808)
);

AND2x2_ASAP7_75t_SL g2809 ( 
.A(n_2551),
.B(n_2142),
.Y(n_2809)
);

NAND2xp33_ASAP7_75t_L g2810 ( 
.A(n_2732),
.B(n_2320),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2361),
.B(n_2243),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2363),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2364),
.Y(n_2813)
);

BUFx6f_ASAP7_75t_SL g2814 ( 
.A(n_2352),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_2610),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2624),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2744),
.B(n_2761),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2624),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2744),
.B(n_2305),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2662),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2761),
.B(n_2305),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2662),
.Y(n_2822)
);

INVx2_ASAP7_75t_SL g2823 ( 
.A(n_2639),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_2461),
.B(n_2292),
.Y(n_2824)
);

INVx2_ASAP7_75t_L g2825 ( 
.A(n_2671),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2671),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2369),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2568),
.B(n_2292),
.Y(n_2828)
);

INVx1_ASAP7_75t_SL g2829 ( 
.A(n_2347),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2682),
.Y(n_2830)
);

INVx2_ASAP7_75t_SL g2831 ( 
.A(n_2546),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2682),
.Y(n_2832)
);

INVx2_ASAP7_75t_L g2833 ( 
.A(n_2726),
.Y(n_2833)
);

INVx1_ASAP7_75t_SL g2834 ( 
.A(n_2360),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2761),
.B(n_2658),
.Y(n_2835)
);

BUFx3_ASAP7_75t_L g2836 ( 
.A(n_2405),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2726),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2733),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2373),
.Y(n_2839)
);

BUFx6f_ASAP7_75t_L g2840 ( 
.A(n_2450),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2733),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2450),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_L g2843 ( 
.A(n_2337),
.B(n_2292),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2374),
.Y(n_2844)
);

NAND3xp33_ASAP7_75t_L g2845 ( 
.A(n_2759),
.B(n_2320),
.C(n_2307),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2382),
.Y(n_2846)
);

INVx3_ASAP7_75t_L g2847 ( 
.A(n_2450),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2384),
.Y(n_2848)
);

BUFx3_ASAP7_75t_L g2849 ( 
.A(n_2512),
.Y(n_2849)
);

AOI21x1_ASAP7_75t_L g2850 ( 
.A1(n_2354),
.A2(n_2367),
.B(n_2365),
.Y(n_2850)
);

OR2x2_ASAP7_75t_L g2851 ( 
.A(n_2515),
.B(n_2330),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2658),
.B(n_1968),
.Y(n_2852)
);

AND2x2_ASAP7_75t_SL g2853 ( 
.A(n_2533),
.B(n_2142),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_SL g2854 ( 
.A(n_2701),
.B(n_2271),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_L g2855 ( 
.A(n_2450),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_2734),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2734),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2658),
.B(n_1968),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2385),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_2337),
.B(n_2235),
.Y(n_2860)
);

INVxp67_ASAP7_75t_SL g2861 ( 
.A(n_2647),
.Y(n_2861)
);

INVx5_ASAP7_75t_L g2862 ( 
.A(n_2548),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2738),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2661),
.B(n_1968),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2387),
.Y(n_2865)
);

INVx2_ASAP7_75t_SL g2866 ( 
.A(n_2546),
.Y(n_2866)
);

OAI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2686),
.A2(n_2724),
.B1(n_2594),
.B2(n_2596),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2738),
.Y(n_2868)
);

INVx2_ASAP7_75t_L g2869 ( 
.A(n_2739),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2739),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2661),
.B(n_2290),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2743),
.Y(n_2872)
);

INVx8_ASAP7_75t_L g2873 ( 
.A(n_2548),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2661),
.B(n_2291),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_SL g2875 ( 
.A(n_2706),
.B(n_2271),
.Y(n_2875)
);

OAI22xp33_ASAP7_75t_L g2876 ( 
.A1(n_2686),
.A2(n_2091),
.B1(n_2266),
.B2(n_2271),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2389),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2339),
.B(n_2241),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_SL g2879 ( 
.A(n_2706),
.B(n_2271),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2625),
.B(n_2637),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2366),
.B(n_2415),
.Y(n_2881)
);

INVx2_ASAP7_75t_L g2882 ( 
.A(n_2743),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2421),
.B(n_2291),
.Y(n_2883)
);

BUFx10_ASAP7_75t_L g2884 ( 
.A(n_2555),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2710),
.B(n_2271),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_SL g2886 ( 
.A(n_2710),
.B(n_2239),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2349),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2748),
.Y(n_2888)
);

INVxp67_ASAP7_75t_SL g2889 ( 
.A(n_2647),
.Y(n_2889)
);

BUFx6f_ASAP7_75t_SL g2890 ( 
.A(n_2352),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2481),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2393),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2394),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2395),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2669),
.B(n_2299),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2401),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2748),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2408),
.Y(n_2898)
);

CKINVDCx6p67_ASAP7_75t_R g2899 ( 
.A(n_2403),
.Y(n_2899)
);

INVx5_ASAP7_75t_L g2900 ( 
.A(n_2548),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2417),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2724),
.A2(n_2073),
.B1(n_2123),
.B2(n_2054),
.Y(n_2902)
);

AOI21x1_ASAP7_75t_L g2903 ( 
.A1(n_2354),
.A2(n_2231),
.B(n_1981),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2417),
.Y(n_2904)
);

INVx8_ASAP7_75t_L g2905 ( 
.A(n_2548),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2430),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2430),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2447),
.B(n_2470),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2402),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2432),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2432),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2438),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2736),
.B(n_2075),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2481),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2713),
.B(n_2239),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_SL g2916 ( 
.A(n_2713),
.B(n_2240),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2410),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_SL g2918 ( 
.A(n_2722),
.B(n_2240),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2438),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2424),
.Y(n_2920)
);

INVxp67_ASAP7_75t_L g2921 ( 
.A(n_2377),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2442),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_SL g2923 ( 
.A(n_2334),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2442),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2425),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2443),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2722),
.B(n_2253),
.Y(n_2927)
);

CKINVDCx5p33_ASAP7_75t_R g2928 ( 
.A(n_2483),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2434),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2443),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_L g2931 ( 
.A(n_2342),
.B(n_2245),
.Y(n_2931)
);

BUFx6f_ASAP7_75t_SL g2932 ( 
.A(n_2334),
.Y(n_2932)
);

INVxp67_ASAP7_75t_L g2933 ( 
.A(n_2460),
.Y(n_2933)
);

INVx8_ASAP7_75t_L g2934 ( 
.A(n_2548),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2451),
.Y(n_2935)
);

CKINVDCx11_ASAP7_75t_R g2936 ( 
.A(n_2403),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2435),
.Y(n_2937)
);

NOR2xp33_ASAP7_75t_L g2938 ( 
.A(n_2356),
.B(n_2245),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2455),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2439),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_2747),
.B(n_2256),
.Y(n_2941)
);

INVx2_ASAP7_75t_L g2942 ( 
.A(n_2455),
.Y(n_2942)
);

BUFx4f_ASAP7_75t_L g2943 ( 
.A(n_2634),
.Y(n_2943)
);

CKINVDCx5p33_ASAP7_75t_R g2944 ( 
.A(n_2378),
.Y(n_2944)
);

BUFx2_ASAP7_75t_L g2945 ( 
.A(n_2349),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2446),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2458),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2694),
.B(n_2122),
.Y(n_2948)
);

INVx8_ASAP7_75t_L g2949 ( 
.A(n_2735),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2458),
.Y(n_2950)
);

INVx1_ASAP7_75t_SL g2951 ( 
.A(n_2605),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2542),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2542),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2452),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2386),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2562),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2562),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2356),
.B(n_2246),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2459),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_SL g2960 ( 
.A(n_2747),
.B(n_2256),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2749),
.B(n_2257),
.Y(n_2961)
);

INVx1_ASAP7_75t_SL g2962 ( 
.A(n_2386),
.Y(n_2962)
);

AOI22xp5_ASAP7_75t_L g2963 ( 
.A1(n_2735),
.A2(n_2751),
.B1(n_2073),
.B2(n_2123),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2577),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_2481),
.Y(n_2965)
);

INVx2_ASAP7_75t_L g2966 ( 
.A(n_2577),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2749),
.B(n_2257),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2467),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2474),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2473),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2474),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2474),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2752),
.B(n_2258),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_SL g2974 ( 
.A(n_2752),
.B(n_2258),
.Y(n_2974)
);

INVx3_ASAP7_75t_L g2975 ( 
.A(n_2481),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2523),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2476),
.Y(n_2977)
);

BUFx6f_ASAP7_75t_L g2978 ( 
.A(n_2489),
.Y(n_2978)
);

INVx2_ASAP7_75t_SL g2979 ( 
.A(n_2690),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2531),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_SL g2981 ( 
.A(n_2758),
.B(n_2263),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2531),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_SL g2983 ( 
.A(n_2758),
.B(n_2762),
.Y(n_2983)
);

XNOR2xp5_ASAP7_75t_L g2984 ( 
.A(n_2525),
.B(n_1655),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2487),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_SL g2986 ( 
.A(n_2762),
.B(n_2263),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_SL g2987 ( 
.A(n_2579),
.B(n_2267),
.Y(n_2987)
);

INVx2_ASAP7_75t_L g2988 ( 
.A(n_2531),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2579),
.B(n_2267),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2566),
.Y(n_2990)
);

INVx2_ASAP7_75t_SL g2991 ( 
.A(n_2690),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2496),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2696),
.B(n_2700),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2566),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2497),
.Y(n_2995)
);

INVx2_ASAP7_75t_SL g2996 ( 
.A(n_2746),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2505),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2594),
.B(n_2301),
.Y(n_2998)
);

INVx2_ASAP7_75t_SL g2999 ( 
.A(n_2746),
.Y(n_2999)
);

OR2x2_ASAP7_75t_L g3000 ( 
.A(n_2695),
.B(n_2272),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2508),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2566),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2341),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2341),
.Y(n_3004)
);

NAND3xp33_ASAP7_75t_L g3005 ( 
.A(n_2567),
.B(n_2606),
.C(n_2580),
.Y(n_3005)
);

CKINVDCx6p67_ASAP7_75t_R g3006 ( 
.A(n_2406),
.Y(n_3006)
);

BUFx2_ASAP7_75t_L g3007 ( 
.A(n_2617),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2517),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_L g3009 ( 
.A(n_2489),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2519),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2358),
.B(n_2247),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2644),
.B(n_2309),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2521),
.Y(n_3013)
);

NAND3xp33_ASAP7_75t_L g3014 ( 
.A(n_2667),
.B(n_2307),
.C(n_2304),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2341),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2370),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2522),
.Y(n_3017)
);

INVx2_ASAP7_75t_SL g3018 ( 
.A(n_2757),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2370),
.Y(n_3019)
);

AND2x4_ASAP7_75t_SL g3020 ( 
.A(n_2634),
.B(n_2142),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2532),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2704),
.B(n_2309),
.Y(n_3022)
);

INVx5_ASAP7_75t_L g3023 ( 
.A(n_2735),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_SL g3024 ( 
.A(n_2596),
.B(n_2310),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2714),
.B(n_2310),
.Y(n_3025)
);

INVx3_ASAP7_75t_L g3026 ( 
.A(n_2489),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2730),
.B(n_2122),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_SL g3028 ( 
.A(n_2598),
.B(n_2247),
.Y(n_3028)
);

INVx3_ASAP7_75t_L g3029 ( 
.A(n_2489),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2370),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2737),
.B(n_2754),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_2397),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2705),
.B(n_2178),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2534),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2409),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_2598),
.B(n_2248),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_SL g3037 ( 
.A(n_2627),
.B(n_2248),
.Y(n_3037)
);

OAI22xp33_ASAP7_75t_L g3038 ( 
.A1(n_2751),
.A2(n_2091),
.B1(n_2266),
.B2(n_2249),
.Y(n_3038)
);

INVx2_ASAP7_75t_SL g3039 ( 
.A(n_2757),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2629),
.B(n_2249),
.Y(n_3040)
);

INVx2_ASAP7_75t_L g3041 ( 
.A(n_2409),
.Y(n_3041)
);

BUFx2_ASAP7_75t_L g3042 ( 
.A(n_2589),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2409),
.Y(n_3043)
);

BUFx6f_ASAP7_75t_L g3044 ( 
.A(n_2493),
.Y(n_3044)
);

NOR2xp33_ASAP7_75t_L g3045 ( 
.A(n_2362),
.B(n_2304),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2428),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2428),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2707),
.B(n_2178),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2428),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2674),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2709),
.B(n_2208),
.Y(n_3051)
);

INVx3_ASAP7_75t_L g3052 ( 
.A(n_2493),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2676),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2493),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2677),
.Y(n_3055)
);

BUFx6f_ASAP7_75t_SL g3056 ( 
.A(n_2334),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2718),
.B(n_2208),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2536),
.Y(n_3058)
);

CKINVDCx6p67_ASAP7_75t_R g3059 ( 
.A(n_2406),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2512),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2355),
.Y(n_3061)
);

INVx3_ASAP7_75t_L g3062 ( 
.A(n_2493),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2563),
.B(n_2322),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2537),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_SL g3065 ( 
.A(n_2575),
.B(n_2322),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2683),
.Y(n_3066)
);

INVx2_ASAP7_75t_SL g3067 ( 
.A(n_2600),
.Y(n_3067)
);

INVx2_ASAP7_75t_L g3068 ( 
.A(n_2685),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2728),
.B(n_2313),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2691),
.Y(n_3070)
);

BUFx6f_ASAP7_75t_L g3071 ( 
.A(n_2495),
.Y(n_3071)
);

INVx2_ASAP7_75t_L g3072 ( 
.A(n_2692),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2544),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2693),
.Y(n_3074)
);

INVx3_ASAP7_75t_L g3075 ( 
.A(n_2495),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2547),
.Y(n_3076)
);

INVx2_ASAP7_75t_SL g3077 ( 
.A(n_2464),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2552),
.Y(n_3078)
);

INVx4_ASAP7_75t_L g3079 ( 
.A(n_2735),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2731),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2560),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_SL g3082 ( 
.A(n_2673),
.B(n_2276),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2561),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2565),
.B(n_2225),
.Y(n_3084)
);

NAND3xp33_ASAP7_75t_L g3085 ( 
.A(n_2338),
.B(n_2324),
.C(n_2276),
.Y(n_3085)
);

OR2x2_ASAP7_75t_L g3086 ( 
.A(n_2711),
.B(n_2272),
.Y(n_3086)
);

BUFx6f_ASAP7_75t_L g3087 ( 
.A(n_2495),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2741),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2745),
.Y(n_3089)
);

INVx1_ASAP7_75t_SL g3090 ( 
.A(n_2755),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2570),
.Y(n_3091)
);

BUFx3_ASAP7_75t_L g3092 ( 
.A(n_2355),
.Y(n_3092)
);

AOI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2684),
.A2(n_2327),
.B1(n_2181),
.B2(n_2195),
.Y(n_3093)
);

NAND2xp33_ASAP7_75t_SL g3094 ( 
.A(n_2440),
.B(n_2142),
.Y(n_3094)
);

INVx4_ASAP7_75t_L g3095 ( 
.A(n_2735),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2495),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2750),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2571),
.Y(n_3098)
);

BUFx6f_ASAP7_75t_L g3099 ( 
.A(n_2574),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2572),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2576),
.Y(n_3101)
);

OAI22xp5_ASAP7_75t_L g3102 ( 
.A1(n_2436),
.A2(n_2045),
.B1(n_2324),
.B2(n_2225),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2756),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2581),
.Y(n_3104)
);

INVx4_ASAP7_75t_L g3105 ( 
.A(n_2735),
.Y(n_3105)
);

INVx2_ASAP7_75t_L g3106 ( 
.A(n_2365),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2583),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_2498),
.B(n_2502),
.Y(n_3108)
);

INVx1_ASAP7_75t_SL g3109 ( 
.A(n_2468),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2367),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2585),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2586),
.Y(n_3112)
);

INVx5_ASAP7_75t_L g3113 ( 
.A(n_2574),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2381),
.B(n_1970),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2371),
.B(n_1670),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2359),
.Y(n_3116)
);

NAND2xp33_ASAP7_75t_L g3117 ( 
.A(n_2660),
.B(n_1952),
.Y(n_3117)
);

NOR2x1p5_ASAP7_75t_L g3118 ( 
.A(n_2503),
.B(n_2331),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2574),
.Y(n_3119)
);

NOR3xp33_ASAP7_75t_L g3120 ( 
.A(n_2509),
.B(n_2238),
.C(n_2069),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_SL g3121 ( 
.A(n_2642),
.B(n_2211),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_SL g3122 ( 
.A(n_2699),
.B(n_2211),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_SL g3123 ( 
.A(n_2702),
.B(n_2211),
.Y(n_3123)
);

BUFx2_ASAP7_75t_L g3124 ( 
.A(n_2712),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2359),
.Y(n_3125)
);

INVx2_ASAP7_75t_L g3126 ( 
.A(n_2359),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2587),
.B(n_2225),
.Y(n_3127)
);

INVx4_ASAP7_75t_L g3128 ( 
.A(n_2574),
.Y(n_3128)
);

INVx2_ASAP7_75t_SL g3129 ( 
.A(n_2376),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2588),
.B(n_2225),
.Y(n_3130)
);

INVx2_ASAP7_75t_SL g3131 ( 
.A(n_2376),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_2578),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2593),
.B(n_1970),
.Y(n_3133)
);

INVx5_ASAP7_75t_L g3134 ( 
.A(n_2578),
.Y(n_3134)
);

NOR2xp33_ASAP7_75t_L g3135 ( 
.A(n_2371),
.B(n_1670),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2597),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_2355),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2609),
.Y(n_3138)
);

AOI22xp5_ASAP7_75t_L g3139 ( 
.A1(n_2614),
.A2(n_2073),
.B1(n_2123),
.B2(n_2054),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2375),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2619),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2623),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2375),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_SL g3144 ( 
.A(n_2720),
.B(n_2211),
.Y(n_3144)
);

BUFx6f_ASAP7_75t_SL g3145 ( 
.A(n_2334),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_SL g3146 ( 
.A(n_2539),
.B(n_2303),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_SL g3147 ( 
.A(n_2539),
.B(n_2303),
.Y(n_3147)
);

INVxp67_ASAP7_75t_SL g3148 ( 
.A(n_2335),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2630),
.B(n_1969),
.Y(n_3149)
);

NAND3xp33_ASAP7_75t_L g3150 ( 
.A(n_2338),
.B(n_2454),
.C(n_2437),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2632),
.B(n_2162),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2633),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_SL g3153 ( 
.A(n_2539),
.B(n_2303),
.Y(n_3153)
);

CKINVDCx5p33_ASAP7_75t_R g3154 ( 
.A(n_2379),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_SL g3155 ( 
.A(n_2613),
.B(n_2303),
.Y(n_3155)
);

INVx3_ASAP7_75t_L g3156 ( 
.A(n_2578),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_2645),
.A2(n_2073),
.B1(n_2123),
.B2(n_2054),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_2388),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2652),
.B(n_2162),
.Y(n_3159)
);

INVx2_ASAP7_75t_L g3160 ( 
.A(n_2392),
.Y(n_3160)
);

AO21x2_ASAP7_75t_L g3161 ( 
.A1(n_2392),
.A2(n_2501),
.B(n_2400),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2654),
.Y(n_3162)
);

CKINVDCx6p67_ASAP7_75t_R g3163 ( 
.A(n_2420),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2400),
.Y(n_3164)
);

INVx2_ASAP7_75t_SL g3165 ( 
.A(n_2376),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2501),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2663),
.B(n_2550),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2514),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2550),
.B(n_2162),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2514),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2518),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2518),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_SL g3173 ( 
.A(n_2678),
.B(n_2098),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_2457),
.B(n_2047),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2472),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2478),
.Y(n_3176)
);

INVx1_ASAP7_75t_L g3177 ( 
.A(n_2478),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_2650),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2650),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2550),
.B(n_2229),
.Y(n_3180)
);

INVx2_ASAP7_75t_L g3181 ( 
.A(n_2650),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2725),
.B(n_2380),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2490),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2499),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2499),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2608),
.Y(n_3186)
);

INVx1_ASAP7_75t_L g3187 ( 
.A(n_2608),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2608),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2615),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2615),
.Y(n_3190)
);

NOR2xp33_ASAP7_75t_L g3191 ( 
.A(n_2379),
.B(n_1676),
.Y(n_3191)
);

NOR2xp33_ASAP7_75t_L g3192 ( 
.A(n_2383),
.B(n_2396),
.Y(n_3192)
);

INVx2_ASAP7_75t_L g3193 ( 
.A(n_2615),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_2646),
.B(n_2229),
.Y(n_3194)
);

BUFx10_ASAP7_75t_L g3195 ( 
.A(n_2555),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2656),
.Y(n_3196)
);

NOR2xp33_ASAP7_75t_L g3197 ( 
.A(n_2383),
.B(n_1676),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_SL g3198 ( 
.A(n_2528),
.B(n_2098),
.Y(n_3198)
);

CKINVDCx6p67_ASAP7_75t_R g3199 ( 
.A(n_2420),
.Y(n_3199)
);

NAND3xp33_ASAP7_75t_L g3200 ( 
.A(n_2742),
.B(n_2261),
.C(n_1944),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_2657),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2657),
.Y(n_3202)
);

CKINVDCx5p33_ASAP7_75t_R g3203 ( 
.A(n_2396),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2670),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2670),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2380),
.B(n_2229),
.Y(n_3206)
);

NOR2x1p5_ASAP7_75t_L g3207 ( 
.A(n_2503),
.B(n_2285),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_SL g3208 ( 
.A(n_2506),
.B(n_2274),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_2670),
.Y(n_3209)
);

AND2x2_ASAP7_75t_SL g3210 ( 
.A(n_2943),
.B(n_2853),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2867),
.B(n_2407),
.Y(n_3211)
);

INVx2_ASAP7_75t_SL g3212 ( 
.A(n_3118),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2766),
.B(n_2116),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2811),
.B(n_2116),
.Y(n_3214)
);

CKINVDCx5p33_ASAP7_75t_R g3215 ( 
.A(n_2936),
.Y(n_3215)
);

NAND2xp33_ASAP7_75t_L g3216 ( 
.A(n_2804),
.B(n_2407),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3149),
.B(n_2116),
.Y(n_3217)
);

OR2x6_ASAP7_75t_L g3218 ( 
.A(n_2873),
.B(n_2905),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2828),
.B(n_2132),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_2913),
.B(n_2612),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2824),
.B(n_2132),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2913),
.B(n_2621),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2793),
.B(n_2132),
.Y(n_3223)
);

AND2x4_ASAP7_75t_L g3224 ( 
.A(n_3118),
.B(n_2679),
.Y(n_3224)
);

CKINVDCx5p33_ASAP7_75t_R g3225 ( 
.A(n_2928),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2791),
.B(n_2135),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2993),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2768),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_2791),
.B(n_2908),
.Y(n_3229)
);

INVx4_ASAP7_75t_L g3230 ( 
.A(n_3113),
.Y(n_3230)
);

OR2x2_ASAP7_75t_L g3231 ( 
.A(n_2834),
.B(n_2411),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3031),
.B(n_2135),
.Y(n_3232)
);

AOI22xp33_ASAP7_75t_L g3233 ( 
.A1(n_2876),
.A2(n_2453),
.B1(n_2716),
.B2(n_2708),
.Y(n_3233)
);

BUFx6f_ASAP7_75t_L g3234 ( 
.A(n_2840),
.Y(n_3234)
);

BUFx3_ASAP7_75t_L g3235 ( 
.A(n_2782),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2787),
.Y(n_3236)
);

AND2x2_ASAP7_75t_L g3237 ( 
.A(n_3108),
.B(n_2411),
.Y(n_3237)
);

NAND2xp33_ASAP7_75t_L g3238 ( 
.A(n_2804),
.B(n_2529),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2774),
.Y(n_3239)
);

NOR2xp33_ASAP7_75t_L g3240 ( 
.A(n_2770),
.B(n_2592),
.Y(n_3240)
);

AND2x6_ASAP7_75t_L g3241 ( 
.A(n_2963),
.B(n_2380),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3108),
.B(n_2582),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2774),
.Y(n_3243)
);

NOR2xp33_ASAP7_75t_L g3244 ( 
.A(n_2770),
.B(n_2494),
.Y(n_3244)
);

BUFx4f_ASAP7_75t_L g3245 ( 
.A(n_2899),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_3174),
.B(n_2513),
.Y(n_3246)
);

AND2x2_ASAP7_75t_L g3247 ( 
.A(n_3174),
.B(n_2541),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2778),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_3194),
.B(n_2681),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2780),
.B(n_2135),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2780),
.B(n_2783),
.Y(n_3251)
);

BUFx10_ASAP7_75t_L g3252 ( 
.A(n_3115),
.Y(n_3252)
);

AND2x6_ASAP7_75t_L g3253 ( 
.A(n_2963),
.B(n_2902),
.Y(n_3253)
);

INVx3_ASAP7_75t_L g3254 ( 
.A(n_2767),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3114),
.B(n_2557),
.Y(n_3255)
);

CKINVDCx20_ASAP7_75t_R g3256 ( 
.A(n_2899),
.Y(n_3256)
);

INVx4_ASAP7_75t_L g3257 ( 
.A(n_3113),
.Y(n_3257)
);

INVx3_ASAP7_75t_L g3258 ( 
.A(n_2767),
.Y(n_3258)
);

AND2x6_ASAP7_75t_L g3259 ( 
.A(n_2902),
.B(n_2418),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2860),
.B(n_1683),
.Y(n_3260)
);

AND2x4_ASAP7_75t_L g3261 ( 
.A(n_3194),
.B(n_2717),
.Y(n_3261)
);

BUFx3_ASAP7_75t_L g3262 ( 
.A(n_3007),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2784),
.Y(n_3263)
);

BUFx6f_ASAP7_75t_L g3264 ( 
.A(n_2840),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_2784),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_2796),
.Y(n_3266)
);

CKINVDCx5p33_ASAP7_75t_R g3267 ( 
.A(n_2928),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2796),
.Y(n_3268)
);

HB1xp67_ASAP7_75t_L g3269 ( 
.A(n_3007),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2799),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2799),
.B(n_2066),
.Y(n_3271)
);

INVxp67_ASAP7_75t_SL g3272 ( 
.A(n_2852),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_L g3273 ( 
.A(n_2803),
.B(n_2156),
.Y(n_3273)
);

BUFx2_ASAP7_75t_L g3274 ( 
.A(n_2951),
.Y(n_3274)
);

INVxp67_ASAP7_75t_SL g3275 ( 
.A(n_2858),
.Y(n_3275)
);

BUFx2_ASAP7_75t_L g3276 ( 
.A(n_2951),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2789),
.Y(n_3277)
);

BUFx6f_ASAP7_75t_L g3278 ( 
.A(n_2840),
.Y(n_3278)
);

BUFx6f_ASAP7_75t_L g3279 ( 
.A(n_2840),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2803),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2812),
.B(n_2156),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_2834),
.B(n_2591),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2812),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2813),
.B(n_2156),
.Y(n_3284)
);

AND2x6_ASAP7_75t_L g3285 ( 
.A(n_3139),
.B(n_2418),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_3194),
.B(n_3129),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2790),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_2790),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_2792),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_3114),
.B(n_2274),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_2813),
.Y(n_3291)
);

OR2x2_ASAP7_75t_L g3292 ( 
.A(n_3000),
.B(n_2602),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2827),
.Y(n_3293)
);

BUFx6f_ASAP7_75t_L g3294 ( 
.A(n_2840),
.Y(n_3294)
);

BUFx6f_ASAP7_75t_L g3295 ( 
.A(n_2855),
.Y(n_3295)
);

AOI22xp33_ASAP7_75t_L g3296 ( 
.A1(n_2764),
.A2(n_2708),
.B1(n_2203),
.B2(n_2643),
.Y(n_3296)
);

NAND2x1p5_ASAP7_75t_L g3297 ( 
.A(n_2943),
.B(n_2355),
.Y(n_3297)
);

BUFx4f_ASAP7_75t_L g3298 ( 
.A(n_3006),
.Y(n_3298)
);

BUFx6f_ASAP7_75t_SL g3299 ( 
.A(n_2884),
.Y(n_3299)
);

AND2x6_ASAP7_75t_L g3300 ( 
.A(n_3139),
.B(n_2418),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2827),
.Y(n_3301)
);

AND2x4_ASAP7_75t_L g3302 ( 
.A(n_3194),
.B(n_2740),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_2878),
.B(n_2688),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_2767),
.Y(n_3304)
);

BUFx3_ASAP7_75t_L g3305 ( 
.A(n_2805),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2839),
.B(n_2045),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_3129),
.B(n_2688),
.Y(n_3307)
);

INVx3_ASAP7_75t_L g3308 ( 
.A(n_2775),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_2839),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_2844),
.Y(n_3310)
);

AND2x6_ASAP7_75t_L g3311 ( 
.A(n_3157),
.B(n_2785),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_2792),
.Y(n_3312)
);

AO22x2_ASAP7_75t_L g3313 ( 
.A1(n_3150),
.A2(n_2326),
.B1(n_2391),
.B2(n_2182),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_2794),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_2772),
.Y(n_3315)
);

INVx1_ASAP7_75t_SL g3316 ( 
.A(n_2772),
.Y(n_3316)
);

INVx3_ASAP7_75t_L g3317 ( 
.A(n_2775),
.Y(n_3317)
);

INVx2_ASAP7_75t_L g3318 ( 
.A(n_2794),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2801),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_2846),
.B(n_2848),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2846),
.B(n_2045),
.Y(n_3321)
);

AND2x4_ASAP7_75t_L g3322 ( 
.A(n_3131),
.B(n_2423),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2848),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_2801),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2859),
.B(n_2334),
.Y(n_3325)
);

AND2x6_ASAP7_75t_L g3326 ( 
.A(n_3157),
.B(n_2423),
.Y(n_3326)
);

BUFx4f_ASAP7_75t_L g3327 ( 
.A(n_3006),
.Y(n_3327)
);

NOR2xp33_ASAP7_75t_L g3328 ( 
.A(n_2931),
.B(n_1715),
.Y(n_3328)
);

NOR2xp33_ASAP7_75t_L g3329 ( 
.A(n_2938),
.B(n_1716),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2865),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2865),
.Y(n_3331)
);

INVx1_ASAP7_75t_SL g3332 ( 
.A(n_2773),
.Y(n_3332)
);

NAND2x1p5_ASAP7_75t_L g3333 ( 
.A(n_2943),
.B(n_2372),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2877),
.B(n_2334),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2877),
.Y(n_3335)
);

AND2x6_ASAP7_75t_L g3336 ( 
.A(n_2785),
.B(n_2775),
.Y(n_3336)
);

INVx5_ASAP7_75t_L g3337 ( 
.A(n_2873),
.Y(n_3337)
);

CKINVDCx5p33_ASAP7_75t_R g3338 ( 
.A(n_3059),
.Y(n_3338)
);

INVx4_ASAP7_75t_SL g3339 ( 
.A(n_2923),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_2958),
.B(n_1716),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3011),
.B(n_2278),
.Y(n_3341)
);

INVx2_ASAP7_75t_SL g3342 ( 
.A(n_2884),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2892),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2892),
.Y(n_3344)
);

NAND2x1p5_ASAP7_75t_L g3345 ( 
.A(n_2795),
.B(n_2372),
.Y(n_3345)
);

INVx1_ASAP7_75t_SL g3346 ( 
.A(n_2773),
.Y(n_3346)
);

INVx1_ASAP7_75t_SL g3347 ( 
.A(n_2829),
.Y(n_3347)
);

INVx2_ASAP7_75t_L g3348 ( 
.A(n_2802),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2893),
.B(n_2894),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2893),
.Y(n_3350)
);

AND2x4_ASAP7_75t_L g3351 ( 
.A(n_3131),
.B(n_2423),
.Y(n_3351)
);

BUFx2_ASAP7_75t_L g3352 ( 
.A(n_2805),
.Y(n_3352)
);

INVx5_ASAP7_75t_L g3353 ( 
.A(n_2873),
.Y(n_3353)
);

NOR2xp33_ASAP7_75t_L g3354 ( 
.A(n_3045),
.B(n_1717),
.Y(n_3354)
);

OR2x2_ASAP7_75t_L g3355 ( 
.A(n_3086),
.B(n_2278),
.Y(n_3355)
);

INVx3_ASAP7_75t_L g3356 ( 
.A(n_2836),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_2894),
.Y(n_3357)
);

INVx2_ASAP7_75t_L g3358 ( 
.A(n_2802),
.Y(n_3358)
);

BUFx2_ASAP7_75t_L g3359 ( 
.A(n_2887),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2815),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_2896),
.Y(n_3361)
);

INVx3_ASAP7_75t_L g3362 ( 
.A(n_2836),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_2896),
.B(n_2296),
.Y(n_3363)
);

INVx1_ASAP7_75t_SL g3364 ( 
.A(n_2829),
.Y(n_3364)
);

BUFx10_ASAP7_75t_L g3365 ( 
.A(n_3135),
.Y(n_3365)
);

BUFx2_ASAP7_75t_L g3366 ( 
.A(n_2887),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2909),
.Y(n_3367)
);

INVx3_ASAP7_75t_L g3368 ( 
.A(n_2836),
.Y(n_3368)
);

INVx1_ASAP7_75t_L g3369 ( 
.A(n_2909),
.Y(n_3369)
);

OR2x2_ASAP7_75t_L g3370 ( 
.A(n_3086),
.B(n_2285),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_2917),
.Y(n_3371)
);

AND2x6_ASAP7_75t_L g3372 ( 
.A(n_2785),
.B(n_2433),
.Y(n_3372)
);

HB1xp67_ASAP7_75t_L g3373 ( 
.A(n_2835),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2917),
.Y(n_3374)
);

BUFx6f_ASAP7_75t_L g3375 ( 
.A(n_2855),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2920),
.Y(n_3376)
);

AND2x2_ASAP7_75t_L g3377 ( 
.A(n_2948),
.B(n_2287),
.Y(n_3377)
);

BUFx6f_ASAP7_75t_L g3378 ( 
.A(n_2855),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2815),
.Y(n_3379)
);

INVx3_ASAP7_75t_L g3380 ( 
.A(n_2849),
.Y(n_3380)
);

AND2x6_ASAP7_75t_L g3381 ( 
.A(n_2785),
.B(n_2433),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2925),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_2816),
.Y(n_3383)
);

INVxp67_ASAP7_75t_L g3384 ( 
.A(n_3148),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2925),
.B(n_2296),
.Y(n_3385)
);

BUFx3_ASAP7_75t_L g3386 ( 
.A(n_3163),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2816),
.Y(n_3387)
);

INVx4_ASAP7_75t_L g3388 ( 
.A(n_3113),
.Y(n_3388)
);

AND2x4_ASAP7_75t_L g3389 ( 
.A(n_3165),
.B(n_2433),
.Y(n_3389)
);

OAI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3038),
.A2(n_2480),
.B1(n_2033),
.B2(n_2641),
.Y(n_3390)
);

INVx1_ASAP7_75t_SL g3391 ( 
.A(n_3090),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2929),
.Y(n_3392)
);

BUFx6f_ASAP7_75t_L g3393 ( 
.A(n_2855),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2929),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_3163),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_2948),
.B(n_2288),
.Y(n_3396)
);

INVx1_ASAP7_75t_SL g3397 ( 
.A(n_3090),
.Y(n_3397)
);

NAND2xp5_ASAP7_75t_L g3398 ( 
.A(n_2937),
.B(n_2296),
.Y(n_3398)
);

INVx2_ASAP7_75t_L g3399 ( 
.A(n_2818),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2937),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2940),
.B(n_2296),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3192),
.B(n_2288),
.Y(n_3402)
);

OR2x2_ASAP7_75t_L g3403 ( 
.A(n_2962),
.B(n_2298),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_2940),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_2946),
.B(n_2315),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_2946),
.Y(n_3406)
);

INVx3_ASAP7_75t_L g3407 ( 
.A(n_2849),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_2954),
.B(n_2315),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_2818),
.Y(n_3409)
);

INVx4_ASAP7_75t_L g3410 ( 
.A(n_3113),
.Y(n_3410)
);

BUFx6f_ASAP7_75t_L g3411 ( 
.A(n_2855),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2954),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2959),
.Y(n_3413)
);

BUFx3_ASAP7_75t_L g3414 ( 
.A(n_3199),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2959),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_2820),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_L g3417 ( 
.A(n_2843),
.B(n_1751),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_2968),
.B(n_2315),
.Y(n_3418)
);

OR2x2_ASAP7_75t_L g3419 ( 
.A(n_2962),
.B(n_2298),
.Y(n_3419)
);

INVx5_ASAP7_75t_L g3420 ( 
.A(n_2873),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2968),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_2970),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_2970),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_2880),
.B(n_2302),
.Y(n_3424)
);

BUFx4f_ASAP7_75t_L g3425 ( 
.A(n_3199),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2820),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_2977),
.B(n_2315),
.Y(n_3427)
);

INVxp33_ASAP7_75t_L g3428 ( 
.A(n_3191),
.Y(n_3428)
);

AO22x2_ASAP7_75t_L g3429 ( 
.A1(n_3150),
.A2(n_2326),
.B1(n_2182),
.B2(n_1958),
.Y(n_3429)
);

BUFx6f_ASAP7_75t_L g3430 ( 
.A(n_2978),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2977),
.B(n_2164),
.Y(n_3431)
);

OR2x6_ASAP7_75t_L g3432 ( 
.A(n_2873),
.B(n_2554),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_2822),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_2822),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2985),
.Y(n_3435)
);

INVx3_ASAP7_75t_L g3436 ( 
.A(n_2849),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_3197),
.B(n_1754),
.Y(n_3437)
);

OR2x6_ASAP7_75t_L g3438 ( 
.A(n_2905),
.B(n_2444),
.Y(n_3438)
);

AND2x4_ASAP7_75t_L g3439 ( 
.A(n_3165),
.B(n_2444),
.Y(n_3439)
);

BUFx2_ASAP7_75t_L g3440 ( 
.A(n_2945),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_2825),
.Y(n_3441)
);

AND2x4_ASAP7_75t_L g3442 ( 
.A(n_3067),
.B(n_2444),
.Y(n_3442)
);

INVx3_ASAP7_75t_L g3443 ( 
.A(n_3060),
.Y(n_3443)
);

INVx3_ASAP7_75t_L g3444 ( 
.A(n_3060),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_2825),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_2851),
.B(n_2955),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2985),
.B(n_2164),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3109),
.B(n_2260),
.Y(n_3448)
);

OR2x2_ASAP7_75t_L g3449 ( 
.A(n_2851),
.B(n_2326),
.Y(n_3449)
);

CKINVDCx5p33_ASAP7_75t_R g3450 ( 
.A(n_3154),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_2992),
.B(n_2164),
.Y(n_3451)
);

INVx3_ASAP7_75t_L g3452 ( 
.A(n_3128),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2992),
.B(n_2164),
.Y(n_3453)
);

CKINVDCx5p33_ASAP7_75t_R g3454 ( 
.A(n_3154),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3203),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_2826),
.Y(n_3456)
);

AND3x4_ASAP7_75t_L g3457 ( 
.A(n_3120),
.B(n_2326),
.C(n_2260),
.Y(n_3457)
);

HB1xp67_ASAP7_75t_L g3458 ( 
.A(n_2817),
.Y(n_3458)
);

AO21x2_ASAP7_75t_L g3459 ( 
.A1(n_2850),
.A2(n_2527),
.B(n_2456),
.Y(n_3459)
);

HB1xp67_ASAP7_75t_L g3460 ( 
.A(n_3169),
.Y(n_3460)
);

AND2x4_ASAP7_75t_L g3461 ( 
.A(n_3067),
.B(n_2486),
.Y(n_3461)
);

INVx5_ASAP7_75t_L g3462 ( 
.A(n_2905),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_2995),
.B(n_2164),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_3109),
.B(n_2260),
.Y(n_3464)
);

BUFx10_ASAP7_75t_L g3465 ( 
.A(n_3203),
.Y(n_3465)
);

AND2x6_ASAP7_75t_L g3466 ( 
.A(n_3061),
.B(n_2486),
.Y(n_3466)
);

INVxp67_ASAP7_75t_SL g3467 ( 
.A(n_2864),
.Y(n_3467)
);

INVx4_ASAP7_75t_L g3468 ( 
.A(n_3134),
.Y(n_3468)
);

AND2x6_ASAP7_75t_L g3469 ( 
.A(n_3061),
.B(n_2486),
.Y(n_3469)
);

AOI22xp33_ASAP7_75t_L g3470 ( 
.A1(n_2923),
.A2(n_2203),
.B1(n_2643),
.B2(n_2641),
.Y(n_3470)
);

NOR3xp33_ASAP7_75t_L g3471 ( 
.A(n_3014),
.B(n_2250),
.C(n_2080),
.Y(n_3471)
);

INVx4_ASAP7_75t_L g3472 ( 
.A(n_3134),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_2995),
.B(n_2997),
.Y(n_3473)
);

XNOR2x2_ASAP7_75t_L g3474 ( 
.A(n_2984),
.B(n_2262),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_2826),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_2997),
.Y(n_3476)
);

NAND2x1p5_ASAP7_75t_L g3477 ( 
.A(n_2795),
.B(n_2372),
.Y(n_3477)
);

AND2x2_ASAP7_75t_SL g3478 ( 
.A(n_2853),
.B(n_2530),
.Y(n_3478)
);

NOR2xp33_ASAP7_75t_L g3479 ( 
.A(n_2921),
.B(n_1754),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_2830),
.Y(n_3480)
);

AND2x4_ASAP7_75t_L g3481 ( 
.A(n_3207),
.B(n_3020),
.Y(n_3481)
);

NOR2xp33_ASAP7_75t_L g3482 ( 
.A(n_2933),
.B(n_1769),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3001),
.Y(n_3483)
);

AOI22xp33_ASAP7_75t_L g3484 ( 
.A1(n_2923),
.A2(n_2095),
.B1(n_2463),
.B2(n_2441),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3008),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_SL g3486 ( 
.A(n_3077),
.B(n_2399),
.Y(n_3486)
);

CKINVDCx20_ASAP7_75t_R g3487 ( 
.A(n_2944),
.Y(n_3487)
);

BUFx10_ASAP7_75t_L g3488 ( 
.A(n_2944),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3008),
.Y(n_3489)
);

NAND2xp33_ASAP7_75t_L g3490 ( 
.A(n_2804),
.B(n_2538),
.Y(n_3490)
);

INVx2_ASAP7_75t_SL g3491 ( 
.A(n_2884),
.Y(n_3491)
);

AND2x2_ASAP7_75t_L g3492 ( 
.A(n_3077),
.B(n_2260),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_2830),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_L g3494 ( 
.A(n_3010),
.B(n_2165),
.Y(n_3494)
);

OAI22xp5_ASAP7_75t_L g3495 ( 
.A1(n_3133),
.A2(n_3013),
.B1(n_3017),
.B2(n_3010),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3013),
.Y(n_3496)
);

INVx4_ASAP7_75t_L g3497 ( 
.A(n_3134),
.Y(n_3497)
);

INVx3_ASAP7_75t_L g3498 ( 
.A(n_3128),
.Y(n_3498)
);

INVx4_ASAP7_75t_L g3499 ( 
.A(n_3134),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_3017),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_3021),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3021),
.B(n_2165),
.Y(n_3502)
);

BUFx6f_ASAP7_75t_L g3503 ( 
.A(n_2978),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3128),
.Y(n_3504)
);

INVx3_ASAP7_75t_L g3505 ( 
.A(n_3128),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3034),
.B(n_2165),
.Y(n_3506)
);

INVx4_ASAP7_75t_L g3507 ( 
.A(n_3134),
.Y(n_3507)
);

BUFx10_ASAP7_75t_L g3508 ( 
.A(n_3032),
.Y(n_3508)
);

INVx4_ASAP7_75t_L g3509 ( 
.A(n_2814),
.Y(n_3509)
);

INVx3_ASAP7_75t_L g3510 ( 
.A(n_3061),
.Y(n_3510)
);

AND2x4_ASAP7_75t_L g3511 ( 
.A(n_3207),
.B(n_2530),
.Y(n_3511)
);

BUFx3_ASAP7_75t_L g3512 ( 
.A(n_3042),
.Y(n_3512)
);

INVx2_ASAP7_75t_SL g3513 ( 
.A(n_3195),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3058),
.B(n_2165),
.Y(n_3514)
);

NAND2x1p5_ASAP7_75t_L g3515 ( 
.A(n_2795),
.B(n_2372),
.Y(n_3515)
);

BUFx4f_ASAP7_75t_L g3516 ( 
.A(n_3124),
.Y(n_3516)
);

BUFx2_ASAP7_75t_L g3517 ( 
.A(n_3124),
.Y(n_3517)
);

OR2x6_ASAP7_75t_L g3518 ( 
.A(n_2905),
.B(n_2530),
.Y(n_3518)
);

INVx4_ASAP7_75t_L g3519 ( 
.A(n_2814),
.Y(n_3519)
);

AOI22xp33_ASAP7_75t_L g3520 ( 
.A1(n_3093),
.A2(n_2631),
.B1(n_2628),
.B2(n_2569),
.Y(n_3520)
);

NOR2xp67_ASAP7_75t_L g3521 ( 
.A(n_2845),
.B(n_2556),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3058),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_2807),
.B(n_3033),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3064),
.Y(n_3524)
);

AO22x2_ASAP7_75t_L g3525 ( 
.A1(n_2845),
.A2(n_2107),
.B1(n_2181),
.B2(n_2160),
.Y(n_3525)
);

OAI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3064),
.A2(n_2033),
.B1(n_2169),
.B2(n_2168),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3073),
.Y(n_3527)
);

BUFx6f_ASAP7_75t_L g3528 ( 
.A(n_2978),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3073),
.B(n_2165),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3076),
.Y(n_3530)
);

OR2x2_ASAP7_75t_L g3531 ( 
.A(n_3048),
.B(n_2558),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3076),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_2832),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_L g3534 ( 
.A(n_2881),
.B(n_1769),
.Y(n_3534)
);

CKINVDCx5p33_ASAP7_75t_R g3535 ( 
.A(n_3032),
.Y(n_3535)
);

INVx5_ASAP7_75t_L g3536 ( 
.A(n_2905),
.Y(n_3536)
);

INVx2_ASAP7_75t_SL g3537 ( 
.A(n_3195),
.Y(n_3537)
);

INVx3_ASAP7_75t_L g3538 ( 
.A(n_3092),
.Y(n_3538)
);

AOI22xp33_ASAP7_75t_L g3539 ( 
.A1(n_2932),
.A2(n_2095),
.B1(n_2181),
.B2(n_2160),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_3078),
.B(n_2171),
.Y(n_3540)
);

AND2x2_ASAP7_75t_L g3541 ( 
.A(n_2807),
.B(n_3051),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_3081),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3027),
.B(n_1787),
.Y(n_3543)
);

AND2x4_ASAP7_75t_L g3544 ( 
.A(n_3020),
.B(n_2448),
.Y(n_3544)
);

INVx4_ASAP7_75t_L g3545 ( 
.A(n_2890),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3081),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_SL g3547 ( 
.A(n_2795),
.B(n_2603),
.Y(n_3547)
);

INVx5_ASAP7_75t_L g3548 ( 
.A(n_2934),
.Y(n_3548)
);

INVx2_ASAP7_75t_L g3549 ( 
.A(n_2832),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_2833),
.Y(n_3550)
);

AND2x6_ASAP7_75t_L g3551 ( 
.A(n_3092),
.B(n_2680),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3083),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3083),
.Y(n_3553)
);

AND2x2_ASAP7_75t_L g3554 ( 
.A(n_3057),
.B(n_2128),
.Y(n_3554)
);

AND2x4_ASAP7_75t_L g3555 ( 
.A(n_3020),
.B(n_3146),
.Y(n_3555)
);

INVx1_ASAP7_75t_SL g3556 ( 
.A(n_2800),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_2833),
.Y(n_3557)
);

AND2x4_ASAP7_75t_L g3558 ( 
.A(n_3147),
.B(n_2491),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3091),
.B(n_2171),
.Y(n_3559)
);

AOI22xp33_ASAP7_75t_L g3560 ( 
.A1(n_2932),
.A2(n_2181),
.B1(n_2195),
.B2(n_2160),
.Y(n_3560)
);

AND2x4_ASAP7_75t_L g3561 ( 
.A(n_3153),
.B(n_2616),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3091),
.B(n_2171),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_2853),
.B(n_2128),
.Y(n_3563)
);

NOR2xp33_ASAP7_75t_L g3564 ( 
.A(n_2883),
.B(n_1793),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3098),
.Y(n_3565)
);

CKINVDCx5p33_ASAP7_75t_R g3566 ( 
.A(n_3195),
.Y(n_3566)
);

BUFx6f_ASAP7_75t_L g3567 ( 
.A(n_2978),
.Y(n_3567)
);

BUFx6f_ASAP7_75t_L g3568 ( 
.A(n_2978),
.Y(n_3568)
);

AO22x1_ASAP7_75t_L g3569 ( 
.A1(n_2806),
.A2(n_2607),
.B1(n_2618),
.B2(n_2604),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_2837),
.Y(n_3570)
);

OR2x6_ASAP7_75t_L g3571 ( 
.A(n_2934),
.B(n_2640),
.Y(n_3571)
);

INVxp67_ASAP7_75t_L g3572 ( 
.A(n_3282),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3315),
.B(n_3069),
.Y(n_3573)
);

NOR2xp33_ASAP7_75t_L g3574 ( 
.A(n_3428),
.B(n_2429),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_SL g3575 ( 
.A(n_3347),
.B(n_2809),
.Y(n_3575)
);

BUFx3_ASAP7_75t_L g3576 ( 
.A(n_3274),
.Y(n_3576)
);

AOI22xp33_ASAP7_75t_L g3577 ( 
.A1(n_3474),
.A2(n_3296),
.B1(n_3233),
.B2(n_3390),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3227),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3229),
.B(n_3098),
.Y(n_3579)
);

OAI22xp5_ASAP7_75t_L g3580 ( 
.A1(n_3495),
.A2(n_3167),
.B1(n_3101),
.B2(n_3104),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_3236),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3229),
.B(n_3100),
.Y(n_3582)
);

NOR2xp33_ASAP7_75t_L g3583 ( 
.A(n_3260),
.B(n_2429),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3228),
.Y(n_3584)
);

OR2x6_ASAP7_75t_L g3585 ( 
.A(n_3218),
.B(n_2934),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_SL g3586 ( 
.A(n_3364),
.B(n_2809),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3213),
.B(n_3100),
.Y(n_3587)
);

NOR2xp33_ASAP7_75t_L g3588 ( 
.A(n_3328),
.B(n_1799),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3213),
.B(n_3272),
.Y(n_3589)
);

A2O1A1Ixp33_ASAP7_75t_L g3590 ( 
.A1(n_3471),
.A2(n_3014),
.B(n_3085),
.C(n_2771),
.Y(n_3590)
);

AOI22xp5_ASAP7_75t_L g3591 ( 
.A1(n_3329),
.A2(n_3354),
.B1(n_3340),
.B2(n_3534),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3272),
.B(n_3101),
.Y(n_3592)
);

INVx2_ASAP7_75t_L g3593 ( 
.A(n_3277),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_SL g3594 ( 
.A(n_3364),
.B(n_2862),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3239),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3287),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3243),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3248),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3275),
.B(n_3467),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3288),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3275),
.B(n_3104),
.Y(n_3601)
);

INVx3_ASAP7_75t_R g3602 ( 
.A(n_3276),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_SL g3603 ( 
.A(n_3402),
.B(n_2862),
.Y(n_3603)
);

BUFx6f_ASAP7_75t_SL g3604 ( 
.A(n_3465),
.Y(n_3604)
);

NOR2xp33_ASAP7_75t_L g3605 ( 
.A(n_3417),
.B(n_1799),
.Y(n_3605)
);

AOI22xp33_ASAP7_75t_L g3606 ( 
.A1(n_3296),
.A2(n_2631),
.B1(n_2564),
.B2(n_2569),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3467),
.B(n_3251),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_SL g3608 ( 
.A(n_3516),
.B(n_2862),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_3289),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3251),
.B(n_3107),
.Y(n_3610)
);

NAND2xp33_ASAP7_75t_L g3611 ( 
.A(n_3336),
.B(n_2804),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3516),
.B(n_3384),
.Y(n_3612)
);

AOI22xp33_ASAP7_75t_L g3613 ( 
.A1(n_3233),
.A2(n_2564),
.B1(n_1830),
.B2(n_1817),
.Y(n_3613)
);

AOI22xp33_ASAP7_75t_L g3614 ( 
.A1(n_3390),
.A2(n_1830),
.B1(n_1817),
.B2(n_2488),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3315),
.B(n_3107),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3263),
.Y(n_3616)
);

OAI22xp5_ASAP7_75t_L g3617 ( 
.A1(n_3495),
.A2(n_3112),
.B1(n_3136),
.B2(n_3111),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3316),
.B(n_3111),
.Y(n_3618)
);

NAND2x1p5_ASAP7_75t_L g3619 ( 
.A(n_3337),
.B(n_2862),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3543),
.A2(n_2668),
.B1(n_3056),
.B2(n_2932),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_SL g3621 ( 
.A(n_3384),
.B(n_2862),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_R g3622 ( 
.A(n_3487),
.B(n_2558),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3312),
.Y(n_3623)
);

AND2x4_ASAP7_75t_L g3624 ( 
.A(n_3339),
.B(n_2831),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3470),
.A2(n_3056),
.B1(n_3145),
.B2(n_2687),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3314),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3265),
.Y(n_3627)
);

OAI22xp33_ASAP7_75t_L g3628 ( 
.A1(n_3231),
.A2(n_3095),
.B1(n_3105),
.B2(n_3079),
.Y(n_3628)
);

NOR2xp33_ASAP7_75t_L g3629 ( 
.A(n_3479),
.B(n_1975),
.Y(n_3629)
);

AOI22xp33_ASAP7_75t_L g3630 ( 
.A1(n_3470),
.A2(n_3564),
.B1(n_3313),
.B2(n_3253),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3266),
.Y(n_3631)
);

AOI22xp5_ASAP7_75t_L g3632 ( 
.A1(n_3437),
.A2(n_2507),
.B1(n_2524),
.B2(n_2504),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3332),
.B(n_3136),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_3244),
.B(n_2900),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3332),
.B(n_3138),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_SL g3636 ( 
.A(n_3240),
.B(n_2900),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3268),
.Y(n_3637)
);

O2A1O1Ixp5_ASAP7_75t_L g3638 ( 
.A1(n_3211),
.A2(n_3221),
.B(n_3219),
.C(n_2779),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3346),
.B(n_3138),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3270),
.Y(n_3640)
);

BUFx3_ASAP7_75t_L g3641 ( 
.A(n_3235),
.Y(n_3641)
);

BUFx3_ASAP7_75t_L g3642 ( 
.A(n_3262),
.Y(n_3642)
);

NOR3xp33_ASAP7_75t_L g3643 ( 
.A(n_3303),
.B(n_3155),
.C(n_2721),
.Y(n_3643)
);

INVxp67_ASAP7_75t_L g3644 ( 
.A(n_3269),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_SL g3645 ( 
.A(n_3442),
.B(n_2900),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3346),
.B(n_3141),
.Y(n_3646)
);

NAND2xp33_ASAP7_75t_L g3647 ( 
.A(n_3336),
.B(n_2804),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3280),
.Y(n_3648)
);

OR2x2_ASAP7_75t_L g3649 ( 
.A(n_3355),
.B(n_3208),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3283),
.Y(n_3650)
);

INVxp67_ASAP7_75t_L g3651 ( 
.A(n_3269),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_L g3652 ( 
.A1(n_3320),
.A2(n_3142),
.B1(n_3152),
.B2(n_3141),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_L g3653 ( 
.A(n_3482),
.B(n_1975),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3291),
.Y(n_3654)
);

BUFx3_ASAP7_75t_L g3655 ( 
.A(n_3305),
.Y(n_3655)
);

INVx1_ASAP7_75t_L g3656 ( 
.A(n_3293),
.Y(n_3656)
);

AND2x4_ASAP7_75t_L g3657 ( 
.A(n_3339),
.B(n_2831),
.Y(n_3657)
);

NOR2xp33_ASAP7_75t_L g3658 ( 
.A(n_3237),
.B(n_2504),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3457),
.A2(n_2524),
.B1(n_2507),
.B2(n_2538),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3301),
.Y(n_3660)
);

A2O1A1Ixp33_ASAP7_75t_L g3661 ( 
.A1(n_3232),
.A2(n_3012),
.B(n_3025),
.C(n_3022),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3377),
.B(n_3162),
.Y(n_3662)
);

OAI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_3349),
.A2(n_3162),
.B1(n_2819),
.B2(n_2821),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3309),
.Y(n_3664)
);

INVxp33_ASAP7_75t_SL g3665 ( 
.A(n_3450),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3396),
.B(n_2895),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3424),
.B(n_2871),
.Y(n_3667)
);

BUFx6f_ASAP7_75t_L g3668 ( 
.A(n_3234),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_SL g3669 ( 
.A(n_3461),
.B(n_3023),
.Y(n_3669)
);

OAI22xp33_ASAP7_75t_L g3670 ( 
.A1(n_3449),
.A2(n_3095),
.B1(n_3105),
.B2(n_3079),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3310),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3290),
.B(n_3523),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3541),
.B(n_2874),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3220),
.B(n_2604),
.Y(n_3674)
);

INVx2_ASAP7_75t_L g3675 ( 
.A(n_3318),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3222),
.B(n_3246),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3247),
.B(n_2607),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3319),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3242),
.B(n_2618),
.Y(n_3679)
);

OR2x6_ASAP7_75t_L g3680 ( 
.A(n_3218),
.B(n_2934),
.Y(n_3680)
);

OR2x6_ASAP7_75t_L g3681 ( 
.A(n_3218),
.B(n_3438),
.Y(n_3681)
);

NAND2xp33_ASAP7_75t_L g3682 ( 
.A(n_3336),
.B(n_2804),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3255),
.B(n_2620),
.Y(n_3683)
);

INVxp67_ASAP7_75t_L g3684 ( 
.A(n_3352),
.Y(n_3684)
);

INVx2_ASAP7_75t_L g3685 ( 
.A(n_3324),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3323),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3531),
.B(n_2549),
.Y(n_3687)
);

NAND2xp5_ASAP7_75t_SL g3688 ( 
.A(n_3556),
.B(n_3023),
.Y(n_3688)
);

AOI22xp33_ASAP7_75t_L g3689 ( 
.A1(n_3313),
.A2(n_3145),
.B1(n_3056),
.B2(n_2449),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3556),
.B(n_3023),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3391),
.B(n_3397),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3348),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3358),
.Y(n_3693)
);

BUFx6f_ASAP7_75t_L g3694 ( 
.A(n_3234),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_L g3695 ( 
.A(n_3391),
.B(n_2620),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3360),
.Y(n_3696)
);

NOR2xp33_ASAP7_75t_L g3697 ( 
.A(n_3454),
.B(n_2553),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3397),
.B(n_2622),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3379),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3448),
.B(n_2622),
.Y(n_3700)
);

INVx2_ASAP7_75t_L g3701 ( 
.A(n_3383),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3387),
.Y(n_3702)
);

BUFx3_ASAP7_75t_L g3703 ( 
.A(n_3245),
.Y(n_3703)
);

AO22x2_ASAP7_75t_L g3704 ( 
.A1(n_3563),
.A2(n_3005),
.B1(n_3053),
.B2(n_3050),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3464),
.B(n_2626),
.Y(n_3705)
);

NOR2xp33_ASAP7_75t_L g3706 ( 
.A(n_3455),
.B(n_2426),
.Y(n_3706)
);

AND2x4_ASAP7_75t_L g3707 ( 
.A(n_3339),
.B(n_2866),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_L g3708 ( 
.A(n_3292),
.B(n_2427),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3370),
.B(n_2626),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3399),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3252),
.B(n_3023),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_SL g3712 ( 
.A(n_3365),
.B(n_3023),
.Y(n_3712)
);

NAND2xp5_ASAP7_75t_L g3713 ( 
.A(n_3458),
.B(n_2635),
.Y(n_3713)
);

INVx3_ASAP7_75t_L g3714 ( 
.A(n_3551),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3458),
.B(n_2635),
.Y(n_3715)
);

NOR2xp67_ASAP7_75t_SL g3716 ( 
.A(n_3215),
.B(n_2427),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3409),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3446),
.B(n_2445),
.Y(n_3718)
);

CKINVDCx5p33_ASAP7_75t_R g3719 ( 
.A(n_3225),
.Y(n_3719)
);

NAND2xp5_ASAP7_75t_L g3720 ( 
.A(n_3373),
.B(n_2636),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3373),
.B(n_2636),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3554),
.B(n_2638),
.Y(n_3722)
);

NOR2xp67_ASAP7_75t_SL g3723 ( 
.A(n_3267),
.B(n_2465),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3330),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3331),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3473),
.B(n_3492),
.Y(n_3726)
);

NOR2xp33_ASAP7_75t_L g3727 ( 
.A(n_3341),
.B(n_2465),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_SL g3728 ( 
.A(n_3365),
.B(n_2983),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_L g3729 ( 
.A(n_3473),
.B(n_2638),
.Y(n_3729)
);

OAI22xp5_ASAP7_75t_L g3730 ( 
.A1(n_3217),
.A2(n_3105),
.B1(n_3095),
.B2(n_3180),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3335),
.Y(n_3731)
);

INVx2_ASAP7_75t_L g3732 ( 
.A(n_3416),
.Y(n_3732)
);

AND2x4_ASAP7_75t_L g3733 ( 
.A(n_3481),
.B(n_2866),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3359),
.B(n_2466),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3403),
.B(n_3419),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3343),
.B(n_2651),
.Y(n_3736)
);

BUFx6f_ASAP7_75t_L g3737 ( 
.A(n_3234),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3426),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3433),
.Y(n_3739)
);

CKINVDCx16_ASAP7_75t_R g3740 ( 
.A(n_3256),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3344),
.B(n_2651),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_3366),
.B(n_2466),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3350),
.B(n_2653),
.Y(n_3743)
);

BUFx5_ASAP7_75t_L g3744 ( 
.A(n_3551),
.Y(n_3744)
);

NAND2xp5_ASAP7_75t_L g3745 ( 
.A(n_3357),
.B(n_2655),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3361),
.B(n_2655),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_3367),
.B(n_2659),
.Y(n_3747)
);

NOR2xp67_ASAP7_75t_L g3748 ( 
.A(n_3509),
.B(n_2559),
.Y(n_3748)
);

NAND2xp5_ASAP7_75t_L g3749 ( 
.A(n_3369),
.B(n_2659),
.Y(n_3749)
);

AND2x4_ASAP7_75t_L g3750 ( 
.A(n_3481),
.B(n_3092),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3371),
.B(n_2666),
.Y(n_3751)
);

AOI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_3429),
.A2(n_2475),
.B1(n_2477),
.B2(n_2479),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3374),
.Y(n_3753)
);

INVxp67_ASAP7_75t_SL g3754 ( 
.A(n_3460),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3376),
.B(n_2666),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_SL g3756 ( 
.A(n_3249),
.B(n_2786),
.Y(n_3756)
);

NOR2xp33_ASAP7_75t_L g3757 ( 
.A(n_3440),
.B(n_2475),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3382),
.B(n_2675),
.Y(n_3758)
);

AOI22xp5_ASAP7_75t_L g3759 ( 
.A1(n_3429),
.A2(n_2477),
.B1(n_2484),
.B2(n_2479),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_3434),
.Y(n_3760)
);

BUFx6f_ASAP7_75t_L g3761 ( 
.A(n_3264),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3217),
.B(n_2952),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_SL g3763 ( 
.A(n_3249),
.B(n_3095),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3232),
.B(n_2952),
.Y(n_3764)
);

BUFx3_ASAP7_75t_L g3765 ( 
.A(n_3245),
.Y(n_3765)
);

INVx2_ASAP7_75t_L g3766 ( 
.A(n_3441),
.Y(n_3766)
);

AND2x2_ASAP7_75t_L g3767 ( 
.A(n_3313),
.B(n_2047),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_L g3768 ( 
.A(n_3214),
.B(n_3226),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3445),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3214),
.B(n_2953),
.Y(n_3770)
);

INVx8_ASAP7_75t_L g3771 ( 
.A(n_3466),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3226),
.B(n_2953),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3392),
.B(n_2956),
.Y(n_3773)
);

NOR2xp33_ASAP7_75t_L g3774 ( 
.A(n_3535),
.B(n_2484),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3394),
.B(n_2956),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_3400),
.Y(n_3776)
);

OAI21xp5_ASAP7_75t_L g3777 ( 
.A1(n_3219),
.A2(n_3005),
.B(n_3102),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3404),
.Y(n_3778)
);

NAND2xp33_ASAP7_75t_L g3779 ( 
.A(n_3336),
.B(n_2934),
.Y(n_3779)
);

INVx2_ASAP7_75t_L g3780 ( 
.A(n_3456),
.Y(n_3780)
);

BUFx6f_ASAP7_75t_SL g3781 ( 
.A(n_3465),
.Y(n_3781)
);

NOR2xp33_ASAP7_75t_L g3782 ( 
.A(n_3517),
.B(n_2500),
.Y(n_3782)
);

AOI22xp5_ASAP7_75t_L g3783 ( 
.A1(n_3429),
.A2(n_2500),
.B1(n_2511),
.B2(n_2510),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3406),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3412),
.B(n_2957),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3475),
.Y(n_3786)
);

INVxp67_ASAP7_75t_SL g3787 ( 
.A(n_3460),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3480),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3493),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_L g3790 ( 
.A(n_3413),
.B(n_2957),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3415),
.B(n_2964),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3421),
.B(n_2964),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3533),
.Y(n_3793)
);

INVx1_ASAP7_75t_SL g3794 ( 
.A(n_3261),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3422),
.Y(n_3795)
);

INVx2_ASAP7_75t_L g3796 ( 
.A(n_3549),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3550),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3423),
.B(n_2966),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_L g3799 ( 
.A(n_3435),
.B(n_2966),
.Y(n_3799)
);

NAND2xp33_ASAP7_75t_SL g3800 ( 
.A(n_3299),
.B(n_3145),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3476),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3483),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_SL g3803 ( 
.A(n_3261),
.B(n_3206),
.Y(n_3803)
);

AND2x2_ASAP7_75t_L g3804 ( 
.A(n_3520),
.B(n_2047),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3557),
.Y(n_3805)
);

OAI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3432),
.A2(n_2516),
.B1(n_2520),
.B2(n_2510),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_SL g3807 ( 
.A(n_3302),
.B(n_3182),
.Y(n_3807)
);

NOR3xp33_ASAP7_75t_L g3808 ( 
.A(n_3216),
.B(n_3082),
.C(n_3040),
.Y(n_3808)
);

INVx2_ASAP7_75t_L g3809 ( 
.A(n_3570),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_SL g3810 ( 
.A(n_3302),
.B(n_3009),
.Y(n_3810)
);

AND2x4_ASAP7_75t_L g3811 ( 
.A(n_3286),
.B(n_3509),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3485),
.B(n_2898),
.Y(n_3812)
);

AND2x2_ASAP7_75t_L g3813 ( 
.A(n_3307),
.B(n_2047),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_SL g3814 ( 
.A(n_3224),
.B(n_3009),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_L g3815 ( 
.A(n_3489),
.B(n_2898),
.Y(n_3815)
);

AOI22xp5_ASAP7_75t_L g3816 ( 
.A1(n_3285),
.A2(n_2526),
.B1(n_2890),
.B2(n_2545),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3496),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_SL g3818 ( 
.A(n_3224),
.B(n_3009),
.Y(n_3818)
);

INVx2_ASAP7_75t_L g3819 ( 
.A(n_3500),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3478),
.B(n_3009),
.Y(n_3820)
);

INVx2_ASAP7_75t_SL g3821 ( 
.A(n_3298),
.Y(n_3821)
);

AOI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_3285),
.A2(n_2526),
.B1(n_2890),
.B2(n_2543),
.Y(n_3822)
);

OR2x6_ASAP7_75t_L g3823 ( 
.A(n_3438),
.B(n_2949),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3501),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3522),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_SL g3826 ( 
.A(n_3286),
.B(n_3009),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_3524),
.B(n_2901),
.Y(n_3827)
);

BUFx6f_ASAP7_75t_L g3828 ( 
.A(n_3264),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3527),
.B(n_2901),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3530),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3532),
.B(n_2904),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_SL g3832 ( 
.A(n_3555),
.B(n_3044),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3542),
.B(n_2904),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_L g3834 ( 
.A(n_3546),
.B(n_2906),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_SL g3835 ( 
.A(n_3210),
.B(n_2949),
.Y(n_3835)
);

HB1xp67_ASAP7_75t_L g3836 ( 
.A(n_3512),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3552),
.Y(n_3837)
);

OR2x6_ASAP7_75t_L g3838 ( 
.A(n_3438),
.B(n_2949),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3555),
.B(n_3044),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_3553),
.B(n_2906),
.Y(n_3840)
);

INVxp67_ASAP7_75t_L g3841 ( 
.A(n_3386),
.Y(n_3841)
);

OR2x6_ASAP7_75t_L g3842 ( 
.A(n_3518),
.B(n_2949),
.Y(n_3842)
);

BUFx5_ASAP7_75t_L g3843 ( 
.A(n_3551),
.Y(n_3843)
);

AOI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3253),
.A2(n_2449),
.B1(n_2482),
.B2(n_2414),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3565),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3431),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_L g3847 ( 
.A(n_3253),
.B(n_2907),
.Y(n_3847)
);

NOR2xp33_ASAP7_75t_L g3848 ( 
.A(n_3511),
.B(n_3028),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3253),
.B(n_3271),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3431),
.Y(n_3850)
);

INVx2_ASAP7_75t_SL g3851 ( 
.A(n_3327),
.Y(n_3851)
);

AO221x1_ASAP7_75t_L g3852 ( 
.A1(n_3525),
.A2(n_742),
.B1(n_815),
.B2(n_693),
.C(n_676),
.Y(n_3852)
);

AND2x4_ASAP7_75t_L g3853 ( 
.A(n_3519),
.B(n_3545),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3447),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_L g3855 ( 
.A(n_3271),
.B(n_2907),
.Y(n_3855)
);

INVx3_ASAP7_75t_L g3856 ( 
.A(n_3551),
.Y(n_3856)
);

INVx5_ASAP7_75t_L g3857 ( 
.A(n_3466),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3511),
.B(n_2082),
.Y(n_3858)
);

AND2x4_ASAP7_75t_L g3859 ( 
.A(n_3519),
.B(n_3137),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3526),
.Y(n_3860)
);

INVxp33_ASAP7_75t_L g3861 ( 
.A(n_3327),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3250),
.B(n_2910),
.Y(n_3862)
);

CKINVDCx5p33_ASAP7_75t_R g3863 ( 
.A(n_3338),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3526),
.Y(n_3864)
);

OAI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3432),
.A2(n_2729),
.B1(n_2723),
.B2(n_2648),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_3486),
.B(n_3036),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3250),
.B(n_2910),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3425),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3273),
.B(n_2911),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3447),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3254),
.B(n_3044),
.Y(n_3871)
);

OAI21xp5_ASAP7_75t_L g3872 ( 
.A1(n_3221),
.A2(n_3223),
.B(n_3200),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_SL g3873 ( 
.A(n_3258),
.B(n_3044),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3484),
.B(n_2082),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3273),
.B(n_2911),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3545),
.B(n_3322),
.Y(n_3876)
);

AOI221xp5_ASAP7_75t_L g3877 ( 
.A1(n_3525),
.A2(n_1456),
.B1(n_1467),
.B2(n_1461),
.C(n_1459),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_3558),
.B(n_3037),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3451),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3281),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3569),
.B(n_3063),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3281),
.Y(n_3882)
);

AND2x4_ASAP7_75t_L g3883 ( 
.A(n_3322),
.B(n_3351),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3484),
.B(n_2082),
.Y(n_3884)
);

INVx2_ASAP7_75t_SL g3885 ( 
.A(n_3425),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3451),
.Y(n_3886)
);

INVx1_ASAP7_75t_L g3887 ( 
.A(n_3284),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3453),
.Y(n_3888)
);

BUFx2_ASAP7_75t_L g3889 ( 
.A(n_3414),
.Y(n_3889)
);

AND2x4_ASAP7_75t_L g3890 ( 
.A(n_3351),
.B(n_3137),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3453),
.Y(n_3891)
);

NAND2x1_ASAP7_75t_L g3892 ( 
.A(n_3230),
.B(n_2842),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_L g3893 ( 
.A(n_3284),
.B(n_3259),
.Y(n_3893)
);

NOR2xp67_ASAP7_75t_L g3894 ( 
.A(n_3342),
.B(n_2573),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3463),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3259),
.B(n_2912),
.Y(n_3896)
);

OR2x2_ASAP7_75t_L g3897 ( 
.A(n_3212),
.B(n_3065),
.Y(n_3897)
);

AND2x4_ASAP7_75t_L g3898 ( 
.A(n_3389),
.B(n_3439),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_L g3899 ( 
.A(n_3539),
.B(n_2043),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3463),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3539),
.B(n_3561),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3488),
.B(n_2043),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3494),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3494),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3819),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3735),
.B(n_3573),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3581),
.Y(n_3907)
);

BUFx6f_ASAP7_75t_L g3908 ( 
.A(n_3771),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3824),
.Y(n_3909)
);

BUFx4f_ASAP7_75t_L g3910 ( 
.A(n_3771),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3825),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3830),
.Y(n_3912)
);

INVx3_ASAP7_75t_L g3913 ( 
.A(n_3714),
.Y(n_3913)
);

AND2x2_ASAP7_75t_L g3914 ( 
.A(n_3849),
.B(n_3525),
.Y(n_3914)
);

OR2x2_ASAP7_75t_L g3915 ( 
.A(n_3849),
.B(n_3363),
.Y(n_3915)
);

INVx3_ASAP7_75t_L g3916 ( 
.A(n_3714),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3860),
.B(n_3510),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3864),
.B(n_3510),
.Y(n_3918)
);

HB1xp67_ASAP7_75t_L g3919 ( 
.A(n_3644),
.Y(n_3919)
);

BUFx3_ASAP7_75t_L g3920 ( 
.A(n_3641),
.Y(n_3920)
);

INVx3_ASAP7_75t_L g3921 ( 
.A(n_3856),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3593),
.Y(n_3922)
);

BUFx6f_ASAP7_75t_L g3923 ( 
.A(n_3771),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3596),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_3672),
.B(n_3572),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3600),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3845),
.B(n_3538),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3584),
.B(n_3538),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3609),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3666),
.B(n_3521),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_L g3931 ( 
.A(n_3662),
.B(n_3558),
.Y(n_3931)
);

INVxp67_ASAP7_75t_SL g3932 ( 
.A(n_3607),
.Y(n_3932)
);

INVx3_ASAP7_75t_L g3933 ( 
.A(n_3856),
.Y(n_3933)
);

BUFx3_ASAP7_75t_L g3934 ( 
.A(n_3642),
.Y(n_3934)
);

AND2x4_ASAP7_75t_L g3935 ( 
.A(n_3681),
.B(n_3304),
.Y(n_3935)
);

INVx4_ASAP7_75t_L g3936 ( 
.A(n_3857),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3623),
.Y(n_3937)
);

BUFx3_ASAP7_75t_L g3938 ( 
.A(n_3655),
.Y(n_3938)
);

BUFx5_ASAP7_75t_L g3939 ( 
.A(n_3880),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3595),
.Y(n_3940)
);

AND2x2_ASAP7_75t_L g3941 ( 
.A(n_3597),
.B(n_3598),
.Y(n_3941)
);

BUFx6f_ASAP7_75t_L g3942 ( 
.A(n_3857),
.Y(n_3942)
);

AND2x2_ASAP7_75t_SL g3943 ( 
.A(n_3611),
.B(n_3238),
.Y(n_3943)
);

INVx5_ASAP7_75t_L g3944 ( 
.A(n_3857),
.Y(n_3944)
);

INVx3_ASAP7_75t_SL g3945 ( 
.A(n_3719),
.Y(n_3945)
);

AND2x4_ASAP7_75t_L g3946 ( 
.A(n_3681),
.B(n_3304),
.Y(n_3946)
);

OR2x2_ASAP7_75t_L g3947 ( 
.A(n_3599),
.B(n_3754),
.Y(n_3947)
);

INVx8_ASAP7_75t_L g3948 ( 
.A(n_3857),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3726),
.B(n_3561),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_3676),
.B(n_3566),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_3615),
.B(n_3618),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3681),
.Y(n_3952)
);

INVx1_ASAP7_75t_SL g3953 ( 
.A(n_3622),
.Y(n_3953)
);

INVx4_ASAP7_75t_L g3954 ( 
.A(n_3823),
.Y(n_3954)
);

AND2x2_ASAP7_75t_L g3955 ( 
.A(n_3616),
.B(n_3259),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_L g3956 ( 
.A(n_3633),
.B(n_3491),
.Y(n_3956)
);

OAI21xp5_ASAP7_75t_L g3957 ( 
.A1(n_3591),
.A2(n_3200),
.B(n_2810),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3627),
.B(n_3259),
.Y(n_3958)
);

OR2x2_ASAP7_75t_L g3959 ( 
.A(n_3599),
.B(n_3363),
.Y(n_3959)
);

AND2x2_ASAP7_75t_L g3960 ( 
.A(n_3631),
.B(n_3308),
.Y(n_3960)
);

INVxp67_ASAP7_75t_SL g3961 ( 
.A(n_3607),
.Y(n_3961)
);

INVx2_ASAP7_75t_L g3962 ( 
.A(n_3626),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3637),
.B(n_3308),
.Y(n_3963)
);

INVx2_ASAP7_75t_SL g3964 ( 
.A(n_3668),
.Y(n_3964)
);

OAI21xp5_ASAP7_75t_L g3965 ( 
.A1(n_3638),
.A2(n_2915),
.B(n_2886),
.Y(n_3965)
);

INVxp67_ASAP7_75t_L g3966 ( 
.A(n_3691),
.Y(n_3966)
);

HB1xp67_ASAP7_75t_L g3967 ( 
.A(n_3651),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3635),
.B(n_3513),
.Y(n_3968)
);

AND2x2_ASAP7_75t_L g3969 ( 
.A(n_3640),
.B(n_3317),
.Y(n_3969)
);

INVx8_ASAP7_75t_L g3970 ( 
.A(n_3585),
.Y(n_3970)
);

AND2x2_ASAP7_75t_SL g3971 ( 
.A(n_3647),
.B(n_3490),
.Y(n_3971)
);

INVx3_ASAP7_75t_SL g3972 ( 
.A(n_3863),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3648),
.B(n_3317),
.Y(n_3973)
);

OR2x2_ASAP7_75t_L g3974 ( 
.A(n_3787),
.B(n_3385),
.Y(n_3974)
);

HB1xp67_ASAP7_75t_L g3975 ( 
.A(n_3684),
.Y(n_3975)
);

OAI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3590),
.A2(n_2918),
.B(n_2916),
.Y(n_3976)
);

INVxp67_ASAP7_75t_L g3977 ( 
.A(n_3576),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3639),
.B(n_3537),
.Y(n_3978)
);

BUFx3_ASAP7_75t_L g3979 ( 
.A(n_3703),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3650),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3654),
.B(n_3356),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_3646),
.B(n_2987),
.Y(n_3982)
);

HB1xp67_ASAP7_75t_L g3983 ( 
.A(n_3836),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3656),
.B(n_3356),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3667),
.B(n_2989),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_SL g3986 ( 
.A(n_3580),
.B(n_3223),
.Y(n_3986)
);

NAND2x1p5_ASAP7_75t_L g3987 ( 
.A(n_3794),
.B(n_3337),
.Y(n_3987)
);

INVx2_ASAP7_75t_SL g3988 ( 
.A(n_3668),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3675),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3660),
.B(n_3362),
.Y(n_3990)
);

BUFx3_ASAP7_75t_L g3991 ( 
.A(n_3765),
.Y(n_3991)
);

INVx2_ASAP7_75t_L g3992 ( 
.A(n_3678),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3664),
.B(n_3362),
.Y(n_3993)
);

BUFx3_ASAP7_75t_L g3994 ( 
.A(n_3868),
.Y(n_3994)
);

AND2x2_ASAP7_75t_L g3995 ( 
.A(n_3671),
.B(n_3368),
.Y(n_3995)
);

BUFx6f_ASAP7_75t_L g3996 ( 
.A(n_3750),
.Y(n_3996)
);

INVxp33_ASAP7_75t_L g3997 ( 
.A(n_3718),
.Y(n_3997)
);

OR2x2_ASAP7_75t_L g3998 ( 
.A(n_3847),
.B(n_3385),
.Y(n_3998)
);

INVx2_ASAP7_75t_SL g3999 ( 
.A(n_3668),
.Y(n_3999)
);

INVx2_ASAP7_75t_SL g4000 ( 
.A(n_3694),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3686),
.B(n_3368),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3673),
.B(n_3439),
.Y(n_4002)
);

AND2x4_ASAP7_75t_L g4003 ( 
.A(n_3585),
.B(n_3680),
.Y(n_4003)
);

AND2x2_ASAP7_75t_SL g4004 ( 
.A(n_3682),
.B(n_3241),
.Y(n_4004)
);

NAND2x1p5_ASAP7_75t_L g4005 ( 
.A(n_3794),
.B(n_3337),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3685),
.Y(n_4006)
);

INVx1_ASAP7_75t_SL g4007 ( 
.A(n_3889),
.Y(n_4007)
);

BUFx6f_ASAP7_75t_L g4008 ( 
.A(n_3750),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3724),
.Y(n_4009)
);

INVx2_ASAP7_75t_SL g4010 ( 
.A(n_3694),
.Y(n_4010)
);

INVx3_ASAP7_75t_L g4011 ( 
.A(n_3744),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3725),
.B(n_3380),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3692),
.Y(n_4013)
);

INVx1_ASAP7_75t_SL g4014 ( 
.A(n_3695),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3731),
.B(n_3380),
.Y(n_4015)
);

OR2x2_ASAP7_75t_L g4016 ( 
.A(n_3847),
.B(n_3398),
.Y(n_4016)
);

INVx3_ASAP7_75t_L g4017 ( 
.A(n_3744),
.Y(n_4017)
);

OAI21xp5_ASAP7_75t_L g4018 ( 
.A1(n_3877),
.A2(n_2941),
.B(n_2927),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3693),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3753),
.B(n_3407),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3696),
.Y(n_4021)
);

BUFx6f_ASAP7_75t_L g4022 ( 
.A(n_3890),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3699),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3776),
.B(n_3407),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_3778),
.B(n_3436),
.Y(n_4025)
);

INVxp67_ASAP7_75t_L g4026 ( 
.A(n_3574),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3784),
.B(n_3436),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3729),
.B(n_2998),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3795),
.B(n_3443),
.Y(n_4029)
);

INVx2_ASAP7_75t_SL g4030 ( 
.A(n_3694),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3801),
.B(n_3443),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3802),
.B(n_3444),
.Y(n_4032)
);

HB1xp67_ASAP7_75t_L g4033 ( 
.A(n_3578),
.Y(n_4033)
);

BUFx3_ASAP7_75t_L g4034 ( 
.A(n_3853),
.Y(n_4034)
);

INVx2_ASAP7_75t_L g4035 ( 
.A(n_3701),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3702),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3817),
.B(n_3444),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3710),
.Y(n_4038)
);

OAI21xp33_ASAP7_75t_L g4039 ( 
.A1(n_3580),
.A2(n_1461),
.B(n_1459),
.Y(n_4039)
);

INVx2_ASAP7_75t_L g4040 ( 
.A(n_3717),
.Y(n_4040)
);

AND2x4_ASAP7_75t_L g4041 ( 
.A(n_3585),
.B(n_3452),
.Y(n_4041)
);

OAI21xp5_ASAP7_75t_L g4042 ( 
.A1(n_3663),
.A2(n_2961),
.B(n_2960),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3579),
.B(n_3024),
.Y(n_4043)
);

AND2x2_ASAP7_75t_SL g4044 ( 
.A(n_3630),
.B(n_3241),
.Y(n_4044)
);

NOR2xp33_ASAP7_75t_SL g4045 ( 
.A(n_3774),
.B(n_2412),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_L g4046 ( 
.A(n_3579),
.B(n_3544),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3582),
.B(n_3544),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3732),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_3680),
.B(n_3452),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_3837),
.B(n_3325),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3846),
.B(n_3325),
.Y(n_4051)
);

OAI21xp33_ASAP7_75t_L g4052 ( 
.A1(n_3605),
.A2(n_1468),
.B(n_1467),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3850),
.B(n_3334),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3854),
.B(n_3334),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3738),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3588),
.B(n_2729),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3739),
.Y(n_4057)
);

INVx3_ASAP7_75t_L g4058 ( 
.A(n_3744),
.Y(n_4058)
);

AND2x6_ASAP7_75t_L g4059 ( 
.A(n_3893),
.B(n_3241),
.Y(n_4059)
);

BUFx3_ASAP7_75t_L g4060 ( 
.A(n_3853),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3582),
.B(n_3050),
.Y(n_4061)
);

INVx2_ASAP7_75t_L g4062 ( 
.A(n_3760),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3766),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_SL g4064 ( 
.A(n_3589),
.B(n_3264),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3769),
.Y(n_4065)
);

INVx4_ASAP7_75t_L g4066 ( 
.A(n_3823),
.Y(n_4066)
);

BUFx6f_ASAP7_75t_L g4067 ( 
.A(n_3890),
.Y(n_4067)
);

INVx1_ASAP7_75t_L g4068 ( 
.A(n_3780),
.Y(n_4068)
);

AND2x4_ASAP7_75t_SL g4069 ( 
.A(n_3680),
.B(n_3488),
.Y(n_4069)
);

INVx3_ASAP7_75t_L g4070 ( 
.A(n_3744),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3589),
.B(n_3278),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_SL g4072 ( 
.A(n_3663),
.B(n_3893),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_3649),
.B(n_3053),
.Y(n_4073)
);

AND2x2_ASAP7_75t_L g4074 ( 
.A(n_3870),
.B(n_3241),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3786),
.Y(n_4075)
);

CKINVDCx5p33_ASAP7_75t_R g4076 ( 
.A(n_3665),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3788),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3789),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3610),
.B(n_3055),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3793),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3652),
.B(n_3278),
.Y(n_4081)
);

OAI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_3661),
.A2(n_2973),
.B(n_2967),
.Y(n_4082)
);

AND2x2_ASAP7_75t_L g4083 ( 
.A(n_3879),
.B(n_3398),
.Y(n_4083)
);

NAND2x1p5_ASAP7_75t_L g4084 ( 
.A(n_3608),
.B(n_3337),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3823),
.B(n_3498),
.Y(n_4085)
);

AND2x2_ASAP7_75t_SL g4086 ( 
.A(n_3835),
.B(n_3560),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3796),
.Y(n_4087)
);

CKINVDCx20_ASAP7_75t_R g4088 ( 
.A(n_3740),
.Y(n_4088)
);

NOR2xp67_ASAP7_75t_L g4089 ( 
.A(n_3821),
.B(n_3395),
.Y(n_4089)
);

AND2x4_ASAP7_75t_L g4090 ( 
.A(n_3838),
.B(n_3498),
.Y(n_4090)
);

NOR2xp33_ASAP7_75t_SL g4091 ( 
.A(n_3723),
.B(n_2412),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_3797),
.Y(n_4092)
);

INVx2_ASAP7_75t_L g4093 ( 
.A(n_3805),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3886),
.B(n_3401),
.Y(n_4094)
);

INVxp67_ASAP7_75t_SL g4095 ( 
.A(n_3592),
.Y(n_4095)
);

INVx1_ASAP7_75t_SL g4096 ( 
.A(n_3698),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3809),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3888),
.Y(n_4098)
);

AND2x2_ASAP7_75t_SL g4099 ( 
.A(n_3835),
.B(n_3779),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_L g4100 ( 
.A(n_3583),
.B(n_2416),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3773),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3891),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3900),
.B(n_3401),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3773),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3767),
.B(n_3405),
.Y(n_4105)
);

BUFx3_ASAP7_75t_L g4106 ( 
.A(n_3811),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_3704),
.B(n_3895),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_3652),
.B(n_3278),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3775),
.Y(n_4109)
);

HB1xp67_ASAP7_75t_L g4110 ( 
.A(n_3592),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3775),
.Y(n_4111)
);

BUFx3_ASAP7_75t_L g4112 ( 
.A(n_3811),
.Y(n_4112)
);

HB1xp67_ASAP7_75t_L g4113 ( 
.A(n_3601),
.Y(n_4113)
);

AND2x2_ASAP7_75t_SL g4114 ( 
.A(n_3689),
.B(n_3560),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_3704),
.B(n_3405),
.Y(n_4115)
);

HB1xp67_ASAP7_75t_L g4116 ( 
.A(n_3601),
.Y(n_4116)
);

BUFx6f_ASAP7_75t_L g4117 ( 
.A(n_3838),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3785),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_3713),
.B(n_3066),
.Y(n_4119)
);

INVx3_ASAP7_75t_L g4120 ( 
.A(n_3744),
.Y(n_4120)
);

INVx2_ASAP7_75t_L g4121 ( 
.A(n_3790),
.Y(n_4121)
);

HB1xp67_ASAP7_75t_L g4122 ( 
.A(n_3617),
.Y(n_4122)
);

INVx2_ASAP7_75t_L g4123 ( 
.A(n_3791),
.Y(n_4123)
);

NOR2xp33_ASAP7_75t_L g4124 ( 
.A(n_3708),
.B(n_2416),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_3903),
.B(n_3408),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_3904),
.B(n_3408),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_3882),
.B(n_3887),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_SL g4128 ( 
.A(n_3843),
.B(n_3279),
.Y(n_4128)
);

BUFx6f_ASAP7_75t_L g4129 ( 
.A(n_3838),
.Y(n_4129)
);

AND2x2_ASAP7_75t_SL g4130 ( 
.A(n_3577),
.B(n_3300),
.Y(n_4130)
);

NOR2xp33_ASAP7_75t_L g4131 ( 
.A(n_3677),
.B(n_2419),
.Y(n_4131)
);

INVx3_ASAP7_75t_L g4132 ( 
.A(n_3843),
.Y(n_4132)
);

BUFx6f_ASAP7_75t_L g4133 ( 
.A(n_3842),
.Y(n_4133)
);

HB1xp67_ASAP7_75t_L g4134 ( 
.A(n_3617),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_3602),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_3715),
.B(n_3066),
.Y(n_4136)
);

HB1xp67_ASAP7_75t_L g4137 ( 
.A(n_3881),
.Y(n_4137)
);

AND2x2_ASAP7_75t_L g4138 ( 
.A(n_3874),
.B(n_3884),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_3842),
.B(n_3504),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3720),
.B(n_3068),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3792),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3721),
.B(n_3709),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3798),
.Y(n_4143)
);

INVx2_ASAP7_75t_SL g4144 ( 
.A(n_3737),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3799),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_3587),
.B(n_3068),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3799),
.Y(n_4147)
);

AND2x2_ASAP7_75t_L g4148 ( 
.A(n_3587),
.B(n_3768),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3812),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_3812),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3737),
.Y(n_4151)
);

AND2x4_ASAP7_75t_L g4152 ( 
.A(n_3842),
.B(n_3504),
.Y(n_4152)
);

INVx3_ASAP7_75t_L g4153 ( 
.A(n_3843),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3813),
.B(n_3070),
.Y(n_4154)
);

BUFx2_ASAP7_75t_L g4155 ( 
.A(n_3859),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3815),
.Y(n_4156)
);

INVx2_ASAP7_75t_SL g4157 ( 
.A(n_3761),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_3815),
.Y(n_4158)
);

BUFx2_ASAP7_75t_L g4159 ( 
.A(n_3859),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_3768),
.B(n_3418),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3827),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3901),
.B(n_3418),
.Y(n_4162)
);

AND2x2_ASAP7_75t_SL g4163 ( 
.A(n_3625),
.B(n_3300),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_SL g4164 ( 
.A(n_3843),
.B(n_3730),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_L g4165 ( 
.A(n_3878),
.B(n_3070),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_3683),
.B(n_3674),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3827),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3829),
.Y(n_4168)
);

INVx2_ASAP7_75t_SL g4169 ( 
.A(n_3761),
.Y(n_4169)
);

NAND2x1p5_ASAP7_75t_L g4170 ( 
.A(n_3612),
.B(n_3353),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_3829),
.B(n_3427),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_3831),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3804),
.B(n_3072),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3831),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_3833),
.B(n_3427),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3700),
.B(n_3074),
.Y(n_4176)
);

INVx4_ASAP7_75t_L g4177 ( 
.A(n_3828),
.Y(n_4177)
);

INVx1_ASAP7_75t_SL g4178 ( 
.A(n_3782),
.Y(n_4178)
);

INVx2_ASAP7_75t_L g4179 ( 
.A(n_3833),
.Y(n_4179)
);

INVxp67_ASAP7_75t_L g4180 ( 
.A(n_3734),
.Y(n_4180)
);

OAI21xp5_ASAP7_75t_L g4181 ( 
.A1(n_3777),
.A2(n_2981),
.B(n_2974),
.Y(n_4181)
);

CKINVDCx20_ASAP7_75t_R g4182 ( 
.A(n_3659),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3834),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_3705),
.B(n_3736),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_3834),
.Y(n_4185)
);

AND2x4_ASAP7_75t_L g4186 ( 
.A(n_3624),
.B(n_3505),
.Y(n_4186)
);

AND2x4_ASAP7_75t_SL g4187 ( 
.A(n_3883),
.B(n_3898),
.Y(n_4187)
);

INVx2_ASAP7_75t_L g4188 ( 
.A(n_3840),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_3741),
.B(n_3743),
.Y(n_4189)
);

NOR2xp33_ASAP7_75t_L g4190 ( 
.A(n_3679),
.B(n_2419),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_3840),
.Y(n_4191)
);

INVx2_ASAP7_75t_L g4192 ( 
.A(n_3764),
.Y(n_4192)
);

AND2x2_ASAP7_75t_L g4193 ( 
.A(n_3855),
.B(n_3300),
.Y(n_4193)
);

NOR2xp67_ASAP7_75t_L g4194 ( 
.A(n_3851),
.B(n_3885),
.Y(n_4194)
);

OAI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_3777),
.A2(n_2986),
.B(n_2788),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_3764),
.Y(n_4196)
);

BUFx2_ASAP7_75t_L g4197 ( 
.A(n_3896),
.Y(n_4197)
);

INVx2_ASAP7_75t_SL g4198 ( 
.A(n_3828),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_L g4199 ( 
.A(n_3658),
.B(n_2469),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_3772),
.Y(n_4200)
);

INVx1_ASAP7_75t_SL g4201 ( 
.A(n_3742),
.Y(n_4201)
);

BUFx6f_ASAP7_75t_L g4202 ( 
.A(n_3828),
.Y(n_4202)
);

NOR2xp33_ASAP7_75t_SL g4203 ( 
.A(n_3697),
.B(n_2648),
.Y(n_4203)
);

HB1xp67_ASAP7_75t_L g4204 ( 
.A(n_3810),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3772),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_3745),
.B(n_3074),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3746),
.B(n_3080),
.Y(n_4207)
);

AND2x4_ASAP7_75t_L g4208 ( 
.A(n_3624),
.B(n_3505),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3747),
.B(n_3080),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_3862),
.Y(n_4210)
);

INVx2_ASAP7_75t_L g4211 ( 
.A(n_3862),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_3855),
.B(n_3326),
.Y(n_4212)
);

NOR2xp67_ASAP7_75t_L g4213 ( 
.A(n_3816),
.B(n_3353),
.Y(n_4213)
);

INVxp33_ASAP7_75t_L g4214 ( 
.A(n_3757),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_SL g4215 ( 
.A(n_3706),
.B(n_2665),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_SL g4216 ( 
.A(n_3730),
.B(n_3279),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_3872),
.B(n_3326),
.Y(n_4217)
);

NAND2xp5_ASAP7_75t_L g4218 ( 
.A(n_3749),
.B(n_3751),
.Y(n_4218)
);

INVx4_ASAP7_75t_L g4219 ( 
.A(n_3657),
.Y(n_4219)
);

BUFx6f_ASAP7_75t_L g4220 ( 
.A(n_3883),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_3755),
.B(n_3088),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_3770),
.B(n_3326),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_3657),
.B(n_3294),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_3867),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_3867),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_3869),
.Y(n_4226)
);

CKINVDCx5p33_ASAP7_75t_R g4227 ( 
.A(n_3604),
.Y(n_4227)
);

INVx1_ASAP7_75t_L g4228 ( 
.A(n_3869),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_3770),
.B(n_3326),
.Y(n_4229)
);

HB1xp67_ASAP7_75t_L g4230 ( 
.A(n_3897),
.Y(n_4230)
);

AND2x2_ASAP7_75t_L g4231 ( 
.A(n_3896),
.B(n_3170),
.Y(n_4231)
);

AND2x4_ASAP7_75t_L g4232 ( 
.A(n_3707),
.B(n_3294),
.Y(n_4232)
);

BUFx3_ASAP7_75t_L g4233 ( 
.A(n_3876),
.Y(n_4233)
);

AND2x2_ASAP7_75t_L g4234 ( 
.A(n_3575),
.B(n_3170),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3586),
.B(n_3762),
.Y(n_4235)
);

BUFx3_ASAP7_75t_L g4236 ( 
.A(n_3876),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3875),
.Y(n_4237)
);

BUFx6f_ASAP7_75t_L g4238 ( 
.A(n_3898),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3758),
.B(n_3089),
.Y(n_4239)
);

BUFx12f_ASAP7_75t_SL g4240 ( 
.A(n_3902),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_SL g4241 ( 
.A(n_3628),
.B(n_3294),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_3762),
.Y(n_4242)
);

AND2x2_ASAP7_75t_L g4243 ( 
.A(n_3634),
.B(n_3171),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_L g4244 ( 
.A(n_3722),
.B(n_3089),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_3899),
.B(n_3176),
.Y(n_4245)
);

AND2x2_ASAP7_75t_SL g4246 ( 
.A(n_3844),
.B(n_3852),
.Y(n_4246)
);

INVxp67_ASAP7_75t_L g4247 ( 
.A(n_3687),
.Y(n_4247)
);

BUFx6f_ASAP7_75t_L g4248 ( 
.A(n_3733),
.Y(n_4248)
);

AND2x2_ASAP7_75t_L g4249 ( 
.A(n_3832),
.B(n_3839),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_3871),
.Y(n_4250)
);

BUFx3_ASAP7_75t_L g4251 ( 
.A(n_3733),
.Y(n_4251)
);

AND2x4_ASAP7_75t_L g4252 ( 
.A(n_3707),
.B(n_3295),
.Y(n_4252)
);

NOR2xp67_ASAP7_75t_L g4253 ( 
.A(n_3822),
.B(n_3353),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3848),
.B(n_3097),
.Y(n_4254)
);

BUFx8_ASAP7_75t_SL g4255 ( 
.A(n_3604),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_3873),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_3858),
.B(n_3176),
.Y(n_4257)
);

INVx3_ASAP7_75t_L g4258 ( 
.A(n_3892),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_3820),
.B(n_3177),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3826),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_3688),
.Y(n_4261)
);

INVx2_ASAP7_75t_L g4262 ( 
.A(n_3690),
.Y(n_4262)
);

OAI21xp5_ASAP7_75t_L g4263 ( 
.A1(n_3986),
.A2(n_3756),
.B(n_3643),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_4148),
.B(n_3866),
.Y(n_4264)
);

OAI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_3986),
.A2(n_3808),
.B(n_3653),
.Y(n_4265)
);

AND2x4_ASAP7_75t_L g4266 ( 
.A(n_4003),
.B(n_3748),
.Y(n_4266)
);

OAI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_4039),
.A2(n_3629),
.B(n_3311),
.Y(n_4267)
);

NAND3xp33_ASAP7_75t_L g4268 ( 
.A(n_3957),
.B(n_3752),
.C(n_3759),
.Y(n_4268)
);

A2O1A1Ixp33_ASAP7_75t_L g4269 ( 
.A1(n_4130),
.A2(n_3727),
.B(n_3620),
.C(n_3783),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_L g4270 ( 
.A(n_4148),
.B(n_3632),
.Y(n_4270)
);

AOI21xp5_ASAP7_75t_L g4271 ( 
.A1(n_4216),
.A2(n_3621),
.B(n_3670),
.Y(n_4271)
);

AOI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_4164),
.A2(n_3603),
.B(n_3636),
.Y(n_4272)
);

NAND3xp33_ASAP7_75t_SL g4273 ( 
.A(n_4052),
.B(n_3614),
.C(n_2469),
.Y(n_4273)
);

NAND2xp5_ASAP7_75t_L g4274 ( 
.A(n_3906),
.B(n_3803),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3966),
.B(n_3728),
.Y(n_4275)
);

NOR2x1p5_ASAP7_75t_SL g4276 ( 
.A(n_3939),
.B(n_2903),
.Y(n_4276)
);

INVxp67_ASAP7_75t_L g4277 ( 
.A(n_3983),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_3951),
.B(n_3807),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4127),
.B(n_3814),
.Y(n_4279)
);

NAND3xp33_ASAP7_75t_L g4280 ( 
.A(n_4122),
.B(n_779),
.C(n_775),
.Y(n_4280)
);

NAND2xp5_ASAP7_75t_L g4281 ( 
.A(n_4127),
.B(n_3818),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_3943),
.A2(n_3763),
.B(n_3506),
.Y(n_4282)
);

NAND2xp5_ASAP7_75t_L g4283 ( 
.A(n_3925),
.B(n_3894),
.Y(n_4283)
);

OAI21xp5_ASAP7_75t_L g4284 ( 
.A1(n_4247),
.A2(n_4082),
.B(n_4134),
.Y(n_4284)
);

AOI21xp5_ASAP7_75t_L g4285 ( 
.A1(n_3943),
.A2(n_3971),
.B(n_4081),
.Y(n_4285)
);

OAI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_3997),
.A2(n_3806),
.B1(n_3841),
.B2(n_3571),
.Y(n_4286)
);

NAND3xp33_ASAP7_75t_L g4287 ( 
.A(n_3976),
.B(n_782),
.C(n_779),
.Y(n_4287)
);

OAI22xp33_ASAP7_75t_L g4288 ( 
.A1(n_3997),
.A2(n_3571),
.B1(n_2665),
.B2(n_3518),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4033),
.Y(n_4289)
);

OAI22xp5_ASAP7_75t_L g4290 ( 
.A1(n_4130),
.A2(n_3571),
.B1(n_3613),
.B2(n_3861),
.Y(n_4290)
);

NOR2xp33_ASAP7_75t_L g4291 ( 
.A(n_4214),
.B(n_2414),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_3919),
.B(n_1041),
.Y(n_4292)
);

BUFx6f_ASAP7_75t_L g4293 ( 
.A(n_3920),
.Y(n_4293)
);

NAND3xp33_ASAP7_75t_L g4294 ( 
.A(n_4042),
.B(n_806),
.C(n_782),
.Y(n_4294)
);

AOI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_4108),
.A2(n_3514),
.B(n_3502),
.Y(n_4295)
);

AOI22xp5_ASAP7_75t_L g4296 ( 
.A1(n_4044),
.A2(n_3865),
.B1(n_2449),
.B2(n_2482),
.Y(n_4296)
);

AOI22xp33_ASAP7_75t_L g4297 ( 
.A1(n_4044),
.A2(n_3606),
.B1(n_2414),
.B2(n_2485),
.Y(n_4297)
);

OAI22xp5_ASAP7_75t_L g4298 ( 
.A1(n_4180),
.A2(n_3781),
.B1(n_3518),
.B2(n_2797),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_3967),
.B(n_1120),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_3905),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_SL g4301 ( 
.A(n_4004),
.B(n_3800),
.Y(n_4301)
);

BUFx4f_ASAP7_75t_L g4302 ( 
.A(n_3908),
.Y(n_4302)
);

NOR2xp33_ASAP7_75t_L g4303 ( 
.A(n_4214),
.B(n_2482),
.Y(n_4303)
);

BUFx6f_ASAP7_75t_L g4304 ( 
.A(n_3920),
.Y(n_4304)
);

AO22x1_ASAP7_75t_L g4305 ( 
.A1(n_4135),
.A2(n_2485),
.B1(n_3469),
.B2(n_3466),
.Y(n_4305)
);

OAI22xp5_ASAP7_75t_L g4306 ( 
.A1(n_4178),
.A2(n_3781),
.B1(n_2808),
.B2(n_2777),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4014),
.B(n_3311),
.Y(n_4307)
);

AOI21xp5_ASAP7_75t_L g4308 ( 
.A1(n_4108),
.A2(n_3529),
.B(n_3514),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4096),
.B(n_3311),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4072),
.A2(n_3540),
.B(n_3529),
.Y(n_4310)
);

NOR2xp67_ASAP7_75t_L g4311 ( 
.A(n_4026),
.B(n_3711),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_SL g4312 ( 
.A(n_4004),
.B(n_3712),
.Y(n_4312)
);

NAND3xp33_ASAP7_75t_L g4313 ( 
.A(n_4072),
.B(n_809),
.C(n_806),
.Y(n_4313)
);

AOI21xp5_ASAP7_75t_L g4314 ( 
.A1(n_4241),
.A2(n_3562),
.B(n_3559),
.Y(n_4314)
);

OAI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_4181),
.A2(n_2875),
.B(n_2854),
.Y(n_4315)
);

NAND2xp5_ASAP7_75t_SL g4316 ( 
.A(n_4213),
.B(n_3295),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4253),
.B(n_3295),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3947),
.B(n_3103),
.Y(n_4318)
);

AND2x4_ASAP7_75t_L g4319 ( 
.A(n_4003),
.B(n_4034),
.Y(n_4319)
);

O2A1O1Ixp33_ASAP7_75t_L g4320 ( 
.A1(n_4018),
.A2(n_2024),
.B(n_811),
.C(n_820),
.Y(n_4320)
);

AOI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_4099),
.A2(n_3540),
.B(n_3594),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_4095),
.A2(n_3117),
.B(n_3177),
.Y(n_4322)
);

INVx2_ASAP7_75t_L g4323 ( 
.A(n_3909),
.Y(n_4323)
);

O2A1O1Ixp33_ASAP7_75t_L g4324 ( 
.A1(n_4189),
.A2(n_811),
.B(n_820),
.C(n_810),
.Y(n_4324)
);

AO21x1_ASAP7_75t_L g4325 ( 
.A1(n_3930),
.A2(n_823),
.B(n_822),
.Y(n_4325)
);

AOI21x1_ASAP7_75t_L g4326 ( 
.A1(n_4128),
.A2(n_2885),
.B(n_2879),
.Y(n_4326)
);

AOI21xp33_ASAP7_75t_L g4327 ( 
.A1(n_4246),
.A2(n_3103),
.B(n_3645),
.Y(n_4327)
);

BUFx6f_ASAP7_75t_L g4328 ( 
.A(n_3934),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_3911),
.Y(n_4329)
);

O2A1O1Ixp33_ASAP7_75t_L g4330 ( 
.A1(n_4218),
.A2(n_823),
.B(n_825),
.C(n_822),
.Y(n_4330)
);

AOI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_3932),
.A2(n_3185),
.B(n_3669),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3975),
.B(n_2485),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_3912),
.Y(n_4333)
);

OAI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_3965),
.A2(n_3094),
.B(n_3173),
.Y(n_4334)
);

OAI22xp5_ASAP7_75t_L g4335 ( 
.A1(n_4201),
.A2(n_3159),
.B1(n_3151),
.B2(n_3121),
.Y(n_4335)
);

AND2x4_ASAP7_75t_SL g4336 ( 
.A(n_4088),
.B(n_3508),
.Y(n_4336)
);

AOI21xp5_ASAP7_75t_L g4337 ( 
.A1(n_3961),
.A2(n_3185),
.B(n_2823),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_3941),
.B(n_3306),
.Y(n_4338)
);

NOR2xp33_ASAP7_75t_L g4339 ( 
.A(n_4045),
.B(n_3716),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_3941),
.B(n_3306),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_4064),
.A2(n_2823),
.B(n_2798),
.Y(n_4341)
);

INVxp67_ASAP7_75t_L g4342 ( 
.A(n_4230),
.Y(n_4342)
);

INVx2_ASAP7_75t_L g4343 ( 
.A(n_4057),
.Y(n_4343)
);

NOR2xp33_ASAP7_75t_L g4344 ( 
.A(n_4203),
.B(n_3508),
.Y(n_4344)
);

INVx3_ASAP7_75t_L g4345 ( 
.A(n_4034),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3940),
.Y(n_4346)
);

INVx2_ASAP7_75t_SL g4347 ( 
.A(n_3934),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_4003),
.B(n_3375),
.Y(n_4348)
);

NOR2xp33_ASAP7_75t_L g4349 ( 
.A(n_4215),
.B(n_1468),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_4110),
.B(n_3321),
.Y(n_4350)
);

NOR2xp33_ASAP7_75t_L g4351 ( 
.A(n_4100),
.B(n_1472),
.Y(n_4351)
);

AOI21xp5_ASAP7_75t_L g4352 ( 
.A1(n_4071),
.A2(n_3110),
.B(n_3106),
.Y(n_4352)
);

NOR3xp33_ASAP7_75t_L g4353 ( 
.A(n_4028),
.B(n_826),
.C(n_825),
.Y(n_4353)
);

OAI22xp5_ASAP7_75t_L g4354 ( 
.A1(n_4182),
.A2(n_3122),
.B1(n_3144),
.B2(n_3123),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_4071),
.A2(n_3110),
.B(n_3106),
.Y(n_4355)
);

CKINVDCx10_ASAP7_75t_R g4356 ( 
.A(n_4255),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_L g4357 ( 
.A(n_4113),
.B(n_1472),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4116),
.B(n_1473),
.Y(n_4358)
);

AOI21xp5_ASAP7_75t_L g4359 ( 
.A1(n_4079),
.A2(n_3172),
.B(n_3175),
.Y(n_4359)
);

OAI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4166),
.A2(n_3127),
.B1(n_3130),
.B2(n_3084),
.Y(n_4360)
);

OAI21xp5_ASAP7_75t_L g4361 ( 
.A1(n_4195),
.A2(n_3198),
.B(n_3372),
.Y(n_4361)
);

O2A1O1Ixp33_ASAP7_75t_L g4362 ( 
.A1(n_4184),
.A2(n_827),
.B(n_828),
.C(n_826),
.Y(n_4362)
);

HB1xp67_ASAP7_75t_L g4363 ( 
.A(n_3960),
.Y(n_4363)
);

NAND2xp5_ASAP7_75t_SL g4364 ( 
.A(n_4246),
.B(n_4041),
.Y(n_4364)
);

OR2x6_ASAP7_75t_L g4365 ( 
.A(n_3948),
.B(n_3619),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_3931),
.B(n_1473),
.Y(n_4366)
);

AND2x4_ASAP7_75t_L g4367 ( 
.A(n_4060),
.B(n_3375),
.Y(n_4367)
);

OAI21xp33_ASAP7_75t_L g4368 ( 
.A1(n_3956),
.A2(n_838),
.B(n_831),
.Y(n_4368)
);

A2O1A1Ixp33_ASAP7_75t_L g4369 ( 
.A1(n_4056),
.A2(n_3547),
.B(n_2195),
.C(n_2204),
.Y(n_4369)
);

BUFx8_ASAP7_75t_L g4370 ( 
.A(n_3938),
.Y(n_4370)
);

AOI21xp5_ASAP7_75t_L g4371 ( 
.A1(n_4146),
.A2(n_3143),
.B(n_3140),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4065),
.Y(n_4372)
);

AOI21xp5_ASAP7_75t_L g4373 ( 
.A1(n_3944),
.A2(n_3143),
.B(n_3140),
.Y(n_4373)
);

AO21x1_ASAP7_75t_L g4374 ( 
.A1(n_3968),
.A2(n_3978),
.B(n_4119),
.Y(n_4374)
);

INVx3_ASAP7_75t_L g4375 ( 
.A(n_4060),
.Y(n_4375)
);

NAND2xp5_ASAP7_75t_L g4376 ( 
.A(n_4073),
.B(n_1475),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_3949),
.B(n_1475),
.Y(n_4377)
);

OAI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_4043),
.A2(n_3381),
.B(n_3372),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4160),
.B(n_1477),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_4124),
.B(n_4131),
.Y(n_4380)
);

AND2x4_ASAP7_75t_L g4381 ( 
.A(n_3955),
.B(n_3375),
.Y(n_4381)
);

OAI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_4206),
.A2(n_3381),
.B(n_3372),
.Y(n_4382)
);

AOI21x1_ASAP7_75t_L g4383 ( 
.A1(n_4254),
.A2(n_3125),
.B(n_3116),
.Y(n_4383)
);

AOI21xp5_ASAP7_75t_L g4384 ( 
.A1(n_3944),
.A2(n_3160),
.B(n_3158),
.Y(n_4384)
);

A2O1A1Ixp33_ASAP7_75t_L g4385 ( 
.A1(n_4163),
.A2(n_2195),
.B(n_2204),
.C(n_2160),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_4160),
.B(n_1477),
.Y(n_4386)
);

NOR2xp33_ASAP7_75t_L g4387 ( 
.A(n_4190),
.B(n_1478),
.Y(n_4387)
);

BUFx6f_ASAP7_75t_L g4388 ( 
.A(n_3938),
.Y(n_4388)
);

AND2x4_ASAP7_75t_L g4389 ( 
.A(n_3955),
.B(n_3378),
.Y(n_4389)
);

AOI21xp5_ASAP7_75t_L g4390 ( 
.A1(n_3944),
.A2(n_3160),
.B(n_3158),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_SL g4391 ( 
.A(n_4041),
.B(n_3378),
.Y(n_4391)
);

AOI21xp5_ASAP7_75t_L g4392 ( 
.A1(n_3944),
.A2(n_3166),
.B(n_3164),
.Y(n_4392)
);

AOI21xp5_ASAP7_75t_L g4393 ( 
.A1(n_3944),
.A2(n_3166),
.B(n_3164),
.Y(n_4393)
);

NOR2xp33_ASAP7_75t_L g4394 ( 
.A(n_4076),
.B(n_1478),
.Y(n_4394)
);

O2A1O1Ixp33_ASAP7_75t_L g4395 ( 
.A1(n_4142),
.A2(n_838),
.B(n_844),
.C(n_842),
.Y(n_4395)
);

AOI21xp33_ASAP7_75t_L g4396 ( 
.A1(n_4114),
.A2(n_2221),
.B(n_3186),
.Y(n_4396)
);

HB1xp67_ASAP7_75t_L g4397 ( 
.A(n_3960),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4046),
.B(n_1481),
.Y(n_4398)
);

AOI21xp5_ASAP7_75t_L g4399 ( 
.A1(n_4163),
.A2(n_3168),
.B(n_3183),
.Y(n_4399)
);

INVx4_ASAP7_75t_L g4400 ( 
.A(n_4202),
.Y(n_4400)
);

INVx3_ASAP7_75t_L g4401 ( 
.A(n_4219),
.Y(n_4401)
);

AOI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4061),
.A2(n_3168),
.B(n_3183),
.Y(n_4402)
);

NAND2xp5_ASAP7_75t_L g4403 ( 
.A(n_4047),
.B(n_1481),
.Y(n_4403)
);

O2A1O1Ixp33_ASAP7_75t_L g4404 ( 
.A1(n_4207),
.A2(n_840),
.B(n_858),
.C(n_844),
.Y(n_4404)
);

NOR2xp33_ASAP7_75t_SL g4405 ( 
.A(n_3936),
.B(n_3420),
.Y(n_4405)
);

INVx3_ASAP7_75t_L g4406 ( 
.A(n_4219),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_3927),
.B(n_1485),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4068),
.Y(n_4408)
);

INVx2_ASAP7_75t_L g4409 ( 
.A(n_4075),
.Y(n_4409)
);

A2O1A1Ixp33_ASAP7_75t_L g4410 ( 
.A1(n_4086),
.A2(n_2207),
.B(n_2204),
.C(n_842),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_3927),
.B(n_1485),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_SL g4412 ( 
.A(n_4041),
.B(n_3378),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4165),
.B(n_1486),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_L g4414 ( 
.A(n_4136),
.B(n_1486),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4077),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_3980),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4078),
.Y(n_4417)
);

INVxp67_ASAP7_75t_L g4418 ( 
.A(n_3950),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4140),
.B(n_3982),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_4244),
.B(n_1490),
.Y(n_4420)
);

O2A1O1Ixp33_ASAP7_75t_L g4421 ( 
.A1(n_4209),
.A2(n_840),
.B(n_867),
.C(n_856),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_3928),
.B(n_1490),
.Y(n_4422)
);

AOI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_3948),
.A2(n_4086),
.B(n_3959),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_3959),
.A2(n_3184),
.B(n_3161),
.Y(n_4424)
);

INVx3_ASAP7_75t_L g4425 ( 
.A(n_4219),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_3910),
.A2(n_4049),
.B(n_4085),
.Y(n_4426)
);

INVxp67_ASAP7_75t_L g4427 ( 
.A(n_4007),
.Y(n_4427)
);

AOI21xp5_ASAP7_75t_L g4428 ( 
.A1(n_3910),
.A2(n_3161),
.B(n_3345),
.Y(n_4428)
);

BUFx2_ASAP7_75t_L g4429 ( 
.A(n_4240),
.Y(n_4429)
);

INVx2_ASAP7_75t_L g4430 ( 
.A(n_4080),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4087),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_L g4432 ( 
.A(n_3928),
.B(n_1495),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_L g4433 ( 
.A(n_3963),
.B(n_1495),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_3963),
.B(n_1496),
.Y(n_4434)
);

BUFx6f_ASAP7_75t_L g4435 ( 
.A(n_4022),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4097),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_3969),
.B(n_1496),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4137),
.B(n_856),
.Y(n_4438)
);

AND2x6_ASAP7_75t_L g4439 ( 
.A(n_4217),
.B(n_3393),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_L g4440 ( 
.A(n_3969),
.B(n_1497),
.Y(n_4440)
);

AOI22xp5_ASAP7_75t_L g4441 ( 
.A1(n_3958),
.A2(n_3469),
.B1(n_3381),
.B2(n_3372),
.Y(n_4441)
);

INVx3_ASAP7_75t_L g4442 ( 
.A(n_3935),
.Y(n_4442)
);

AOI21xp5_ASAP7_75t_L g4443 ( 
.A1(n_4049),
.A2(n_4090),
.B(n_4085),
.Y(n_4443)
);

AOI21xp5_ASAP7_75t_L g4444 ( 
.A1(n_4049),
.A2(n_3515),
.B(n_3477),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_3973),
.B(n_1497),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_3973),
.B(n_1498),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_3981),
.B(n_1498),
.Y(n_4447)
);

OR2x2_ASAP7_75t_L g4448 ( 
.A(n_4105),
.B(n_858),
.Y(n_4448)
);

OAI22xp5_ASAP7_75t_L g4449 ( 
.A1(n_3977),
.A2(n_1504),
.B1(n_1509),
.B2(n_1501),
.Y(n_4449)
);

O2A1O1Ixp33_ASAP7_75t_L g4450 ( 
.A1(n_4221),
.A2(n_869),
.B(n_870),
.C(n_867),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_L g4451 ( 
.A(n_3981),
.B(n_1501),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_3984),
.B(n_1504),
.Y(n_4452)
);

AOI22xp5_ASAP7_75t_L g4453 ( 
.A1(n_3958),
.A2(n_3469),
.B1(n_3381),
.B2(n_2207),
.Y(n_4453)
);

O2A1O1Ixp33_ASAP7_75t_L g4454 ( 
.A1(n_4239),
.A2(n_870),
.B(n_880),
.C(n_869),
.Y(n_4454)
);

AO32x2_ASAP7_75t_L g4455 ( 
.A1(n_3954),
.A2(n_2996),
.A3(n_2999),
.B1(n_2991),
.B2(n_2979),
.Y(n_4455)
);

CKINVDCx5p33_ASAP7_75t_R g4456 ( 
.A(n_4255),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_L g4457 ( 
.A(n_3990),
.B(n_1515),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_L g4458 ( 
.A(n_3990),
.B(n_1516),
.Y(n_4458)
);

OAI22xp5_ASAP7_75t_L g4459 ( 
.A1(n_4089),
.A2(n_4227),
.B1(n_4199),
.B2(n_3985),
.Y(n_4459)
);

OAI22xp5_ASAP7_75t_L g4460 ( 
.A1(n_4227),
.A2(n_1520),
.B1(n_1523),
.B2(n_1519),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_3993),
.B(n_1520),
.Y(n_4461)
);

AOI21xp5_ASAP7_75t_L g4462 ( 
.A1(n_4090),
.A2(n_3071),
.B(n_3044),
.Y(n_4462)
);

AOI21xp5_ASAP7_75t_L g4463 ( 
.A1(n_4139),
.A2(n_3087),
.B(n_3071),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4009),
.Y(n_4464)
);

NAND2xp5_ASAP7_75t_L g4465 ( 
.A(n_3993),
.B(n_1523),
.Y(n_4465)
);

OR2x6_ASAP7_75t_SL g4466 ( 
.A(n_4173),
.B(n_848),
.Y(n_4466)
);

AOI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_4139),
.A2(n_3087),
.B(n_3071),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_L g4468 ( 
.A(n_3995),
.B(n_1529),
.Y(n_4468)
);

NAND3xp33_ASAP7_75t_L g4469 ( 
.A(n_4260),
.B(n_889),
.C(n_880),
.Y(n_4469)
);

NOR3xp33_ASAP7_75t_L g4470 ( 
.A(n_4176),
.B(n_898),
.C(n_889),
.Y(n_4470)
);

INVx3_ASAP7_75t_L g4471 ( 
.A(n_3935),
.Y(n_4471)
);

OAI22xp5_ASAP7_75t_L g4472 ( 
.A1(n_4069),
.A2(n_1531),
.B1(n_1533),
.B2(n_1529),
.Y(n_4472)
);

AOI21xp5_ASAP7_75t_L g4473 ( 
.A1(n_4152),
.A2(n_3974),
.B(n_3970),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4098),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_SL g4475 ( 
.A(n_4152),
.B(n_3393),
.Y(n_4475)
);

BUFx6f_ASAP7_75t_L g4476 ( 
.A(n_4022),
.Y(n_4476)
);

O2A1O1Ixp33_ASAP7_75t_L g4477 ( 
.A1(n_4154),
.A2(n_912),
.B(n_915),
.C(n_900),
.Y(n_4477)
);

O2A1O1Ixp33_ASAP7_75t_L g4478 ( 
.A1(n_4091),
.A2(n_912),
.B(n_915),
.C(n_910),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4138),
.B(n_910),
.Y(n_4479)
);

INVx2_ASAP7_75t_L g4480 ( 
.A(n_3907),
.Y(n_4480)
);

OAI21xp5_ASAP7_75t_L g4481 ( 
.A1(n_4256),
.A2(n_2061),
.B(n_1985),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4098),
.Y(n_4482)
);

O2A1O1Ixp33_ASAP7_75t_L g4483 ( 
.A1(n_3953),
.A2(n_923),
.B(n_924),
.C(n_921),
.Y(n_4483)
);

O2A1O1Ixp33_ASAP7_75t_L g4484 ( 
.A1(n_4204),
.A2(n_923),
.B(n_924),
.C(n_921),
.Y(n_4484)
);

NOR2xp33_ASAP7_75t_L g4485 ( 
.A(n_3945),
.B(n_1533),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_L g4486 ( 
.A(n_4001),
.B(n_1535),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_4012),
.B(n_1535),
.Y(n_4487)
);

NOR2xp33_ASAP7_75t_L g4488 ( 
.A(n_3945),
.B(n_1537),
.Y(n_4488)
);

AOI21xp5_ASAP7_75t_L g4489 ( 
.A1(n_3970),
.A2(n_3099),
.B(n_3096),
.Y(n_4489)
);

O2A1O1Ixp33_ASAP7_75t_L g4490 ( 
.A1(n_3979),
.A2(n_939),
.B(n_944),
.C(n_925),
.Y(n_4490)
);

AOI22xp33_ASAP7_75t_L g4491 ( 
.A1(n_4138),
.A2(n_2177),
.B1(n_2179),
.B2(n_2169),
.Y(n_4491)
);

INVx1_ASAP7_75t_L g4492 ( 
.A(n_4102),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_SL g4493 ( 
.A(n_3939),
.B(n_3393),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_4012),
.B(n_1537),
.Y(n_4494)
);

OAI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_3917),
.A2(n_3333),
.B(n_3297),
.Y(n_4495)
);

NOR2xp33_ASAP7_75t_L g4496 ( 
.A(n_3972),
.B(n_1542),
.Y(n_4496)
);

AOI21xp5_ASAP7_75t_L g4497 ( 
.A1(n_3970),
.A2(n_3099),
.B(n_3096),
.Y(n_4497)
);

AOI21xp5_ASAP7_75t_L g4498 ( 
.A1(n_3970),
.A2(n_3946),
.B(n_3935),
.Y(n_4498)
);

O2A1O1Ixp33_ASAP7_75t_L g4499 ( 
.A1(n_3991),
.A2(n_939),
.B(n_944),
.C(n_925),
.Y(n_4499)
);

AOI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4059),
.A2(n_2207),
.B1(n_2204),
.B2(n_2134),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4015),
.B(n_4020),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_L g4502 ( 
.A(n_4015),
.B(n_1544),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4102),
.Y(n_4503)
);

AOI21xp5_ASAP7_75t_L g4504 ( 
.A1(n_3946),
.A2(n_3099),
.B(n_3096),
.Y(n_4504)
);

NOR2xp33_ASAP7_75t_L g4505 ( 
.A(n_3972),
.B(n_1545),
.Y(n_4505)
);

BUFx4f_ASAP7_75t_L g4506 ( 
.A(n_3908),
.Y(n_4506)
);

AOI21xp5_ASAP7_75t_L g4507 ( 
.A1(n_3946),
.A2(n_3132),
.B(n_3099),
.Y(n_4507)
);

AOI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4186),
.A2(n_3132),
.B(n_3099),
.Y(n_4508)
);

AOI22xp5_ASAP7_75t_L g4509 ( 
.A1(n_4059),
.A2(n_2207),
.B1(n_2134),
.B2(n_2143),
.Y(n_4509)
);

INVx5_ASAP7_75t_L g4510 ( 
.A(n_3942),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4020),
.B(n_1547),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_L g4512 ( 
.A(n_4024),
.B(n_1547),
.Y(n_4512)
);

BUFx2_ASAP7_75t_SL g4513 ( 
.A(n_4194),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4024),
.B(n_1548),
.Y(n_4514)
);

O2A1O1Ixp5_ASAP7_75t_L g4515 ( 
.A1(n_3913),
.A2(n_2847),
.B(n_2891),
.C(n_2842),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4025),
.B(n_1548),
.Y(n_4516)
);

BUFx6f_ASAP7_75t_L g4517 ( 
.A(n_4022),
.Y(n_4517)
);

O2A1O1Ixp33_ASAP7_75t_L g4518 ( 
.A1(n_3991),
.A2(n_948),
.B(n_950),
.C(n_946),
.Y(n_4518)
);

AOI21xp5_ASAP7_75t_L g4519 ( 
.A1(n_4208),
.A2(n_3619),
.B(n_3430),
.Y(n_4519)
);

NAND2x1p5_ASAP7_75t_L g4520 ( 
.A(n_3936),
.B(n_3420),
.Y(n_4520)
);

AOI21xp5_ASAP7_75t_L g4521 ( 
.A1(n_4208),
.A2(n_3430),
.B(n_3411),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_3987),
.A2(n_3430),
.B(n_3411),
.Y(n_4522)
);

O2A1O1Ixp33_ASAP7_75t_L g4523 ( 
.A1(n_3994),
.A2(n_948),
.B(n_950),
.C(n_946),
.Y(n_4523)
);

AOI21x1_ASAP7_75t_L g4524 ( 
.A1(n_4250),
.A2(n_3126),
.B(n_3178),
.Y(n_4524)
);

OAI22xp5_ASAP7_75t_L g4525 ( 
.A1(n_3994),
.A2(n_1558),
.B1(n_1561),
.B2(n_1549),
.Y(n_4525)
);

O2A1O1Ixp33_ASAP7_75t_L g4526 ( 
.A1(n_4170),
.A2(n_954),
.B(n_956),
.C(n_951),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_3987),
.A2(n_3411),
.B(n_3503),
.Y(n_4527)
);

OAI22xp5_ASAP7_75t_L g4528 ( 
.A1(n_4257),
.A2(n_1558),
.B1(n_1563),
.B2(n_1549),
.Y(n_4528)
);

CKINVDCx6p67_ASAP7_75t_R g4529 ( 
.A(n_4202),
.Y(n_4529)
);

OAI321xp33_ASAP7_75t_L g4530 ( 
.A1(n_3914),
.A2(n_959),
.A3(n_954),
.B1(n_961),
.B2(n_956),
.C(n_951),
.Y(n_4530)
);

INVx1_ASAP7_75t_L g4531 ( 
.A(n_4121),
.Y(n_4531)
);

O2A1O1Ixp33_ASAP7_75t_L g4532 ( 
.A1(n_4170),
.A2(n_961),
.B(n_967),
.C(n_959),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4025),
.B(n_1563),
.Y(n_4533)
);

BUFx4f_ASAP7_75t_L g4534 ( 
.A(n_3908),
.Y(n_4534)
);

NAND3xp33_ASAP7_75t_L g4535 ( 
.A(n_4027),
.B(n_967),
.C(n_963),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_SL g4536 ( 
.A(n_3939),
.B(n_3503),
.Y(n_4536)
);

NOR2xp33_ASAP7_75t_L g4537 ( 
.A(n_4240),
.B(n_1567),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_4005),
.A2(n_3528),
.B(n_3567),
.Y(n_4538)
);

AND2x2_ASAP7_75t_L g4539 ( 
.A(n_4155),
.B(n_963),
.Y(n_4539)
);

INVx2_ASAP7_75t_SL g4540 ( 
.A(n_4022),
.Y(n_4540)
);

A2O1A1Ixp33_ASAP7_75t_L g4541 ( 
.A1(n_3914),
.A2(n_976),
.B(n_979),
.C(n_969),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4029),
.B(n_1569),
.Y(n_4542)
);

NOR2xp33_ASAP7_75t_L g4543 ( 
.A(n_4159),
.B(n_1569),
.Y(n_4543)
);

AOI21xp5_ASAP7_75t_L g4544 ( 
.A1(n_4222),
.A2(n_3568),
.B(n_3567),
.Y(n_4544)
);

AOI22xp33_ASAP7_75t_L g4545 ( 
.A1(n_4105),
.A2(n_2179),
.B1(n_2180),
.B2(n_2177),
.Y(n_4545)
);

AOI21xp5_ASAP7_75t_L g4546 ( 
.A1(n_4229),
.A2(n_3568),
.B(n_3462),
.Y(n_4546)
);

OA22x2_ASAP7_75t_L g4547 ( 
.A1(n_4002),
.A2(n_2134),
.B1(n_2143),
.B2(n_2101),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4031),
.B(n_969),
.Y(n_4548)
);

OA22x2_ASAP7_75t_L g4549 ( 
.A1(n_4187),
.A2(n_2143),
.B1(n_2149),
.B2(n_2101),
.Y(n_4549)
);

AO22x1_ASAP7_75t_L g4550 ( 
.A1(n_4059),
.A2(n_3462),
.B1(n_3548),
.B2(n_3536),
.Y(n_4550)
);

INVx3_ASAP7_75t_L g4551 ( 
.A(n_4202),
.Y(n_4551)
);

AOI21xp5_ASAP7_75t_L g4552 ( 
.A1(n_4229),
.A2(n_3568),
.B(n_3462),
.Y(n_4552)
);

BUFx3_ASAP7_75t_L g4553 ( 
.A(n_4067),
.Y(n_4553)
);

AND2x2_ASAP7_75t_L g4554 ( 
.A(n_4032),
.B(n_976),
.Y(n_4554)
);

OAI21xp5_ASAP7_75t_L g4555 ( 
.A1(n_3917),
.A2(n_2061),
.B(n_1985),
.Y(n_4555)
);

INVx4_ASAP7_75t_L g4556 ( 
.A(n_4202),
.Y(n_4556)
);

OAI22xp5_ASAP7_75t_L g4557 ( 
.A1(n_4257),
.A2(n_3333),
.B1(n_3297),
.B2(n_3536),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_SL g4558 ( 
.A(n_3939),
.B(n_3195),
.Y(n_4558)
);

INVx3_ASAP7_75t_L g4559 ( 
.A(n_4177),
.Y(n_4559)
);

AOI21xp5_ASAP7_75t_L g4560 ( 
.A1(n_3916),
.A2(n_3462),
.B(n_3420),
.Y(n_4560)
);

AO32x1_ASAP7_75t_L g4561 ( 
.A1(n_4107),
.A2(n_3181),
.A3(n_3179),
.B1(n_2781),
.B2(n_2919),
.Y(n_4561)
);

AOI21xp5_ASAP7_75t_L g4562 ( 
.A1(n_3916),
.A2(n_3536),
.B(n_3420),
.Y(n_4562)
);

BUFx4f_ASAP7_75t_L g4563 ( 
.A(n_3908),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_4032),
.B(n_979),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4037),
.B(n_982),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_3922),
.Y(n_4566)
);

OAI21xp33_ASAP7_75t_L g4567 ( 
.A1(n_3918),
.A2(n_985),
.B(n_982),
.Y(n_4567)
);

AOI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_3921),
.A2(n_3548),
.B(n_2971),
.Y(n_4568)
);

INVx11_ASAP7_75t_L g4569 ( 
.A(n_4059),
.Y(n_4569)
);

O2A1O1Ixp33_ASAP7_75t_SL g4570 ( 
.A1(n_4258),
.A2(n_991),
.B(n_992),
.C(n_985),
.Y(n_4570)
);

INVx1_ASAP7_75t_SL g4571 ( 
.A(n_4197),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4123),
.Y(n_4572)
);

OAI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_3918),
.A2(n_1004),
.B(n_997),
.Y(n_4573)
);

O2A1O1Ixp33_ASAP7_75t_L g4574 ( 
.A1(n_3933),
.A2(n_1004),
.B(n_1005),
.C(n_997),
.Y(n_4574)
);

NOR2xp33_ASAP7_75t_L g4575 ( 
.A(n_4067),
.B(n_849),
.Y(n_4575)
);

NOR2xp33_ASAP7_75t_L g4576 ( 
.A(n_4067),
.B(n_851),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_3924),
.Y(n_4577)
);

NOR2x1_ASAP7_75t_L g4578 ( 
.A(n_4177),
.B(n_3257),
.Y(n_4578)
);

OAI21xp33_ASAP7_75t_SL g4579 ( 
.A1(n_4177),
.A2(n_1006),
.B(n_1005),
.Y(n_4579)
);

OR2x6_ASAP7_75t_L g4580 ( 
.A(n_3954),
.B(n_4066),
.Y(n_4580)
);

AOI21xp5_ASAP7_75t_L g4581 ( 
.A1(n_3933),
.A2(n_3548),
.B(n_2971),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_SL g4582 ( 
.A(n_3939),
.B(n_3257),
.Y(n_4582)
);

AO21x1_ASAP7_75t_L g4583 ( 
.A1(n_4101),
.A2(n_1008),
.B(n_1006),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_3936),
.A2(n_2972),
.B(n_2969),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_3926),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4200),
.B(n_1011),
.Y(n_4586)
);

BUFx6f_ASAP7_75t_L g4587 ( 
.A(n_4067),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4125),
.A2(n_2972),
.B(n_2969),
.Y(n_4588)
);

INVx2_ASAP7_75t_SL g4589 ( 
.A(n_3996),
.Y(n_4589)
);

HB1xp67_ASAP7_75t_L g4590 ( 
.A(n_4234),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4205),
.B(n_1015),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_SL g4592 ( 
.A(n_3939),
.B(n_3942),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4224),
.B(n_4225),
.Y(n_4593)
);

INVx2_ASAP7_75t_L g4594 ( 
.A(n_3926),
.Y(n_4594)
);

AOI21xp5_ASAP7_75t_L g4595 ( 
.A1(n_4126),
.A2(n_2980),
.B(n_2976),
.Y(n_4595)
);

AOI22xp5_ASAP7_75t_L g4596 ( 
.A1(n_4193),
.A2(n_2101),
.B1(n_2151),
.B2(n_2149),
.Y(n_4596)
);

BUFx3_ASAP7_75t_L g4597 ( 
.A(n_4370),
.Y(n_4597)
);

OAI22x1_ASAP7_75t_L g4598 ( 
.A1(n_4296),
.A2(n_4193),
.B1(n_4212),
.B2(n_4107),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4419),
.B(n_4235),
.Y(n_4599)
);

NOR2xp67_ASAP7_75t_L g4600 ( 
.A(n_4339),
.B(n_3954),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4264),
.B(n_4235),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4342),
.B(n_4245),
.Y(n_4602)
);

A2O1A1Ixp33_ASAP7_75t_L g4603 ( 
.A1(n_4269),
.A2(n_4115),
.B(n_1036),
.C(n_1045),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_L g4604 ( 
.A(n_4277),
.B(n_4245),
.Y(n_4604)
);

AOI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_4265),
.A2(n_4017),
.B(n_4011),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_SL g4606 ( 
.A(n_4265),
.B(n_3942),
.Y(n_4606)
);

AND2x6_ASAP7_75t_L g4607 ( 
.A(n_4319),
.B(n_3952),
.Y(n_4607)
);

INVx5_ASAP7_75t_L g4608 ( 
.A(n_4293),
.Y(n_4608)
);

INVx1_ASAP7_75t_SL g4609 ( 
.A(n_4571),
.Y(n_4609)
);

AOI22xp33_ASAP7_75t_L g4610 ( 
.A1(n_4273),
.A2(n_4162),
.B1(n_4074),
.B2(n_4115),
.Y(n_4610)
);

NOR2xp33_ASAP7_75t_R g4611 ( 
.A(n_4456),
.B(n_4233),
.Y(n_4611)
);

INVx1_ASAP7_75t_SL g4612 ( 
.A(n_4571),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4363),
.B(n_4397),
.Y(n_4613)
);

AOI21xp5_ASAP7_75t_L g4614 ( 
.A1(n_4263),
.A2(n_4070),
.B(n_4058),
.Y(n_4614)
);

INVx2_ASAP7_75t_L g4615 ( 
.A(n_4300),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4289),
.Y(n_4616)
);

AND2x2_ASAP7_75t_SL g4617 ( 
.A(n_4429),
.B(n_4066),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4284),
.B(n_4228),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_SL g4619 ( 
.A(n_4293),
.B(n_3942),
.Y(n_4619)
);

OAI22xp5_ASAP7_75t_L g4620 ( 
.A1(n_4268),
.A2(n_4251),
.B1(n_4236),
.B2(n_4233),
.Y(n_4620)
);

INVxp67_ASAP7_75t_L g4621 ( 
.A(n_4283),
.Y(n_4621)
);

NOR3xp33_ASAP7_75t_SL g4622 ( 
.A(n_4351),
.B(n_854),
.C(n_853),
.Y(n_4622)
);

INVx4_ASAP7_75t_L g4623 ( 
.A(n_4293),
.Y(n_4623)
);

AOI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4263),
.A2(n_4070),
.B(n_4058),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_SL g4625 ( 
.A(n_4304),
.B(n_3939),
.Y(n_4625)
);

BUFx6f_ASAP7_75t_L g4626 ( 
.A(n_4304),
.Y(n_4626)
);

AOI21x1_ASAP7_75t_L g4627 ( 
.A1(n_4325),
.A2(n_4252),
.B(n_4232),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4323),
.Y(n_4628)
);

NOR2xp33_ASAP7_75t_L g4629 ( 
.A(n_4380),
.B(n_7),
.Y(n_4629)
);

AOI21xp5_ASAP7_75t_L g4630 ( 
.A1(n_4287),
.A2(n_4070),
.B(n_4058),
.Y(n_4630)
);

OR2x4_ASAP7_75t_L g4631 ( 
.A(n_4304),
.B(n_3923),
.Y(n_4631)
);

NAND3xp33_ASAP7_75t_L g4632 ( 
.A(n_4353),
.B(n_1036),
.C(n_1015),
.Y(n_4632)
);

AOI21xp5_ASAP7_75t_L g4633 ( 
.A1(n_4287),
.A2(n_4313),
.B(n_4592),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4329),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_SL g4635 ( 
.A(n_4328),
.B(n_4223),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4554),
.B(n_4050),
.Y(n_4636)
);

O2A1O1Ixp33_ASAP7_75t_L g4637 ( 
.A1(n_4267),
.A2(n_1051),
.B(n_1057),
.C(n_1045),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4333),
.Y(n_4638)
);

OR2x2_ASAP7_75t_L g4639 ( 
.A(n_4590),
.B(n_3915),
.Y(n_4639)
);

INVx1_ASAP7_75t_L g4640 ( 
.A(n_4346),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4343),
.Y(n_4641)
);

INVx2_ASAP7_75t_L g4642 ( 
.A(n_4372),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4408),
.Y(n_4643)
);

AOI21xp5_ASAP7_75t_L g4644 ( 
.A1(n_4294),
.A2(n_4132),
.B(n_4120),
.Y(n_4644)
);

NAND2xp5_ASAP7_75t_SL g4645 ( 
.A(n_4328),
.B(n_4223),
.Y(n_4645)
);

INVx3_ASAP7_75t_L g4646 ( 
.A(n_4328),
.Y(n_4646)
);

NAND2x1p5_ASAP7_75t_L g4647 ( 
.A(n_4510),
.B(n_4316),
.Y(n_4647)
);

OAI21xp33_ASAP7_75t_SL g4648 ( 
.A1(n_4569),
.A2(n_3988),
.B(n_3964),
.Y(n_4648)
);

NOR2xp33_ASAP7_75t_L g4649 ( 
.A(n_4387),
.B(n_8),
.Y(n_4649)
);

O2A1O1Ixp33_ASAP7_75t_L g4650 ( 
.A1(n_4267),
.A2(n_1057),
.B(n_1068),
.C(n_1051),
.Y(n_4650)
);

A2O1A1Ixp33_ASAP7_75t_L g4651 ( 
.A1(n_4324),
.A2(n_1076),
.B(n_1085),
.C(n_1068),
.Y(n_4651)
);

O2A1O1Ixp33_ASAP7_75t_L g4652 ( 
.A1(n_4330),
.A2(n_1085),
.B(n_1090),
.C(n_1076),
.Y(n_4652)
);

AOI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_4271),
.A2(n_4153),
.B(n_4171),
.Y(n_4653)
);

OR2x2_ASAP7_75t_L g4654 ( 
.A(n_4501),
.B(n_3915),
.Y(n_4654)
);

CKINVDCx5p33_ASAP7_75t_R g4655 ( 
.A(n_4356),
.Y(n_4655)
);

AOI22xp5_ASAP7_75t_L g4656 ( 
.A1(n_4290),
.A2(n_4249),
.B1(n_4248),
.B2(n_4112),
.Y(n_4656)
);

NOR2xp33_ASAP7_75t_R g4657 ( 
.A(n_4370),
.B(n_4106),
.Y(n_4657)
);

NOR2xp67_ASAP7_75t_L g4658 ( 
.A(n_4459),
.B(n_3999),
.Y(n_4658)
);

CKINVDCx5p33_ASAP7_75t_R g4659 ( 
.A(n_4336),
.Y(n_4659)
);

OAI22xp5_ASAP7_75t_L g4660 ( 
.A1(n_4280),
.A2(n_4106),
.B1(n_1090),
.B2(n_1101),
.Y(n_4660)
);

A2O1A1Ixp33_ASAP7_75t_L g4661 ( 
.A1(n_4395),
.A2(n_1101),
.B(n_1103),
.C(n_1094),
.Y(n_4661)
);

OAI21x1_ASAP7_75t_L g4662 ( 
.A1(n_4322),
.A2(n_4153),
.B(n_4084),
.Y(n_4662)
);

AOI21x1_ASAP7_75t_L g4663 ( 
.A1(n_4374),
.A2(n_4591),
.B(n_4586),
.Y(n_4663)
);

AOI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4428),
.A2(n_4175),
.B(n_4171),
.Y(n_4664)
);

BUFx6f_ASAP7_75t_L g4665 ( 
.A(n_4388),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4479),
.B(n_4231),
.Y(n_4666)
);

O2A1O1Ixp33_ASAP7_75t_SL g4667 ( 
.A1(n_4349),
.A2(n_1103),
.B(n_1105),
.C(n_1094),
.Y(n_4667)
);

NAND2xp5_ASAP7_75t_SL g4668 ( 
.A(n_4388),
.B(n_4223),
.Y(n_4668)
);

INVx2_ASAP7_75t_SL g4669 ( 
.A(n_4347),
.Y(n_4669)
);

AND2x4_ASAP7_75t_L g4670 ( 
.A(n_4442),
.B(n_3952),
.Y(n_4670)
);

BUFx6f_ASAP7_75t_L g4671 ( 
.A(n_4435),
.Y(n_4671)
);

INVx1_ASAP7_75t_L g4672 ( 
.A(n_4416),
.Y(n_4672)
);

BUFx3_ASAP7_75t_L g4673 ( 
.A(n_4553),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4270),
.B(n_4104),
.Y(n_4674)
);

NOR2xp33_ASAP7_75t_L g4675 ( 
.A(n_4485),
.B(n_8),
.Y(n_4675)
);

OAI22xp5_ASAP7_75t_L g4676 ( 
.A1(n_4385),
.A2(n_4248),
.B1(n_3923),
.B2(n_3952),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4427),
.B(n_4109),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_SL g4678 ( 
.A(n_4311),
.B(n_4232),
.Y(n_4678)
);

NOR2xp33_ASAP7_75t_L g4679 ( 
.A(n_4488),
.B(n_9),
.Y(n_4679)
);

NOR2xp33_ASAP7_75t_L g4680 ( 
.A(n_4496),
.B(n_10),
.Y(n_4680)
);

AOI22xp5_ASAP7_75t_L g4681 ( 
.A1(n_4280),
.A2(n_4249),
.B1(n_4248),
.B2(n_3952),
.Y(n_4681)
);

OR2x6_ASAP7_75t_L g4682 ( 
.A(n_4423),
.B(n_4117),
.Y(n_4682)
);

O2A1O1Ixp5_ASAP7_75t_L g4683 ( 
.A1(n_4364),
.A2(n_1112),
.B(n_1117),
.C(n_1105),
.Y(n_4683)
);

INVx2_ASAP7_75t_L g4684 ( 
.A(n_4409),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4415),
.Y(n_4685)
);

INVx2_ASAP7_75t_L g4686 ( 
.A(n_4417),
.Y(n_4686)
);

OAI22xp5_ASAP7_75t_L g4687 ( 
.A1(n_4500),
.A2(n_4248),
.B1(n_3923),
.B2(n_4129),
.Y(n_4687)
);

BUFx3_ASAP7_75t_L g4688 ( 
.A(n_4394),
.Y(n_4688)
);

A2O1A1Ixp33_ASAP7_75t_SL g4689 ( 
.A1(n_4505),
.A2(n_1117),
.B(n_1118),
.C(n_1112),
.Y(n_4689)
);

O2A1O1Ixp33_ASAP7_75t_L g4690 ( 
.A1(n_4362),
.A2(n_1118),
.B(n_2183),
.C(n_2180),
.Y(n_4690)
);

NOR2xp33_ASAP7_75t_L g4691 ( 
.A(n_4418),
.B(n_11),
.Y(n_4691)
);

AOI21xp5_ASAP7_75t_L g4692 ( 
.A1(n_4337),
.A2(n_4000),
.B(n_3999),
.Y(n_4692)
);

OAI22xp5_ASAP7_75t_L g4693 ( 
.A1(n_4509),
.A2(n_3923),
.B1(n_4129),
.B2(n_4117),
.Y(n_4693)
);

AOI22xp5_ASAP7_75t_L g4694 ( 
.A1(n_4470),
.A2(n_4243),
.B1(n_4053),
.B2(n_4054),
.Y(n_4694)
);

O2A1O1Ixp33_ASAP7_75t_L g4695 ( 
.A1(n_4320),
.A2(n_2186),
.B(n_2188),
.C(n_2183),
.Y(n_4695)
);

BUFx12f_ASAP7_75t_L g4696 ( 
.A(n_4448),
.Y(n_4696)
);

AOI21xp5_ASAP7_75t_L g4697 ( 
.A1(n_4314),
.A2(n_4030),
.B(n_4010),
.Y(n_4697)
);

INVx3_ASAP7_75t_L g4698 ( 
.A(n_4345),
.Y(n_4698)
);

BUFx6f_ASAP7_75t_L g4699 ( 
.A(n_4435),
.Y(n_4699)
);

NOR2xp33_ASAP7_75t_L g4700 ( 
.A(n_4379),
.B(n_11),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_4338),
.B(n_4111),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_SL g4702 ( 
.A(n_4285),
.B(n_4232),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_SL g4703 ( 
.A(n_4266),
.B(n_4426),
.Y(n_4703)
);

OAI22xp5_ASAP7_75t_L g4704 ( 
.A1(n_4410),
.A2(n_4369),
.B1(n_4466),
.B2(n_4297),
.Y(n_4704)
);

NOR2xp33_ASAP7_75t_SL g4705 ( 
.A(n_4510),
.B(n_4117),
.Y(n_4705)
);

A2O1A1Ixp33_ASAP7_75t_L g4706 ( 
.A1(n_4404),
.A2(n_4187),
.B(n_4053),
.C(n_4054),
.Y(n_4706)
);

AOI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4310),
.A2(n_4151),
.B(n_4144),
.Y(n_4707)
);

BUFx2_ASAP7_75t_L g4708 ( 
.A(n_4345),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4340),
.B(n_4350),
.Y(n_4709)
);

AOI22x1_ASAP7_75t_L g4710 ( 
.A1(n_4513),
.A2(n_857),
.B1(n_860),
.B2(n_855),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4464),
.Y(n_4711)
);

AND2x4_ASAP7_75t_L g4712 ( 
.A(n_4471),
.B(n_4129),
.Y(n_4712)
);

A2O1A1Ixp33_ASAP7_75t_L g4713 ( 
.A1(n_4421),
.A2(n_4051),
.B(n_4259),
.C(n_4141),
.Y(n_4713)
);

OAI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4535),
.A2(n_4016),
.B1(n_3998),
.B2(n_4118),
.Y(n_4714)
);

NOR2xp33_ASAP7_75t_L g4715 ( 
.A(n_4386),
.B(n_12),
.Y(n_4715)
);

AOI21xp5_ASAP7_75t_L g4716 ( 
.A1(n_4493),
.A2(n_4151),
.B(n_4144),
.Y(n_4716)
);

NAND2xp5_ASAP7_75t_SL g4717 ( 
.A(n_4435),
.B(n_4157),
.Y(n_4717)
);

A2O1A1Ixp33_ASAP7_75t_SL g4718 ( 
.A1(n_4344),
.A2(n_2188),
.B(n_2198),
.C(n_2186),
.Y(n_4718)
);

BUFx6f_ASAP7_75t_L g4719 ( 
.A(n_4476),
.Y(n_4719)
);

NOR2xp33_ASAP7_75t_L g4720 ( 
.A(n_4537),
.B(n_13),
.Y(n_4720)
);

CKINVDCx5p33_ASAP7_75t_R g4721 ( 
.A(n_4275),
.Y(n_4721)
);

NOR2xp33_ASAP7_75t_L g4722 ( 
.A(n_4332),
.B(n_13),
.Y(n_4722)
);

AND2x6_ASAP7_75t_L g4723 ( 
.A(n_4441),
.B(n_4133),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4430),
.Y(n_4724)
);

NOR2xp33_ASAP7_75t_R g4725 ( 
.A(n_4302),
.B(n_4157),
.Y(n_4725)
);

NAND2x1p5_ASAP7_75t_L g4726 ( 
.A(n_4510),
.B(n_4133),
.Y(n_4726)
);

INVx1_ASAP7_75t_SL g4727 ( 
.A(n_4375),
.Y(n_4727)
);

AOI22xp33_ASAP7_75t_L g4728 ( 
.A1(n_4396),
.A2(n_4051),
.B1(n_3937),
.B2(n_3962),
.Y(n_4728)
);

BUFx6f_ASAP7_75t_L g4729 ( 
.A(n_4476),
.Y(n_4729)
);

INVx1_ASAP7_75t_L g4730 ( 
.A(n_4431),
.Y(n_4730)
);

NOR2xp33_ASAP7_75t_L g4731 ( 
.A(n_4543),
.B(n_15),
.Y(n_4731)
);

NOR2xp33_ASAP7_75t_L g4732 ( 
.A(n_4366),
.B(n_15),
.Y(n_4732)
);

AOI21xp5_ASAP7_75t_L g4733 ( 
.A1(n_4536),
.A2(n_4198),
.B(n_4169),
.Y(n_4733)
);

O2A1O1Ixp33_ASAP7_75t_L g4734 ( 
.A1(n_4490),
.A2(n_2202),
.B(n_2206),
.C(n_2198),
.Y(n_4734)
);

OAI21xp33_ASAP7_75t_L g4735 ( 
.A1(n_4357),
.A2(n_4358),
.B(n_4413),
.Y(n_4735)
);

AND2x4_ASAP7_75t_L g4736 ( 
.A(n_4471),
.B(n_4133),
.Y(n_4736)
);

NOR2xp33_ASAP7_75t_L g4737 ( 
.A(n_4291),
.B(n_16),
.Y(n_4737)
);

INVx1_ASAP7_75t_L g4738 ( 
.A(n_4436),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4593),
.Y(n_4739)
);

O2A1O1Ixp33_ASAP7_75t_L g4740 ( 
.A1(n_4499),
.A2(n_2206),
.B(n_2214),
.C(n_2202),
.Y(n_4740)
);

A2O1A1Ixp33_ASAP7_75t_L g4741 ( 
.A1(n_4450),
.A2(n_4259),
.B(n_4167),
.C(n_4191),
.Y(n_4741)
);

OAI22xp33_ASAP7_75t_L g4742 ( 
.A1(n_4453),
.A2(n_4238),
.B1(n_4220),
.B2(n_3996),
.Y(n_4742)
);

AOI222xp33_ASAP7_75t_L g4743 ( 
.A1(n_4530),
.A2(n_2155),
.B1(n_2151),
.B2(n_2152),
.C1(n_2149),
.C2(n_871),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_4318),
.B(n_4143),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4279),
.B(n_4145),
.Y(n_4745)
);

NOR2xp33_ASAP7_75t_L g4746 ( 
.A(n_4303),
.B(n_17),
.Y(n_4746)
);

A2O1A1Ixp33_ASAP7_75t_L g4747 ( 
.A1(n_4454),
.A2(n_4183),
.B(n_4149),
.C(n_4156),
.Y(n_4747)
);

A2O1A1Ixp33_ASAP7_75t_L g4748 ( 
.A1(n_4477),
.A2(n_4158),
.B(n_4161),
.C(n_4147),
.Y(n_4748)
);

OAI22xp5_ASAP7_75t_L g4749 ( 
.A1(n_4535),
.A2(n_4016),
.B1(n_3998),
.B2(n_4168),
.Y(n_4749)
);

NOR2xp33_ASAP7_75t_L g4750 ( 
.A(n_4377),
.B(n_18),
.Y(n_4750)
);

NOR2xp33_ASAP7_75t_L g4751 ( 
.A(n_4407),
.B(n_4411),
.Y(n_4751)
);

AOI21xp5_ASAP7_75t_L g4752 ( 
.A1(n_4582),
.A2(n_4198),
.B(n_4084),
.Y(n_4752)
);

AOI21xp5_ASAP7_75t_L g4753 ( 
.A1(n_4282),
.A2(n_4262),
.B(n_4261),
.Y(n_4753)
);

NOR2xp33_ASAP7_75t_L g4754 ( 
.A(n_4398),
.B(n_20),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4281),
.B(n_4174),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_SL g4756 ( 
.A(n_4517),
.B(n_3996),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_SL g4757 ( 
.A(n_4517),
.B(n_3996),
.Y(n_4757)
);

OAI22xp5_ASAP7_75t_L g4758 ( 
.A1(n_4596),
.A2(n_4238),
.B1(n_4220),
.B2(n_4008),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4548),
.B(n_4192),
.Y(n_4759)
);

INVx2_ASAP7_75t_SL g4760 ( 
.A(n_4517),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4531),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4564),
.B(n_4192),
.Y(n_4762)
);

BUFx4f_ASAP7_75t_SL g4763 ( 
.A(n_4529),
.Y(n_4763)
);

OAI22xp5_ASAP7_75t_L g4764 ( 
.A1(n_4469),
.A2(n_4238),
.B1(n_4220),
.B2(n_4008),
.Y(n_4764)
);

AOI21xp5_ASAP7_75t_L g4765 ( 
.A1(n_4360),
.A2(n_4211),
.B(n_4210),
.Y(n_4765)
);

AOI22xp5_ASAP7_75t_L g4766 ( 
.A1(n_4549),
.A2(n_4008),
.B1(n_2151),
.B2(n_2152),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_SL g4767 ( 
.A(n_4587),
.B(n_4473),
.Y(n_4767)
);

INVx1_ASAP7_75t_L g4768 ( 
.A(n_4572),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4474),
.Y(n_4769)
);

HB1xp67_ASAP7_75t_L g4770 ( 
.A(n_4565),
.Y(n_4770)
);

INVx2_ASAP7_75t_L g4771 ( 
.A(n_4480),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4482),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4492),
.Y(n_4773)
);

INVx2_ASAP7_75t_SL g4774 ( 
.A(n_4587),
.Y(n_4774)
);

AOI21xp5_ASAP7_75t_L g4775 ( 
.A1(n_4295),
.A2(n_4211),
.B(n_4210),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4503),
.Y(n_4776)
);

BUFx6f_ASAP7_75t_L g4777 ( 
.A(n_4302),
.Y(n_4777)
);

NOR2xp33_ASAP7_75t_L g4778 ( 
.A(n_4403),
.B(n_20),
.Y(n_4778)
);

NAND2xp5_ASAP7_75t_SL g4779 ( 
.A(n_4443),
.B(n_4123),
.Y(n_4779)
);

BUFx6f_ASAP7_75t_L g4780 ( 
.A(n_4506),
.Y(n_4780)
);

AOI21xp5_ASAP7_75t_L g4781 ( 
.A1(n_4308),
.A2(n_4237),
.B(n_4226),
.Y(n_4781)
);

OAI22xp5_ASAP7_75t_L g4782 ( 
.A1(n_4414),
.A2(n_2965),
.B1(n_2975),
.B2(n_2914),
.Y(n_4782)
);

NAND2xp5_ASAP7_75t_SL g4783 ( 
.A(n_4401),
.B(n_4406),
.Y(n_4783)
);

AOI21xp5_ASAP7_75t_L g4784 ( 
.A1(n_4558),
.A2(n_4237),
.B(n_4226),
.Y(n_4784)
);

A2O1A1Ixp33_ASAP7_75t_L g4785 ( 
.A1(n_4526),
.A2(n_2151),
.B(n_2152),
.C(n_2149),
.Y(n_4785)
);

OAI22x1_ASAP7_75t_L g4786 ( 
.A1(n_4301),
.A2(n_4196),
.B1(n_4242),
.B2(n_4150),
.Y(n_4786)
);

NOR2xp33_ASAP7_75t_L g4787 ( 
.A(n_4420),
.B(n_21),
.Y(n_4787)
);

OAI22xp5_ASAP7_75t_L g4788 ( 
.A1(n_4286),
.A2(n_2965),
.B1(n_2975),
.B2(n_2914),
.Y(n_4788)
);

A2O1A1Ixp33_ASAP7_75t_L g4789 ( 
.A1(n_4532),
.A2(n_2155),
.B(n_2152),
.C(n_863),
.Y(n_4789)
);

NOR2xp33_ASAP7_75t_L g4790 ( 
.A(n_4422),
.B(n_22),
.Y(n_4790)
);

OAI21x1_ASAP7_75t_L g4791 ( 
.A1(n_4524),
.A2(n_4383),
.B(n_4424),
.Y(n_4791)
);

O2A1O1Ixp33_ASAP7_75t_L g4792 ( 
.A1(n_4518),
.A2(n_2233),
.B(n_2065),
.C(n_2068),
.Y(n_4792)
);

BUFx2_ASAP7_75t_L g4793 ( 
.A(n_4559),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_SL g4794 ( 
.A(n_4401),
.B(n_4150),
.Y(n_4794)
);

AOI21xp5_ASAP7_75t_L g4795 ( 
.A1(n_4317),
.A2(n_4179),
.B(n_4172),
.Y(n_4795)
);

AOI21xp5_ASAP7_75t_L g4796 ( 
.A1(n_4550),
.A2(n_4179),
.B(n_4172),
.Y(n_4796)
);

NOR2xp33_ASAP7_75t_L g4797 ( 
.A(n_4432),
.B(n_22),
.Y(n_4797)
);

NOR2xp33_ASAP7_75t_L g4798 ( 
.A(n_4433),
.B(n_24),
.Y(n_4798)
);

AOI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4321),
.A2(n_4188),
.B(n_4185),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_SL g4800 ( 
.A(n_4406),
.B(n_4185),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_SL g4801 ( 
.A(n_4425),
.B(n_4083),
.Y(n_4801)
);

BUFx12f_ASAP7_75t_L g4802 ( 
.A(n_4539),
.Y(n_4802)
);

CKINVDCx5p33_ASAP7_75t_R g4803 ( 
.A(n_4292),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4566),
.Y(n_4804)
);

A2O1A1Ixp33_ASAP7_75t_L g4805 ( 
.A1(n_4523),
.A2(n_2155),
.B(n_864),
.C(n_872),
.Y(n_4805)
);

INVx2_ASAP7_75t_L g4806 ( 
.A(n_4577),
.Y(n_4806)
);

NAND2xp5_ASAP7_75t_SL g4807 ( 
.A(n_4425),
.B(n_4083),
.Y(n_4807)
);

CKINVDCx5p33_ASAP7_75t_R g4808 ( 
.A(n_4299),
.Y(n_4808)
);

BUFx6f_ASAP7_75t_L g4809 ( 
.A(n_4506),
.Y(n_4809)
);

CKINVDCx16_ASAP7_75t_R g4810 ( 
.A(n_4438),
.Y(n_4810)
);

OAI21xp5_ASAP7_75t_L g4811 ( 
.A1(n_4469),
.A2(n_4103),
.B(n_4094),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4573),
.B(n_4094),
.Y(n_4812)
);

INVx2_ASAP7_75t_SL g4813 ( 
.A(n_4534),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_SL g4814 ( 
.A(n_4307),
.B(n_4103),
.Y(n_4814)
);

A2O1A1Ixp33_ASAP7_75t_L g4815 ( 
.A1(n_4484),
.A2(n_2155),
.B(n_873),
.C(n_876),
.Y(n_4815)
);

BUFx2_ASAP7_75t_L g4816 ( 
.A(n_4559),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4381),
.B(n_3929),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4573),
.B(n_3989),
.Y(n_4818)
);

BUFx4f_ASAP7_75t_L g4819 ( 
.A(n_4367),
.Y(n_4819)
);

O2A1O1Ixp33_ASAP7_75t_L g4820 ( 
.A1(n_4541),
.A2(n_2077),
.B(n_2078),
.C(n_2064),
.Y(n_4820)
);

BUFx2_ASAP7_75t_L g4821 ( 
.A(n_4439),
.Y(n_4821)
);

OAI21xp33_ASAP7_75t_SL g4822 ( 
.A1(n_4434),
.A2(n_3410),
.B(n_3388),
.Y(n_4822)
);

OAI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_4491),
.A2(n_952),
.B1(n_833),
.B2(n_693),
.Y(n_4823)
);

AOI22xp33_ASAP7_75t_L g4824 ( 
.A1(n_4547),
.A2(n_3992),
.B1(n_4006),
.B2(n_3989),
.Y(n_4824)
);

CKINVDCx16_ASAP7_75t_R g4825 ( 
.A(n_4439),
.Y(n_4825)
);

AND2x2_ASAP7_75t_L g4826 ( 
.A(n_4381),
.B(n_4389),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4585),
.Y(n_4827)
);

NAND3xp33_ASAP7_75t_SL g4828 ( 
.A(n_4478),
.B(n_878),
.C(n_862),
.Y(n_4828)
);

NAND2xp5_ASAP7_75t_L g4829 ( 
.A(n_4278),
.B(n_3992),
.Y(n_4829)
);

CKINVDCx5p33_ASAP7_75t_R g4830 ( 
.A(n_4437),
.Y(n_4830)
);

BUFx6f_ASAP7_75t_L g4831 ( 
.A(n_4534),
.Y(n_4831)
);

AOI22xp33_ASAP7_75t_L g4832 ( 
.A1(n_4327),
.A2(n_4013),
.B1(n_4019),
.B2(n_4006),
.Y(n_4832)
);

INVx3_ASAP7_75t_SL g4833 ( 
.A(n_4367),
.Y(n_4833)
);

AOI22xp5_ASAP7_75t_L g4834 ( 
.A1(n_4288),
.A2(n_2073),
.B1(n_2123),
.B2(n_2054),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4594),
.Y(n_4835)
);

BUFx6f_ASAP7_75t_L g4836 ( 
.A(n_4563),
.Y(n_4836)
);

OR2x2_ASAP7_75t_L g4837 ( 
.A(n_4309),
.B(n_4013),
.Y(n_4837)
);

AOI221xp5_ASAP7_75t_SL g4838 ( 
.A1(n_4483),
.A2(n_742),
.B1(n_815),
.B2(n_693),
.C(n_676),
.Y(n_4838)
);

NOR2xp33_ASAP7_75t_SL g4839 ( 
.A(n_4382),
.B(n_3468),
.Y(n_4839)
);

A2O1A1Ixp33_ASAP7_75t_L g4840 ( 
.A1(n_4530),
.A2(n_882),
.B(n_883),
.C(n_881),
.Y(n_4840)
);

NOR2xp33_ASAP7_75t_L g4841 ( 
.A(n_4440),
.B(n_24),
.Y(n_4841)
);

A2O1A1Ixp33_ASAP7_75t_L g4842 ( 
.A1(n_4368),
.A2(n_885),
.B(n_887),
.C(n_884),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4274),
.B(n_4021),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_R g4844 ( 
.A(n_4563),
.B(n_26),
.Y(n_4844)
);

AOI21xp5_ASAP7_75t_L g4845 ( 
.A1(n_4272),
.A2(n_3497),
.B(n_3472),
.Y(n_4845)
);

NAND2xp5_ASAP7_75t_L g4846 ( 
.A(n_4376),
.B(n_4021),
.Y(n_4846)
);

NOR2xp33_ASAP7_75t_L g4847 ( 
.A(n_4445),
.B(n_4446),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_SL g4848 ( 
.A(n_4400),
.B(n_4023),
.Y(n_4848)
);

OAI21xp33_ASAP7_75t_L g4849 ( 
.A1(n_4528),
.A2(n_693),
.B(n_676),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4455),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4455),
.Y(n_4851)
);

CKINVDCx14_ASAP7_75t_R g4852 ( 
.A(n_4460),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_SL g4853 ( 
.A(n_4400),
.B(n_4023),
.Y(n_4853)
);

NOR2xp33_ASAP7_75t_L g4854 ( 
.A(n_4447),
.B(n_27),
.Y(n_4854)
);

BUFx2_ASAP7_75t_L g4855 ( 
.A(n_4439),
.Y(n_4855)
);

A2O1A1Ixp33_ASAP7_75t_L g4856 ( 
.A1(n_4567),
.A2(n_891),
.B(n_892),
.C(n_888),
.Y(n_4856)
);

OAI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4451),
.A2(n_2965),
.B1(n_2975),
.B2(n_2914),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4452),
.B(n_4048),
.Y(n_4858)
);

BUFx6f_ASAP7_75t_L g4859 ( 
.A(n_4348),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_SL g4860 ( 
.A(n_4556),
.B(n_4035),
.Y(n_4860)
);

A2O1A1Ixp33_ASAP7_75t_L g4861 ( 
.A1(n_4574),
.A2(n_894),
.B(n_895),
.C(n_890),
.Y(n_4861)
);

BUFx6f_ASAP7_75t_L g4862 ( 
.A(n_4348),
.Y(n_4862)
);

INVx3_ASAP7_75t_SL g4863 ( 
.A(n_4556),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4455),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4457),
.B(n_4458),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4561),
.Y(n_4866)
);

AO32x2_ASAP7_75t_L g4867 ( 
.A1(n_4540),
.A2(n_4589),
.A3(n_4298),
.B1(n_4306),
.B2(n_4557),
.Y(n_4867)
);

NOR2xp33_ASAP7_75t_L g4868 ( 
.A(n_4461),
.B(n_29),
.Y(n_4868)
);

O2A1O1Ixp5_ASAP7_75t_L g4869 ( 
.A1(n_4583),
.A2(n_2078),
.B(n_2084),
.C(n_2081),
.Y(n_4869)
);

OAI22xp5_ASAP7_75t_L g4870 ( 
.A1(n_4545),
.A2(n_1016),
.B1(n_742),
.B2(n_815),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4465),
.B(n_4035),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4468),
.B(n_4036),
.Y(n_4872)
);

AO31x2_ASAP7_75t_L g4873 ( 
.A1(n_4359),
.A2(n_4038),
.A3(n_4040),
.B(n_4036),
.Y(n_4873)
);

AOI21xp5_ASAP7_75t_L g4874 ( 
.A1(n_4568),
.A2(n_3507),
.B(n_3499),
.Y(n_4874)
);

BUFx2_ASAP7_75t_L g4875 ( 
.A(n_4551),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4389),
.B(n_4038),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4561),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_SL g4878 ( 
.A(n_4498),
.B(n_4040),
.Y(n_4878)
);

AO21x1_ASAP7_75t_L g4879 ( 
.A1(n_4486),
.A2(n_2043),
.B(n_2093),
.Y(n_4879)
);

A2O1A1Ixp33_ASAP7_75t_L g4880 ( 
.A1(n_4382),
.A2(n_896),
.B(n_899),
.C(n_893),
.Y(n_4880)
);

OA21x2_ASAP7_75t_L g4881 ( 
.A1(n_4331),
.A2(n_4055),
.B(n_4048),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_SL g4882 ( 
.A(n_4378),
.B(n_4055),
.Y(n_4882)
);

AOI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_4581),
.A2(n_3507),
.B(n_3499),
.Y(n_4883)
);

OAI22xp5_ASAP7_75t_L g4884 ( 
.A1(n_4487),
.A2(n_4502),
.B1(n_4511),
.B2(n_4494),
.Y(n_4884)
);

OAI22xp5_ASAP7_75t_SL g4885 ( 
.A1(n_4512),
.A2(n_901),
.B1(n_902),
.B2(n_897),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4514),
.B(n_4063),
.Y(n_4886)
);

OAI21xp5_ASAP7_75t_L g4887 ( 
.A1(n_4579),
.A2(n_2073),
.B(n_2054),
.Y(n_4887)
);

OAI22xp5_ASAP7_75t_L g4888 ( 
.A1(n_4516),
.A2(n_940),
.B1(n_742),
.B2(n_815),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_SL g4889 ( 
.A(n_4378),
.B(n_4533),
.Y(n_4889)
);

INVx3_ASAP7_75t_L g4890 ( 
.A(n_4580),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_SL g4891 ( 
.A(n_4542),
.B(n_4062),
.Y(n_4891)
);

AOI22xp33_ASAP7_75t_L g4892 ( 
.A1(n_4555),
.A2(n_4092),
.B1(n_4093),
.B2(n_4062),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_SL g4893 ( 
.A(n_4495),
.B(n_4092),
.Y(n_4893)
);

NOR2xp33_ASAP7_75t_L g4894 ( 
.A(n_4449),
.B(n_30),
.Y(n_4894)
);

INVx2_ASAP7_75t_L g4895 ( 
.A(n_4561),
.Y(n_4895)
);

AOI21xp5_ASAP7_75t_L g4896 ( 
.A1(n_4515),
.A2(n_2980),
.B(n_2976),
.Y(n_4896)
);

A2O1A1Ixp33_ASAP7_75t_L g4897 ( 
.A1(n_4575),
.A2(n_908),
.B(n_911),
.C(n_909),
.Y(n_4897)
);

INVx2_ASAP7_75t_L g4898 ( 
.A(n_4326),
.Y(n_4898)
);

AOI21xp5_ASAP7_75t_L g4899 ( 
.A1(n_4334),
.A2(n_2988),
.B(n_2982),
.Y(n_4899)
);

A2O1A1Ixp33_ASAP7_75t_L g4900 ( 
.A1(n_4576),
.A2(n_914),
.B(n_917),
.C(n_916),
.Y(n_4900)
);

AOI21xp5_ASAP7_75t_L g4901 ( 
.A1(n_4560),
.A2(n_2988),
.B(n_2982),
.Y(n_4901)
);

HB1xp67_ASAP7_75t_L g4902 ( 
.A(n_4495),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4562),
.A2(n_2994),
.B(n_2990),
.Y(n_4903)
);

BUFx3_ASAP7_75t_L g4904 ( 
.A(n_4580),
.Y(n_4904)
);

BUFx2_ASAP7_75t_L g4905 ( 
.A(n_4365),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4588),
.B(n_4093),
.Y(n_4906)
);

INVx2_ASAP7_75t_L g4907 ( 
.A(n_4391),
.Y(n_4907)
);

NOR2xp33_ASAP7_75t_L g4908 ( 
.A(n_4525),
.B(n_30),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4412),
.Y(n_4909)
);

NOR3xp33_ASAP7_75t_SL g4910 ( 
.A(n_4472),
.B(n_920),
.C(n_906),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_SL g4911 ( 
.A(n_4521),
.B(n_3137),
.Y(n_4911)
);

INVx3_ASAP7_75t_L g4912 ( 
.A(n_4365),
.Y(n_4912)
);

AOI22xp5_ASAP7_75t_L g4913 ( 
.A1(n_4312),
.A2(n_2073),
.B1(n_2123),
.B2(n_2054),
.Y(n_4913)
);

NOR2xp33_ASAP7_75t_L g4914 ( 
.A(n_4475),
.B(n_31),
.Y(n_4914)
);

A2O1A1Ixp33_ASAP7_75t_L g4915 ( 
.A1(n_4481),
.A2(n_929),
.B(n_931),
.C(n_926),
.Y(n_4915)
);

AOI21xp5_ASAP7_75t_L g4916 ( 
.A1(n_4341),
.A2(n_3002),
.B(n_2889),
.Y(n_4916)
);

BUFx6f_ASAP7_75t_L g4917 ( 
.A(n_4365),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4520),
.Y(n_4918)
);

AND2x4_ASAP7_75t_L g4919 ( 
.A(n_4276),
.B(n_3459),
.Y(n_4919)
);

BUFx6f_ASAP7_75t_L g4920 ( 
.A(n_4626),
.Y(n_4920)
);

AOI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4633),
.A2(n_4405),
.B(n_4489),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_4709),
.B(n_4595),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_SL g4923 ( 
.A(n_4658),
.B(n_4546),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4609),
.B(n_4544),
.Y(n_4924)
);

AOI21x1_ASAP7_75t_L g4925 ( 
.A1(n_4663),
.A2(n_4527),
.B(n_4522),
.Y(n_4925)
);

OAI21xp5_ASAP7_75t_L g4926 ( 
.A1(n_4629),
.A2(n_4570),
.B(n_4335),
.Y(n_4926)
);

NAND3x1_ASAP7_75t_L g4927 ( 
.A(n_4649),
.B(n_4361),
.C(n_4552),
.Y(n_4927)
);

AND3x1_ASAP7_75t_SL g4928 ( 
.A(n_4852),
.B(n_32),
.C(n_33),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4609),
.B(n_4352),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4612),
.B(n_4355),
.Y(n_4930)
);

AOI21xp5_ASAP7_75t_L g4931 ( 
.A1(n_4603),
.A2(n_4405),
.B(n_4497),
.Y(n_4931)
);

AO31x2_ASAP7_75t_L g4932 ( 
.A1(n_4786),
.A2(n_4399),
.A3(n_4402),
.B(n_4371),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4612),
.B(n_4618),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4615),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_SL g4935 ( 
.A(n_4825),
.B(n_4519),
.Y(n_4935)
);

INVx5_ASAP7_75t_L g4936 ( 
.A(n_4723),
.Y(n_4936)
);

OAI21x1_ASAP7_75t_L g4937 ( 
.A1(n_4791),
.A2(n_4538),
.B(n_4384),
.Y(n_4937)
);

O2A1O1Ixp5_ASAP7_75t_L g4938 ( 
.A1(n_4889),
.A2(n_4315),
.B(n_4354),
.C(n_4305),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4613),
.B(n_4578),
.Y(n_4939)
);

OAI21xp5_ASAP7_75t_L g4940 ( 
.A1(n_4675),
.A2(n_4463),
.B(n_4462),
.Y(n_4940)
);

INVx1_ASAP7_75t_SL g4941 ( 
.A(n_4688),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4640),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4628),
.Y(n_4943)
);

INVx5_ASAP7_75t_L g4944 ( 
.A(n_4723),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4739),
.B(n_4467),
.Y(n_4945)
);

OAI21x1_ASAP7_75t_L g4946 ( 
.A1(n_4697),
.A2(n_4390),
.B(n_4373),
.Y(n_4946)
);

BUFx4f_ASAP7_75t_SL g4947 ( 
.A(n_4597),
.Y(n_4947)
);

OAI21xp5_ASAP7_75t_L g4948 ( 
.A1(n_4679),
.A2(n_4508),
.B(n_4507),
.Y(n_4948)
);

AO21x2_ASAP7_75t_L g4949 ( 
.A1(n_4866),
.A2(n_4393),
.B(n_4392),
.Y(n_4949)
);

AOI21x1_ASAP7_75t_SL g4950 ( 
.A1(n_4865),
.A2(n_2043),
.B(n_2093),
.Y(n_4950)
);

AOI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4718),
.A2(n_4444),
.B(n_4504),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4677),
.B(n_4584),
.Y(n_4952)
);

OAI21x1_ASAP7_75t_SL g4953 ( 
.A1(n_4669),
.A2(n_4604),
.B(n_4602),
.Y(n_4953)
);

AO31x2_ASAP7_75t_L g4954 ( 
.A1(n_4898),
.A2(n_3181),
.A3(n_3179),
.B(n_2769),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4621),
.B(n_693),
.Y(n_4955)
);

INVx4_ASAP7_75t_L g4956 ( 
.A(n_4763),
.Y(n_4956)
);

INVx2_ASAP7_75t_L g4957 ( 
.A(n_4634),
.Y(n_4957)
);

OA22x2_ASAP7_75t_L g4958 ( 
.A1(n_4598),
.A2(n_933),
.B1(n_935),
.B2(n_930),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4599),
.B(n_742),
.Y(n_4959)
);

OAI21xp5_ASAP7_75t_L g4960 ( 
.A1(n_4680),
.A2(n_937),
.B(n_936),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4770),
.B(n_815),
.Y(n_4961)
);

CKINVDCx5p33_ASAP7_75t_R g4962 ( 
.A(n_4655),
.Y(n_4962)
);

OAI21x1_ASAP7_75t_L g4963 ( 
.A1(n_4707),
.A2(n_2769),
.B(n_2765),
.Y(n_4963)
);

NAND3xp33_ASAP7_75t_SL g4964 ( 
.A(n_4844),
.B(n_943),
.C(n_941),
.Y(n_4964)
);

AOI21xp5_ASAP7_75t_L g4965 ( 
.A1(n_4606),
.A2(n_3002),
.B(n_3026),
.Y(n_4965)
);

OAI21xp33_ASAP7_75t_SL g4966 ( 
.A1(n_4617),
.A2(n_3189),
.B(n_3187),
.Y(n_4966)
);

AOI21xp5_ASAP7_75t_L g4967 ( 
.A1(n_4625),
.A2(n_3029),
.B(n_3026),
.Y(n_4967)
);

BUFx12f_ASAP7_75t_L g4968 ( 
.A(n_4659),
.Y(n_4968)
);

OAI21x1_ASAP7_75t_L g4969 ( 
.A1(n_4692),
.A2(n_2769),
.B(n_2765),
.Y(n_4969)
);

AOI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4653),
.A2(n_4624),
.B(n_4614),
.Y(n_4970)
);

O2A1O1Ixp33_ASAP7_75t_L g4971 ( 
.A1(n_4667),
.A2(n_2103),
.B(n_2114),
.C(n_2090),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_L g4972 ( 
.A(n_4654),
.B(n_833),
.Y(n_4972)
);

NOR2xp67_ASAP7_75t_L g4973 ( 
.A(n_4648),
.B(n_32),
.Y(n_4973)
);

OAI22xp5_ASAP7_75t_L g4974 ( 
.A1(n_4704),
.A2(n_4746),
.B1(n_4737),
.B2(n_4880),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4638),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4701),
.B(n_833),
.Y(n_4976)
);

NAND2xp33_ASAP7_75t_L g4977 ( 
.A(n_4611),
.B(n_4777),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4641),
.Y(n_4978)
);

OAI21xp5_ASAP7_75t_L g4979 ( 
.A1(n_4908),
.A2(n_4894),
.B(n_4731),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4605),
.A2(n_3052),
.B(n_3029),
.Y(n_4980)
);

INVx2_ASAP7_75t_L g4981 ( 
.A(n_4642),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4601),
.B(n_833),
.Y(n_4982)
);

BUFx12f_ASAP7_75t_L g4983 ( 
.A(n_4803),
.Y(n_4983)
);

NOR2xp67_ASAP7_75t_SL g4984 ( 
.A(n_4802),
.B(n_940),
.Y(n_4984)
);

AO31x2_ASAP7_75t_L g4985 ( 
.A1(n_4850),
.A2(n_2919),
.A3(n_2922),
.B(n_2781),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_SL g4986 ( 
.A(n_4600),
.B(n_940),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4639),
.B(n_940),
.Y(n_4987)
);

NAND2x1p5_ASAP7_75t_L g4988 ( 
.A(n_4608),
.B(n_3052),
.Y(n_4988)
);

O2A1O1Ixp5_ASAP7_75t_L g4989 ( 
.A1(n_4767),
.A2(n_4702),
.B(n_4703),
.C(n_4691),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4674),
.B(n_940),
.Y(n_4990)
);

NOR2x1_ASAP7_75t_SL g4991 ( 
.A(n_4608),
.B(n_3459),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4664),
.B(n_952),
.Y(n_4992)
);

NAND2xp5_ASAP7_75t_L g4993 ( 
.A(n_4745),
.B(n_952),
.Y(n_4993)
);

A2O1A1Ixp33_ASAP7_75t_L g4994 ( 
.A1(n_4720),
.A2(n_964),
.B(n_986),
.C(n_958),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_SL g4995 ( 
.A(n_4810),
.B(n_952),
.Y(n_4995)
);

AOI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4845),
.A2(n_3062),
.B(n_3054),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4755),
.B(n_952),
.Y(n_4997)
);

OAI21xp5_ASAP7_75t_L g4998 ( 
.A1(n_4632),
.A2(n_949),
.B(n_947),
.Y(n_4998)
);

AOI31xp67_ASAP7_75t_L g4999 ( 
.A1(n_4895),
.A2(n_2125),
.A3(n_2126),
.B(n_2119),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4616),
.B(n_1016),
.Y(n_5000)
);

NOR2x1_ASAP7_75t_L g5001 ( 
.A(n_4623),
.B(n_3054),
.Y(n_5001)
);

OAI21x1_ASAP7_75t_L g5002 ( 
.A1(n_4753),
.A2(n_2919),
.B(n_2781),
.Y(n_5002)
);

AOI22xp33_ASAP7_75t_L g5003 ( 
.A1(n_4696),
.A2(n_2838),
.B1(n_2841),
.B2(n_2837),
.Y(n_5003)
);

AND2x2_ASAP7_75t_L g5004 ( 
.A(n_4708),
.B(n_1016),
.Y(n_5004)
);

OAI21x1_ASAP7_75t_L g5005 ( 
.A1(n_4662),
.A2(n_2924),
.B(n_2922),
.Y(n_5005)
);

AOI21x1_ASAP7_75t_L g5006 ( 
.A1(n_4891),
.A2(n_2125),
.B(n_2119),
.Y(n_5006)
);

NOR2xp67_ASAP7_75t_SL g5007 ( 
.A(n_4608),
.B(n_1047),
.Y(n_5007)
);

AOI21x1_ASAP7_75t_L g5008 ( 
.A1(n_4877),
.A2(n_2130),
.B(n_2126),
.Y(n_5008)
);

A2O1A1Ixp33_ASAP7_75t_L g5009 ( 
.A1(n_4754),
.A2(n_984),
.B(n_996),
.C(n_960),
.Y(n_5009)
);

INVx2_ASAP7_75t_L g5010 ( 
.A(n_4643),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4672),
.Y(n_5011)
);

INVx3_ASAP7_75t_L g5012 ( 
.A(n_4626),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_SL g5013 ( 
.A(n_4626),
.B(n_1047),
.Y(n_5013)
);

AO31x2_ASAP7_75t_L g5014 ( 
.A1(n_4851),
.A2(n_2922),
.A3(n_2926),
.B(n_2924),
.Y(n_5014)
);

AOI21xp5_ASAP7_75t_L g5015 ( 
.A1(n_4644),
.A2(n_3062),
.B(n_3054),
.Y(n_5015)
);

AOI21xp5_ASAP7_75t_L g5016 ( 
.A1(n_4630),
.A2(n_3062),
.B(n_3054),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_SL g5017 ( 
.A(n_4665),
.B(n_1047),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_L g5018 ( 
.A(n_4666),
.B(n_1047),
.Y(n_5018)
);

AO31x2_ASAP7_75t_L g5019 ( 
.A1(n_4864),
.A2(n_2924),
.A3(n_2930),
.B(n_2926),
.Y(n_5019)
);

A2O1A1Ixp33_ASAP7_75t_L g5020 ( 
.A1(n_4778),
.A2(n_4750),
.B(n_4732),
.C(n_4787),
.Y(n_5020)
);

AO31x2_ASAP7_75t_L g5021 ( 
.A1(n_4796),
.A2(n_2926),
.A3(n_2935),
.B(n_2930),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4711),
.Y(n_5022)
);

NOR2xp33_ASAP7_75t_L g5023 ( 
.A(n_4735),
.B(n_33),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4636),
.B(n_1047),
.Y(n_5024)
);

NOR2xp33_ASAP7_75t_SL g5025 ( 
.A(n_4808),
.B(n_3062),
.Y(n_5025)
);

AOI21xp5_ASAP7_75t_L g5026 ( 
.A1(n_4874),
.A2(n_3119),
.B(n_3075),
.Y(n_5026)
);

O2A1O1Ixp5_ASAP7_75t_L g5027 ( 
.A1(n_4794),
.A2(n_3119),
.B(n_3156),
.C(n_3075),
.Y(n_5027)
);

AOI22x1_ASAP7_75t_L g5028 ( 
.A1(n_4863),
.A2(n_4830),
.B1(n_4813),
.B2(n_4816),
.Y(n_5028)
);

CKINVDCx8_ASAP7_75t_R g5029 ( 
.A(n_4721),
.Y(n_5029)
);

A2O1A1Ixp33_ASAP7_75t_L g5030 ( 
.A1(n_4700),
.A2(n_972),
.B(n_989),
.C(n_957),
.Y(n_5030)
);

NAND2xp5_ASAP7_75t_SL g5031 ( 
.A(n_4665),
.B(n_3075),
.Y(n_5031)
);

AOI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_4883),
.A2(n_3119),
.B(n_3075),
.Y(n_5032)
);

OAI21x1_ASAP7_75t_SL g5033 ( 
.A1(n_4716),
.A2(n_2136),
.B(n_2130),
.Y(n_5033)
);

BUFx2_ASAP7_75t_L g5034 ( 
.A(n_4646),
.Y(n_5034)
);

AOI21xp5_ASAP7_75t_L g5035 ( 
.A1(n_4714),
.A2(n_3156),
.B(n_3119),
.Y(n_5035)
);

AOI21xp5_ASAP7_75t_L g5036 ( 
.A1(n_4749),
.A2(n_3156),
.B(n_2861),
.Y(n_5036)
);

AO31x2_ASAP7_75t_L g5037 ( 
.A1(n_4906),
.A2(n_4781),
.A3(n_4775),
.B(n_4799),
.Y(n_5037)
);

OAI21x1_ASAP7_75t_L g5038 ( 
.A1(n_4752),
.A2(n_2939),
.B(n_3156),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_4858),
.B(n_832),
.Y(n_5039)
);

AOI221x1_ASAP7_75t_L g5040 ( 
.A1(n_4884),
.A2(n_1510),
.B1(n_1512),
.B2(n_1365),
.C(n_1350),
.Y(n_5040)
);

CKINVDCx5p33_ASAP7_75t_R g5041 ( 
.A(n_4657),
.Y(n_5041)
);

AOI22xp33_ASAP7_75t_L g5042 ( 
.A1(n_4743),
.A2(n_2838),
.B1(n_2856),
.B2(n_2841),
.Y(n_5042)
);

AOI22xp5_ASAP7_75t_L g5043 ( 
.A1(n_4849),
.A2(n_2123),
.B1(n_2138),
.B2(n_2054),
.Y(n_5043)
);

INVx3_ASAP7_75t_L g5044 ( 
.A(n_4665),
.Y(n_5044)
);

INVx2_ASAP7_75t_L g5045 ( 
.A(n_4684),
.Y(n_5045)
);

OAI21x1_ASAP7_75t_L g5046 ( 
.A1(n_4765),
.A2(n_2431),
.B(n_2136),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4871),
.B(n_875),
.Y(n_5047)
);

AND2x4_ASAP7_75t_L g5048 ( 
.A(n_4890),
.B(n_1350),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_L g5049 ( 
.A(n_4872),
.B(n_875),
.Y(n_5049)
);

INVx2_ASAP7_75t_L g5050 ( 
.A(n_4685),
.Y(n_5050)
);

INVxp67_ASAP7_75t_L g5051 ( 
.A(n_4875),
.Y(n_5051)
);

AND2x4_ASAP7_75t_L g5052 ( 
.A(n_4890),
.B(n_1350),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4886),
.B(n_875),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_L g5054 ( 
.A1(n_4764),
.A2(n_3193),
.B(n_3188),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4761),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4727),
.B(n_875),
.Y(n_5056)
);

OAI22xp33_ASAP7_75t_L g5057 ( 
.A1(n_4839),
.A2(n_3189),
.B1(n_3190),
.B2(n_3187),
.Y(n_5057)
);

INVx2_ASAP7_75t_L g5058 ( 
.A(n_4686),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_4768),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_4744),
.B(n_875),
.Y(n_5060)
);

NOR2xp33_ASAP7_75t_L g5061 ( 
.A(n_4884),
.B(n_34),
.Y(n_5061)
);

OAI21x1_ASAP7_75t_SL g5062 ( 
.A1(n_4733),
.A2(n_3188),
.B(n_3186),
.Y(n_5062)
);

NOR2x1_ASAP7_75t_SL g5063 ( 
.A(n_4682),
.B(n_3190),
.Y(n_5063)
);

OAI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_4888),
.A2(n_974),
.B(n_962),
.Y(n_5064)
);

OAI22xp5_ASAP7_75t_L g5065 ( 
.A1(n_4706),
.A2(n_4610),
.B1(n_4834),
.B2(n_4713),
.Y(n_5065)
);

AO22x2_ASAP7_75t_L g5066 ( 
.A1(n_4724),
.A2(n_2942),
.B1(n_2947),
.B2(n_2912),
.Y(n_5066)
);

AOI22xp33_ASAP7_75t_L g5067 ( 
.A1(n_4743),
.A2(n_2857),
.B1(n_2863),
.B2(n_2856),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_4784),
.B(n_4846),
.Y(n_5068)
);

AOI22xp5_ASAP7_75t_L g5069 ( 
.A1(n_4839),
.A2(n_2138),
.B1(n_2093),
.B2(n_3201),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_SL g5070 ( 
.A(n_4821),
.B(n_2171),
.Y(n_5070)
);

INVx5_ASAP7_75t_L g5071 ( 
.A(n_4723),
.Y(n_5071)
);

AOI21x1_ASAP7_75t_L g5072 ( 
.A1(n_4919),
.A2(n_2093),
.B(n_3201),
.Y(n_5072)
);

OAI21xp5_ASAP7_75t_L g5073 ( 
.A1(n_4715),
.A2(n_978),
.B(n_977),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4769),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_4698),
.B(n_875),
.Y(n_5075)
);

AO31x2_ASAP7_75t_L g5076 ( 
.A1(n_4795),
.A2(n_2947),
.A3(n_2950),
.B(n_2942),
.Y(n_5076)
);

OA21x2_ASAP7_75t_L g5077 ( 
.A1(n_4779),
.A2(n_981),
.B(n_980),
.Y(n_5077)
);

OAI22xp5_ASAP7_75t_L g5078 ( 
.A1(n_4766),
.A2(n_4660),
.B1(n_4694),
.B2(n_4840),
.Y(n_5078)
);

INVx4_ASAP7_75t_L g5079 ( 
.A(n_4671),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4907),
.B(n_875),
.Y(n_5080)
);

INVx5_ASAP7_75t_L g5081 ( 
.A(n_4723),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4909),
.B(n_905),
.Y(n_5082)
);

OAI21xp5_ASAP7_75t_L g5083 ( 
.A1(n_4637),
.A2(n_990),
.B(n_987),
.Y(n_5083)
);

AO31x2_ASAP7_75t_L g5084 ( 
.A1(n_4747),
.A2(n_2868),
.A3(n_2869),
.B(n_2857),
.Y(n_5084)
);

AOI22xp5_ASAP7_75t_L g5085 ( 
.A1(n_4676),
.A2(n_2138),
.B1(n_3204),
.B2(n_3202),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_L g5086 ( 
.A(n_4759),
.B(n_905),
.Y(n_5086)
);

AOI22xp5_ASAP7_75t_L g5087 ( 
.A1(n_4660),
.A2(n_2138),
.B1(n_3204),
.B2(n_3202),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4762),
.B(n_905),
.Y(n_5088)
);

OAI21x1_ASAP7_75t_L g5089 ( 
.A1(n_4726),
.A2(n_3196),
.B(n_3193),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4772),
.Y(n_5090)
);

OAI21x1_ASAP7_75t_L g5091 ( 
.A1(n_4811),
.A2(n_3209),
.B(n_3205),
.Y(n_5091)
);

AOI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4741),
.A2(n_3039),
.B(n_3018),
.Y(n_5092)
);

AND2x2_ASAP7_75t_L g5093 ( 
.A(n_4698),
.B(n_905),
.Y(n_5093)
);

CKINVDCx20_ASAP7_75t_R g5094 ( 
.A(n_4673),
.Y(n_5094)
);

NOR2xp67_ASAP7_75t_SL g5095 ( 
.A(n_4780),
.B(n_2390),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4619),
.A2(n_3039),
.B(n_3209),
.Y(n_5096)
);

OR2x6_ASAP7_75t_L g5097 ( 
.A(n_4855),
.B(n_3003),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_SL g5098 ( 
.A(n_4725),
.B(n_2171),
.Y(n_5098)
);

BUFx2_ASAP7_75t_L g5099 ( 
.A(n_4631),
.Y(n_5099)
);

OAI21x1_ASAP7_75t_L g5100 ( 
.A1(n_4647),
.A2(n_2870),
.B(n_2869),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_L g5101 ( 
.A1(n_4869),
.A2(n_2776),
.B(n_3003),
.Y(n_5101)
);

INVx3_ASAP7_75t_L g5102 ( 
.A(n_4793),
.Y(n_5102)
);

OAI22xp5_ASAP7_75t_L g5103 ( 
.A1(n_4790),
.A2(n_994),
.B1(n_995),
.B2(n_993),
.Y(n_5103)
);

AOI21xp5_ASAP7_75t_L g5104 ( 
.A1(n_4800),
.A2(n_2776),
.B(n_3004),
.Y(n_5104)
);

BUFx2_ASAP7_75t_L g5105 ( 
.A(n_4631),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_4902),
.B(n_905),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4773),
.Y(n_5107)
);

AOI21xp5_ASAP7_75t_SL g5108 ( 
.A1(n_4748),
.A2(n_1000),
.B(n_999),
.Y(n_5108)
);

NAND2xp5_ASAP7_75t_L g5109 ( 
.A(n_4801),
.B(n_905),
.Y(n_5109)
);

OAI21x1_ASAP7_75t_L g5110 ( 
.A1(n_4647),
.A2(n_2872),
.B(n_2870),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_4833),
.B(n_905),
.Y(n_5111)
);

NAND3xp33_ASAP7_75t_SL g5112 ( 
.A(n_4879),
.B(n_1009),
.C(n_1007),
.Y(n_5112)
);

OAI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_4650),
.A2(n_1017),
.B(n_1013),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4788),
.A2(n_2776),
.B(n_3004),
.Y(n_5114)
);

AOI21xp33_ASAP7_75t_L g5115 ( 
.A1(n_4914),
.A2(n_1019),
.B(n_1018),
.Y(n_5115)
);

CKINVDCx12_ASAP7_75t_R g5116 ( 
.A(n_4885),
.Y(n_5116)
);

INVx1_ASAP7_75t_SL g5117 ( 
.A(n_4826),
.Y(n_5117)
);

A2O1A1Ixp33_ASAP7_75t_L g5118 ( 
.A1(n_4797),
.A2(n_1033),
.B(n_1048),
.C(n_1020),
.Y(n_5118)
);

AOI21xp5_ASAP7_75t_L g5119 ( 
.A1(n_4783),
.A2(n_3016),
.B(n_3015),
.Y(n_5119)
);

AO31x2_ASAP7_75t_L g5120 ( 
.A1(n_4818),
.A2(n_2882),
.A3(n_2888),
.B(n_2872),
.Y(n_5120)
);

OAI21x1_ASAP7_75t_SL g5121 ( 
.A1(n_4760),
.A2(n_36),
.B(n_37),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_4807),
.B(n_905),
.Y(n_5122)
);

OR2x2_ASAP7_75t_L g5123 ( 
.A(n_4837),
.B(n_1365),
.Y(n_5123)
);

INVx4_ASAP7_75t_L g5124 ( 
.A(n_4671),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_4904),
.B(n_905),
.Y(n_5125)
);

OAI21xp5_ASAP7_75t_L g5126 ( 
.A1(n_4798),
.A2(n_1024),
.B(n_1023),
.Y(n_5126)
);

INVx4_ASAP7_75t_L g5127 ( 
.A(n_4671),
.Y(n_5127)
);

OAI22xp5_ASAP7_75t_L g5128 ( 
.A1(n_4841),
.A2(n_1028),
.B1(n_1029),
.B2(n_1025),
.Y(n_5128)
);

NAND2x1p5_ASAP7_75t_L g5129 ( 
.A(n_4780),
.B(n_2390),
.Y(n_5129)
);

BUFx6f_ASAP7_75t_L g5130 ( 
.A(n_4780),
.Y(n_5130)
);

AOI22xp5_ASAP7_75t_L g5131 ( 
.A1(n_4758),
.A2(n_2138),
.B1(n_2196),
.B2(n_2193),
.Y(n_5131)
);

OAI21x1_ASAP7_75t_SL g5132 ( 
.A1(n_4774),
.A2(n_36),
.B(n_38),
.Y(n_5132)
);

NAND2xp5_ASAP7_75t_L g5133 ( 
.A(n_4829),
.B(n_1030),
.Y(n_5133)
);

AND2x4_ASAP7_75t_L g5134 ( 
.A(n_4712),
.B(n_1365),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_4843),
.B(n_1031),
.Y(n_5135)
);

AOI21xp5_ASAP7_75t_L g5136 ( 
.A1(n_4899),
.A2(n_4911),
.B(n_4887),
.Y(n_5136)
);

NAND2xp5_ASAP7_75t_L g5137 ( 
.A(n_4847),
.B(n_1034),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4776),
.Y(n_5138)
);

AO31x2_ASAP7_75t_L g5139 ( 
.A1(n_4693),
.A2(n_2897),
.A3(n_1989),
.B(n_1993),
.Y(n_5139)
);

AOI21xp5_ASAP7_75t_L g5140 ( 
.A1(n_4887),
.A2(n_3016),
.B(n_3015),
.Y(n_5140)
);

NAND2xp5_ASAP7_75t_L g5141 ( 
.A(n_4751),
.B(n_1035),
.Y(n_5141)
);

A2O1A1Ixp33_ASAP7_75t_L g5142 ( 
.A1(n_4854),
.A2(n_1074),
.B(n_1086),
.C(n_1043),
.Y(n_5142)
);

BUFx6f_ASAP7_75t_L g5143 ( 
.A(n_4809),
.Y(n_5143)
);

AND2x4_ASAP7_75t_L g5144 ( 
.A(n_4712),
.B(n_1365),
.Y(n_5144)
);

AND2x2_ASAP7_75t_L g5145 ( 
.A(n_4736),
.B(n_38),
.Y(n_5145)
);

OAI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4868),
.A2(n_4838),
.B(n_4661),
.Y(n_5146)
);

AND2x2_ASAP7_75t_L g5147 ( 
.A(n_4736),
.B(n_39),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_4814),
.B(n_1037),
.Y(n_5148)
);

OAI21x1_ASAP7_75t_L g5149 ( 
.A1(n_4627),
.A2(n_3030),
.B(n_3019),
.Y(n_5149)
);

A2O1A1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_4652),
.A2(n_1065),
.B(n_1079),
.C(n_1050),
.Y(n_5150)
);

OAI21x1_ASAP7_75t_SL g5151 ( 
.A1(n_4620),
.A2(n_39),
.B(n_41),
.Y(n_5151)
);

NAND2xp5_ASAP7_75t_L g5152 ( 
.A(n_4730),
.B(n_1038),
.Y(n_5152)
);

AOI21xp5_ASAP7_75t_L g5153 ( 
.A1(n_4848),
.A2(n_3030),
.B(n_3019),
.Y(n_5153)
);

OAI21xp5_ASAP7_75t_SL g5154 ( 
.A1(n_4722),
.A2(n_44),
.B(n_46),
.Y(n_5154)
);

AO32x2_ASAP7_75t_L g5155 ( 
.A1(n_4687),
.A2(n_49),
.A3(n_44),
.B1(n_46),
.B2(n_51),
.Y(n_5155)
);

AND2x2_ASAP7_75t_L g5156 ( 
.A(n_4905),
.B(n_49),
.Y(n_5156)
);

NAND3xp33_ASAP7_75t_L g5157 ( 
.A(n_4838),
.B(n_1044),
.C(n_1042),
.Y(n_5157)
);

INVx1_ASAP7_75t_L g5158 ( 
.A(n_4738),
.Y(n_5158)
);

CKINVDCx20_ASAP7_75t_R g5159 ( 
.A(n_4622),
.Y(n_5159)
);

NAND2xp5_ASAP7_75t_L g5160 ( 
.A(n_4812),
.B(n_1049),
.Y(n_5160)
);

OAI21xp5_ASAP7_75t_L g5161 ( 
.A1(n_4651),
.A2(n_1053),
.B(n_1052),
.Y(n_5161)
);

OAI21x1_ASAP7_75t_SL g5162 ( 
.A1(n_4782),
.A2(n_51),
.B(n_52),
.Y(n_5162)
);

AOI211x1_ASAP7_75t_L g5163 ( 
.A1(n_4857),
.A2(n_55),
.B(n_52),
.C(n_54),
.Y(n_5163)
);

INVx2_ASAP7_75t_L g5164 ( 
.A(n_4771),
.Y(n_5164)
);

OAI22xp5_ASAP7_75t_L g5165 ( 
.A1(n_4681),
.A2(n_1059),
.B1(n_1061),
.B2(n_1055),
.Y(n_5165)
);

A2O1A1Ixp33_ASAP7_75t_L g5166 ( 
.A1(n_4683),
.A2(n_1089),
.B(n_1106),
.C(n_1072),
.Y(n_5166)
);

OA21x2_ASAP7_75t_L g5167 ( 
.A1(n_4878),
.A2(n_1066),
.B(n_1062),
.Y(n_5167)
);

AOI21xp5_ASAP7_75t_L g5168 ( 
.A1(n_4853),
.A2(n_4860),
.B(n_4822),
.Y(n_5168)
);

AO22x2_ASAP7_75t_L g5169 ( 
.A1(n_4835),
.A2(n_3035),
.B1(n_3043),
.B2(n_3041),
.Y(n_5169)
);

AND2x2_ASAP7_75t_L g5170 ( 
.A(n_4670),
.B(n_56),
.Y(n_5170)
);

OA22x2_ASAP7_75t_L g5171 ( 
.A1(n_4656),
.A2(n_1069),
.B1(n_1075),
.B2(n_1067),
.Y(n_5171)
);

OAI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_4915),
.A2(n_1078),
.B(n_1077),
.Y(n_5172)
);

AND2x2_ASAP7_75t_L g5173 ( 
.A(n_4670),
.B(n_56),
.Y(n_5173)
);

OAI21xp33_ASAP7_75t_L g5174 ( 
.A1(n_4897),
.A2(n_1083),
.B(n_1080),
.Y(n_5174)
);

AOI22xp5_ASAP7_75t_L g5175 ( 
.A1(n_4882),
.A2(n_2138),
.B1(n_2196),
.B2(n_2193),
.Y(n_5175)
);

CKINVDCx20_ASAP7_75t_R g5176 ( 
.A(n_4635),
.Y(n_5176)
);

AOI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_4916),
.A2(n_3046),
.B(n_3043),
.Y(n_5177)
);

OAI21x1_ASAP7_75t_L g5178 ( 
.A1(n_4881),
.A2(n_3047),
.B(n_3046),
.Y(n_5178)
);

NAND2xp5_ASAP7_75t_L g5179 ( 
.A(n_4817),
.B(n_1084),
.Y(n_5179)
);

AOI21xp5_ASAP7_75t_L g5180 ( 
.A1(n_4705),
.A2(n_3049),
.B(n_3047),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_4876),
.B(n_1088),
.Y(n_5181)
);

OAI21xp5_ASAP7_75t_L g5182 ( 
.A1(n_4900),
.A2(n_1095),
.B(n_1092),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_4705),
.A2(n_3049),
.B(n_2413),
.Y(n_5183)
);

NAND2xp5_ASAP7_75t_L g5184 ( 
.A(n_4918),
.B(n_1096),
.Y(n_5184)
);

OAI22xp5_ASAP7_75t_L g5185 ( 
.A1(n_4805),
.A2(n_1102),
.B1(n_1104),
.B2(n_1100),
.Y(n_5185)
);

OAI21xp5_ASAP7_75t_L g5186 ( 
.A1(n_4842),
.A2(n_1113),
.B(n_1108),
.Y(n_5186)
);

OAI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_4856),
.A2(n_1115),
.B(n_2138),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_4896),
.A2(n_2413),
.B(n_2390),
.Y(n_5188)
);

INVx2_ASAP7_75t_L g5189 ( 
.A(n_5123),
.Y(n_5189)
);

NAND2x1p5_ASAP7_75t_L g5190 ( 
.A(n_4936),
.B(n_4912),
.Y(n_5190)
);

BUFx12f_ASAP7_75t_L g5191 ( 
.A(n_4962),
.Y(n_5191)
);

BUFx8_ASAP7_75t_L g5192 ( 
.A(n_4968),
.Y(n_5192)
);

NAND2xp5_ASAP7_75t_L g5193 ( 
.A(n_4933),
.B(n_4804),
.Y(n_5193)
);

INVx2_ASAP7_75t_L g5194 ( 
.A(n_5090),
.Y(n_5194)
);

AND2x4_ASAP7_75t_L g5195 ( 
.A(n_5099),
.B(n_4682),
.Y(n_5195)
);

AO21x2_ASAP7_75t_L g5196 ( 
.A1(n_5106),
.A2(n_4893),
.B(n_4717),
.Y(n_5196)
);

OAI21xp5_ASAP7_75t_L g5197 ( 
.A1(n_4979),
.A2(n_4823),
.B(n_4870),
.Y(n_5197)
);

INVx5_ASAP7_75t_SL g5198 ( 
.A(n_5130),
.Y(n_5198)
);

AND2x2_ASAP7_75t_L g5199 ( 
.A(n_4939),
.B(n_4699),
.Y(n_5199)
);

OA21x2_ASAP7_75t_L g5200 ( 
.A1(n_4970),
.A2(n_4832),
.B(n_4892),
.Y(n_5200)
);

BUFx2_ASAP7_75t_SL g5201 ( 
.A(n_5094),
.Y(n_5201)
);

AOI21x1_ASAP7_75t_L g5202 ( 
.A1(n_4955),
.A2(n_4668),
.B(n_4645),
.Y(n_5202)
);

OAI21x1_ASAP7_75t_L g5203 ( 
.A1(n_4925),
.A2(n_4728),
.B(n_4756),
.Y(n_5203)
);

INVx2_ASAP7_75t_L g5204 ( 
.A(n_5090),
.Y(n_5204)
);

AO21x2_ASAP7_75t_L g5205 ( 
.A1(n_4961),
.A2(n_4903),
.B(n_4901),
.Y(n_5205)
);

OAI21x1_ASAP7_75t_L g5206 ( 
.A1(n_5168),
.A2(n_4757),
.B(n_4678),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5107),
.Y(n_5207)
);

BUFx2_ASAP7_75t_R g5208 ( 
.A(n_5029),
.Y(n_5208)
);

BUFx12f_ASAP7_75t_L g5209 ( 
.A(n_4983),
.Y(n_5209)
);

OA21x2_ASAP7_75t_L g5210 ( 
.A1(n_5068),
.A2(n_4824),
.B(n_4806),
.Y(n_5210)
);

INVxp67_ASAP7_75t_SL g5211 ( 
.A(n_4992),
.Y(n_5211)
);

BUFx3_ASAP7_75t_L g5212 ( 
.A(n_4947),
.Y(n_5212)
);

INVx2_ASAP7_75t_L g5213 ( 
.A(n_5107),
.Y(n_5213)
);

INVx2_ASAP7_75t_L g5214 ( 
.A(n_5138),
.Y(n_5214)
);

INVx1_ASAP7_75t_SL g5215 ( 
.A(n_4941),
.Y(n_5215)
);

CKINVDCx20_ASAP7_75t_R g5216 ( 
.A(n_5159),
.Y(n_5216)
);

BUFx5_ASAP7_75t_L g5217 ( 
.A(n_5048),
.Y(n_5217)
);

NAND2xp5_ASAP7_75t_L g5218 ( 
.A(n_4945),
.B(n_4827),
.Y(n_5218)
);

INVx3_ASAP7_75t_L g5219 ( 
.A(n_5102),
.Y(n_5219)
);

INVx2_ASAP7_75t_L g5220 ( 
.A(n_5138),
.Y(n_5220)
);

INVx1_ASAP7_75t_SL g5221 ( 
.A(n_5034),
.Y(n_5221)
);

AO21x2_ASAP7_75t_L g5222 ( 
.A1(n_5000),
.A2(n_5082),
.B(n_5080),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4937),
.A2(n_4710),
.B(n_4823),
.Y(n_5223)
);

BUFx2_ASAP7_75t_SL g5224 ( 
.A(n_4956),
.Y(n_5224)
);

HB1xp67_ASAP7_75t_L g5225 ( 
.A(n_4987),
.Y(n_5225)
);

INVx8_ASAP7_75t_L g5226 ( 
.A(n_5041),
.Y(n_5226)
);

CKINVDCx8_ASAP7_75t_R g5227 ( 
.A(n_5130),
.Y(n_5227)
);

BUFx12f_ASAP7_75t_L g5228 ( 
.A(n_4956),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_5011),
.Y(n_5229)
);

OAI21xp5_ASAP7_75t_L g5230 ( 
.A1(n_4938),
.A2(n_4870),
.B(n_4689),
.Y(n_5230)
);

INVx1_ASAP7_75t_SL g5231 ( 
.A(n_5004),
.Y(n_5231)
);

OAI21x1_ASAP7_75t_L g5232 ( 
.A1(n_4923),
.A2(n_4867),
.B(n_4690),
.Y(n_5232)
);

NAND2xp5_ASAP7_75t_L g5233 ( 
.A(n_5022),
.B(n_4873),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_5022),
.Y(n_5234)
);

AO21x2_ASAP7_75t_L g5235 ( 
.A1(n_4993),
.A2(n_4997),
.B(n_5086),
.Y(n_5235)
);

OA21x2_ASAP7_75t_L g5236 ( 
.A1(n_4989),
.A2(n_4867),
.B(n_4861),
.Y(n_5236)
);

NOR2xp33_ASAP7_75t_L g5237 ( 
.A(n_5020),
.B(n_4699),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5158),
.Y(n_5238)
);

OAI21x1_ASAP7_75t_L g5239 ( 
.A1(n_4946),
.A2(n_4867),
.B(n_4695),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_L g5240 ( 
.A(n_4922),
.B(n_4873),
.Y(n_5240)
);

OAI21xp5_ASAP7_75t_L g5241 ( 
.A1(n_5061),
.A2(n_4789),
.B(n_4815),
.Y(n_5241)
);

BUFx2_ASAP7_75t_R g5242 ( 
.A(n_4995),
.Y(n_5242)
);

INVx1_ASAP7_75t_SL g5243 ( 
.A(n_5111),
.Y(n_5243)
);

BUFx3_ASAP7_75t_L g5244 ( 
.A(n_5156),
.Y(n_5244)
);

NOR2xp33_ASAP7_75t_L g5245 ( 
.A(n_5137),
.B(n_4719),
.Y(n_5245)
);

INVxp67_ASAP7_75t_SL g5246 ( 
.A(n_4952),
.Y(n_5246)
);

AO21x2_ASAP7_75t_L g5247 ( 
.A1(n_5088),
.A2(n_5060),
.B(n_4990),
.Y(n_5247)
);

INVx3_ASAP7_75t_L g5248 ( 
.A(n_5102),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5158),
.Y(n_5249)
);

AND2x2_ASAP7_75t_L g5250 ( 
.A(n_5051),
.B(n_4719),
.Y(n_5250)
);

AOI21xp5_ASAP7_75t_L g5251 ( 
.A1(n_5114),
.A2(n_4742),
.B(n_4785),
.Y(n_5251)
);

BUFx3_ASAP7_75t_L g5252 ( 
.A(n_5145),
.Y(n_5252)
);

AO21x2_ASAP7_75t_L g5253 ( 
.A1(n_5039),
.A2(n_4828),
.B(n_4910),
.Y(n_5253)
);

AND2x4_ASAP7_75t_L g5254 ( 
.A(n_5105),
.B(n_4719),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_SL g5255 ( 
.A(n_5028),
.B(n_4729),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_4942),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5055),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_5059),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_5074),
.B(n_4729),
.Y(n_5259)
);

BUFx6f_ASAP7_75t_L g5260 ( 
.A(n_5134),
.Y(n_5260)
);

OAI21xp5_ASAP7_75t_L g5261 ( 
.A1(n_4926),
.A2(n_4913),
.B(n_4819),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5056),
.Y(n_5262)
);

BUFx3_ASAP7_75t_L g5263 ( 
.A(n_5147),
.Y(n_5263)
);

NAND2x1p5_ASAP7_75t_L g5264 ( 
.A(n_4936),
.B(n_4917),
.Y(n_5264)
);

CKINVDCx5p33_ASAP7_75t_R g5265 ( 
.A(n_5116),
.Y(n_5265)
);

NAND2x1p5_ASAP7_75t_L g5266 ( 
.A(n_4936),
.B(n_4917),
.Y(n_5266)
);

BUFx2_ASAP7_75t_SL g5267 ( 
.A(n_4973),
.Y(n_5267)
);

BUFx3_ASAP7_75t_L g5268 ( 
.A(n_5170),
.Y(n_5268)
);

BUFx2_ASAP7_75t_L g5269 ( 
.A(n_4924),
.Y(n_5269)
);

OAI21x1_ASAP7_75t_L g5270 ( 
.A1(n_4927),
.A2(n_4740),
.B(n_4734),
.Y(n_5270)
);

AND2x4_ASAP7_75t_L g5271 ( 
.A(n_5097),
.B(n_4859),
.Y(n_5271)
);

CKINVDCx5p33_ASAP7_75t_R g5272 ( 
.A(n_5028),
.Y(n_5272)
);

INVx2_ASAP7_75t_L g5273 ( 
.A(n_4934),
.Y(n_5273)
);

INVx1_ASAP7_75t_SL g5274 ( 
.A(n_4972),
.Y(n_5274)
);

INVx6_ASAP7_75t_L g5275 ( 
.A(n_5143),
.Y(n_5275)
);

BUFx12f_ASAP7_75t_L g5276 ( 
.A(n_5173),
.Y(n_5276)
);

OAI21x1_ASAP7_75t_L g5277 ( 
.A1(n_5008),
.A2(n_4792),
.B(n_4820),
.Y(n_5277)
);

INVx4_ASAP7_75t_L g5278 ( 
.A(n_5143),
.Y(n_5278)
);

BUFx12f_ASAP7_75t_L g5279 ( 
.A(n_5125),
.Y(n_5279)
);

AND2x4_ASAP7_75t_L g5280 ( 
.A(n_5097),
.B(n_5063),
.Y(n_5280)
);

INVxp67_ASAP7_75t_SL g5281 ( 
.A(n_4929),
.Y(n_5281)
);

HB1xp67_ASAP7_75t_L g5282 ( 
.A(n_4930),
.Y(n_5282)
);

CKINVDCx6p67_ASAP7_75t_R g5283 ( 
.A(n_5141),
.Y(n_5283)
);

NOR2xp67_ASAP7_75t_L g5284 ( 
.A(n_4944),
.B(n_4917),
.Y(n_5284)
);

INVx2_ASAP7_75t_L g5285 ( 
.A(n_4943),
.Y(n_5285)
);

AOI22xp33_ASAP7_75t_L g5286 ( 
.A1(n_4958),
.A2(n_4607),
.B1(n_4862),
.B2(n_4859),
.Y(n_5286)
);

BUFx2_ASAP7_75t_R g5287 ( 
.A(n_4935),
.Y(n_5287)
);

AOI22xp5_ASAP7_75t_L g5288 ( 
.A1(n_5078),
.A2(n_4607),
.B1(n_4862),
.B2(n_4836),
.Y(n_5288)
);

HB1xp67_ASAP7_75t_L g5289 ( 
.A(n_5075),
.Y(n_5289)
);

OAI21x1_ASAP7_75t_L g5290 ( 
.A1(n_4921),
.A2(n_4607),
.B(n_4862),
.Y(n_5290)
);

BUFx6f_ASAP7_75t_L g5291 ( 
.A(n_5144),
.Y(n_5291)
);

BUFx2_ASAP7_75t_SL g5292 ( 
.A(n_5176),
.Y(n_5292)
);

AOI22x1_ASAP7_75t_L g5293 ( 
.A1(n_5073),
.A2(n_4831),
.B1(n_59),
.B2(n_57),
.Y(n_5293)
);

OR2x6_ASAP7_75t_L g5294 ( 
.A(n_5136),
.B(n_4607),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5047),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5049),
.Y(n_5296)
);

OA21x2_ASAP7_75t_L g5297 ( 
.A1(n_4953),
.A2(n_1543),
.B(n_1541),
.Y(n_5297)
);

HB1xp67_ASAP7_75t_L g5298 ( 
.A(n_4949),
.Y(n_5298)
);

AOI22x1_ASAP7_75t_L g5299 ( 
.A1(n_5126),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_5299)
);

AOI22x1_ASAP7_75t_L g5300 ( 
.A1(n_4960),
.A2(n_61),
.B1(n_58),
.B2(n_60),
.Y(n_5300)
);

INVx5_ASAP7_75t_L g5301 ( 
.A(n_5052),
.Y(n_5301)
);

INVx3_ASAP7_75t_L g5302 ( 
.A(n_5079),
.Y(n_5302)
);

OA21x2_ASAP7_75t_L g5303 ( 
.A1(n_5053),
.A2(n_1543),
.B(n_1541),
.Y(n_5303)
);

OAI21x1_ASAP7_75t_L g5304 ( 
.A1(n_4940),
.A2(n_2727),
.B(n_2703),
.Y(n_5304)
);

CKINVDCx5p33_ASAP7_75t_R g5305 ( 
.A(n_5179),
.Y(n_5305)
);

OAI21x1_ASAP7_75t_L g5306 ( 
.A1(n_4948),
.A2(n_2753),
.B(n_2727),
.Y(n_5306)
);

AOI22x1_ASAP7_75t_L g5307 ( 
.A1(n_5124),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_5307)
);

OA21x2_ASAP7_75t_L g5308 ( 
.A1(n_4976),
.A2(n_1566),
.B(n_2038),
.Y(n_5308)
);

INVx2_ASAP7_75t_SL g5309 ( 
.A(n_5117),
.Y(n_5309)
);

OAI21xp5_ASAP7_75t_L g5310 ( 
.A1(n_4974),
.A2(n_626),
.B(n_609),
.Y(n_5310)
);

INVx1_ASAP7_75t_L g5311 ( 
.A(n_4957),
.Y(n_5311)
);

INVx2_ASAP7_75t_L g5312 ( 
.A(n_4975),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_4978),
.Y(n_5313)
);

NAND2x1p5_ASAP7_75t_L g5314 ( 
.A(n_4944),
.B(n_2413),
.Y(n_5314)
);

OAI21x1_ASAP7_75t_L g5315 ( 
.A1(n_5104),
.A2(n_2753),
.B(n_2727),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_4981),
.Y(n_5316)
);

NOR2xp33_ASAP7_75t_L g5317 ( 
.A(n_5154),
.B(n_63),
.Y(n_5317)
);

INVx2_ASAP7_75t_SL g5318 ( 
.A(n_5012),
.Y(n_5318)
);

NOR2xp33_ASAP7_75t_SL g5319 ( 
.A(n_5071),
.B(n_2413),
.Y(n_5319)
);

INVx5_ASAP7_75t_L g5320 ( 
.A(n_5144),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_4959),
.B(n_1365),
.Y(n_5321)
);

OAI21x1_ASAP7_75t_L g5322 ( 
.A1(n_5188),
.A2(n_2763),
.B(n_2753),
.Y(n_5322)
);

CKINVDCx20_ASAP7_75t_R g5323 ( 
.A(n_4928),
.Y(n_5323)
);

AO21x2_ASAP7_75t_L g5324 ( 
.A1(n_4982),
.A2(n_2048),
.B(n_2041),
.Y(n_5324)
);

BUFx3_ASAP7_75t_L g5325 ( 
.A(n_5181),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5018),
.B(n_1510),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_5010),
.Y(n_5327)
);

OAI21x1_ASAP7_75t_L g5328 ( 
.A1(n_5046),
.A2(n_2763),
.B(n_2050),
.Y(n_5328)
);

NAND2x1p5_ASAP7_75t_L g5329 ( 
.A(n_5071),
.B(n_5081),
.Y(n_5329)
);

INVx4_ASAP7_75t_L g5330 ( 
.A(n_5093),
.Y(n_5330)
);

OAI21x1_ASAP7_75t_L g5331 ( 
.A1(n_4951),
.A2(n_2050),
.B(n_2040),
.Y(n_5331)
);

OR2x6_ASAP7_75t_L g5332 ( 
.A(n_4931),
.B(n_2193),
.Y(n_5332)
);

AO21x2_ASAP7_75t_L g5333 ( 
.A1(n_5024),
.A2(n_2052),
.B(n_2048),
.Y(n_5333)
);

INVx2_ASAP7_75t_L g5334 ( 
.A(n_5045),
.Y(n_5334)
);

OAI21x1_ASAP7_75t_L g5335 ( 
.A1(n_5044),
.A2(n_2053),
.B(n_2040),
.Y(n_5335)
);

BUFx2_ASAP7_75t_L g5336 ( 
.A(n_5044),
.Y(n_5336)
);

INVx2_ASAP7_75t_L g5337 ( 
.A(n_5050),
.Y(n_5337)
);

AOI22x1_ASAP7_75t_L g5338 ( 
.A1(n_5124),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_5338)
);

INVx3_ASAP7_75t_L g5339 ( 
.A(n_5127),
.Y(n_5339)
);

AND2x4_ASAP7_75t_L g5340 ( 
.A(n_5081),
.B(n_5127),
.Y(n_5340)
);

BUFx6f_ASAP7_75t_L g5341 ( 
.A(n_4920),
.Y(n_5341)
);

INVx5_ASAP7_75t_L g5342 ( 
.A(n_4920),
.Y(n_5342)
);

CKINVDCx11_ASAP7_75t_R g5343 ( 
.A(n_5103),
.Y(n_5343)
);

NAND2x1p5_ASAP7_75t_L g5344 ( 
.A(n_5007),
.B(n_2578),
.Y(n_5344)
);

CKINVDCx8_ASAP7_75t_R g5345 ( 
.A(n_5023),
.Y(n_5345)
);

BUFx5_ASAP7_75t_L g5346 ( 
.A(n_4991),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5058),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_4977),
.B(n_66),
.Y(n_5348)
);

OAI21x1_ASAP7_75t_L g5349 ( 
.A1(n_5178),
.A2(n_2053),
.B(n_2040),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5169),
.Y(n_5350)
);

AOI22x1_ASAP7_75t_L g5351 ( 
.A1(n_5151),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_5351)
);

OAI21x1_ASAP7_75t_L g5352 ( 
.A1(n_5054),
.A2(n_2053),
.B(n_2052),
.Y(n_5352)
);

AOI21xp5_ASAP7_75t_L g5353 ( 
.A1(n_5108),
.A2(n_2595),
.B(n_2584),
.Y(n_5353)
);

AND2x2_ASAP7_75t_L g5354 ( 
.A(n_4949),
.B(n_69),
.Y(n_5354)
);

HB1xp67_ASAP7_75t_L g5355 ( 
.A(n_5037),
.Y(n_5355)
);

BUFx3_ASAP7_75t_L g5356 ( 
.A(n_5184),
.Y(n_5356)
);

CKINVDCx14_ASAP7_75t_R g5357 ( 
.A(n_4964),
.Y(n_5357)
);

OAI21x1_ASAP7_75t_L g5358 ( 
.A1(n_5072),
.A2(n_2053),
.B(n_2055),
.Y(n_5358)
);

BUFx12f_ASAP7_75t_L g5359 ( 
.A(n_5129),
.Y(n_5359)
);

BUFx2_ASAP7_75t_L g5360 ( 
.A(n_4966),
.Y(n_5360)
);

OAI21x1_ASAP7_75t_L g5361 ( 
.A1(n_5006),
.A2(n_2056),
.B(n_2055),
.Y(n_5361)
);

BUFx2_ASAP7_75t_R g5362 ( 
.A(n_4986),
.Y(n_5362)
);

OA21x2_ASAP7_75t_L g5363 ( 
.A1(n_5109),
.A2(n_1566),
.B(n_2056),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_5169),
.Y(n_5364)
);

INVx6_ASAP7_75t_L g5365 ( 
.A(n_4984),
.Y(n_5365)
);

INVx2_ASAP7_75t_L g5366 ( 
.A(n_5164),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_5037),
.B(n_1510),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5037),
.Y(n_5368)
);

AO21x2_ASAP7_75t_L g5369 ( 
.A1(n_5133),
.A2(n_1982),
.B(n_1158),
.Y(n_5369)
);

AOI22xp5_ASAP7_75t_L g5370 ( 
.A1(n_5065),
.A2(n_2193),
.B1(n_2205),
.B2(n_2196),
.Y(n_5370)
);

INVx2_ASAP7_75t_L g5371 ( 
.A(n_5021),
.Y(n_5371)
);

OAI21xp5_ASAP7_75t_L g5372 ( 
.A1(n_5146),
.A2(n_654),
.B(n_633),
.Y(n_5372)
);

NAND2x1p5_ASAP7_75t_L g5373 ( 
.A(n_5098),
.B(n_2584),
.Y(n_5373)
);

BUFx2_ASAP7_75t_L g5374 ( 
.A(n_5122),
.Y(n_5374)
);

OAI21x1_ASAP7_75t_L g5375 ( 
.A1(n_4963),
.A2(n_1961),
.B(n_1976),
.Y(n_5375)
);

NAND2x1p5_ASAP7_75t_L g5376 ( 
.A(n_5070),
.B(n_2584),
.Y(n_5376)
);

AO21x2_ASAP7_75t_L g5377 ( 
.A1(n_5135),
.A2(n_1158),
.B(n_1155),
.Y(n_5377)
);

INVx6_ASAP7_75t_L g5378 ( 
.A(n_5025),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_5160),
.B(n_4932),
.Y(n_5379)
);

AND2x2_ASAP7_75t_L g5380 ( 
.A(n_4932),
.B(n_70),
.Y(n_5380)
);

AO21x2_ASAP7_75t_L g5381 ( 
.A1(n_5152),
.A2(n_1196),
.B(n_1155),
.Y(n_5381)
);

INVx2_ASAP7_75t_L g5382 ( 
.A(n_5021),
.Y(n_5382)
);

BUFx2_ASAP7_75t_L g5383 ( 
.A(n_5001),
.Y(n_5383)
);

OAI21x1_ASAP7_75t_L g5384 ( 
.A1(n_5038),
.A2(n_1961),
.B(n_1976),
.Y(n_5384)
);

OAI21x1_ASAP7_75t_L g5385 ( 
.A1(n_5062),
.A2(n_1961),
.B(n_1976),
.Y(n_5385)
);

AO21x1_ASAP7_75t_L g5386 ( 
.A1(n_5128),
.A2(n_71),
.B(n_72),
.Y(n_5386)
);

AOI22x1_ASAP7_75t_L g5387 ( 
.A1(n_5121),
.A2(n_75),
.B1(n_71),
.B2(n_74),
.Y(n_5387)
);

INVx3_ASAP7_75t_SL g5388 ( 
.A(n_5171),
.Y(n_5388)
);

OAI21x1_ASAP7_75t_L g5389 ( 
.A1(n_5183),
.A2(n_1961),
.B(n_1983),
.Y(n_5389)
);

BUFx6f_ASAP7_75t_L g5390 ( 
.A(n_5155),
.Y(n_5390)
);

BUFx6f_ASAP7_75t_L g5391 ( 
.A(n_5155),
.Y(n_5391)
);

BUFx6f_ASAP7_75t_L g5392 ( 
.A(n_5155),
.Y(n_5392)
);

AND2x2_ASAP7_75t_L g5393 ( 
.A(n_4932),
.B(n_75),
.Y(n_5393)
);

INVxp67_ASAP7_75t_SL g5394 ( 
.A(n_5091),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_4985),
.Y(n_5395)
);

BUFx8_ASAP7_75t_L g5396 ( 
.A(n_5115),
.Y(n_5396)
);

AO21x2_ASAP7_75t_L g5397 ( 
.A1(n_5033),
.A2(n_1206),
.B(n_1196),
.Y(n_5397)
);

OAI21x1_ASAP7_75t_L g5398 ( 
.A1(n_4969),
.A2(n_1983),
.B(n_1211),
.Y(n_5398)
);

AOI22x1_ASAP7_75t_L g5399 ( 
.A1(n_5132),
.A2(n_79),
.B1(n_76),
.B2(n_77),
.Y(n_5399)
);

INVx4_ASAP7_75t_L g5400 ( 
.A(n_5077),
.Y(n_5400)
);

OAI21x1_ASAP7_75t_L g5401 ( 
.A1(n_5027),
.A2(n_1983),
.B(n_1211),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_4985),
.Y(n_5402)
);

OAI21x1_ASAP7_75t_L g5403 ( 
.A1(n_5005),
.A2(n_1213),
.B(n_1206),
.Y(n_5403)
);

CKINVDCx16_ASAP7_75t_R g5404 ( 
.A(n_5112),
.Y(n_5404)
);

INVx5_ASAP7_75t_L g5405 ( 
.A(n_4950),
.Y(n_5405)
);

CKINVDCx11_ASAP7_75t_R g5406 ( 
.A(n_5165),
.Y(n_5406)
);

AO21x2_ASAP7_75t_L g5407 ( 
.A1(n_5101),
.A2(n_1224),
.B(n_1213),
.Y(n_5407)
);

OAI21x1_ASAP7_75t_L g5408 ( 
.A1(n_5002),
.A2(n_1231),
.B(n_1224),
.Y(n_5408)
);

INVx2_ASAP7_75t_SL g5409 ( 
.A(n_4988),
.Y(n_5409)
);

OAI21x1_ASAP7_75t_SL g5410 ( 
.A1(n_5077),
.A2(n_76),
.B(n_79),
.Y(n_5410)
);

AOI21xp5_ASAP7_75t_L g5411 ( 
.A1(n_5236),
.A2(n_5017),
.B(n_5013),
.Y(n_5411)
);

INVx2_ASAP7_75t_SL g5412 ( 
.A(n_5226),
.Y(n_5412)
);

O2A1O1Ixp33_ASAP7_75t_L g5413 ( 
.A1(n_5310),
.A2(n_4994),
.B(n_5009),
.C(n_5030),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_SL g5414 ( 
.A(n_5272),
.B(n_5057),
.Y(n_5414)
);

OAI22xp5_ASAP7_75t_L g5415 ( 
.A1(n_5390),
.A2(n_5163),
.B1(n_5167),
.B2(n_5118),
.Y(n_5415)
);

BUFx8_ASAP7_75t_L g5416 ( 
.A(n_5228),
.Y(n_5416)
);

NAND2x1p5_ASAP7_75t_L g5417 ( 
.A(n_5255),
.B(n_5095),
.Y(n_5417)
);

AOI221xp5_ASAP7_75t_L g5418 ( 
.A1(n_5390),
.A2(n_5392),
.B1(n_5391),
.B2(n_5379),
.C(n_5354),
.Y(n_5418)
);

OAI22xp5_ASAP7_75t_L g5419 ( 
.A1(n_5391),
.A2(n_5142),
.B1(n_5085),
.B2(n_5157),
.Y(n_5419)
);

OAI21xp5_ASAP7_75t_L g5420 ( 
.A1(n_5310),
.A2(n_5064),
.B(n_5148),
.Y(n_5420)
);

OA21x2_ASAP7_75t_L g5421 ( 
.A1(n_5240),
.A2(n_5040),
.B(n_5149),
.Y(n_5421)
);

NOR2xp33_ASAP7_75t_L g5422 ( 
.A(n_5208),
.B(n_5174),
.Y(n_5422)
);

BUFx8_ASAP7_75t_L g5423 ( 
.A(n_5209),
.Y(n_5423)
);

OA21x2_ASAP7_75t_L g5424 ( 
.A1(n_5240),
.A2(n_5110),
.B(n_5100),
.Y(n_5424)
);

NOR2xp33_ASAP7_75t_L g5425 ( 
.A(n_5208),
.B(n_4998),
.Y(n_5425)
);

A2O1A1Ixp33_ASAP7_75t_L g5426 ( 
.A1(n_5391),
.A2(n_5187),
.B(n_5182),
.C(n_5113),
.Y(n_5426)
);

INVxp67_ASAP7_75t_SL g5427 ( 
.A(n_5298),
.Y(n_5427)
);

NAND2x1p5_ASAP7_75t_L g5428 ( 
.A(n_5215),
.B(n_5031),
.Y(n_5428)
);

AO21x2_ASAP7_75t_L g5429 ( 
.A1(n_5367),
.A2(n_5162),
.B(n_4980),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_5196),
.Y(n_5430)
);

INVx2_ASAP7_75t_L g5431 ( 
.A(n_5194),
.Y(n_5431)
);

OAI22xp5_ASAP7_75t_L g5432 ( 
.A1(n_5392),
.A2(n_5323),
.B1(n_5360),
.B2(n_5287),
.Y(n_5432)
);

INVx3_ASAP7_75t_L g5433 ( 
.A(n_5330),
.Y(n_5433)
);

NAND3xp33_ASAP7_75t_SL g5434 ( 
.A(n_5345),
.B(n_5069),
.C(n_5131),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5204),
.Y(n_5435)
);

BUFx2_ASAP7_75t_SL g5436 ( 
.A(n_5212),
.Y(n_5436)
);

BUFx3_ASAP7_75t_L g5437 ( 
.A(n_5192),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5207),
.Y(n_5438)
);

OAI21x1_ASAP7_75t_L g5439 ( 
.A1(n_5329),
.A2(n_5203),
.B(n_5290),
.Y(n_5439)
);

AOI221xp5_ASAP7_75t_L g5440 ( 
.A1(n_5392),
.A2(n_5172),
.B1(n_5185),
.B2(n_5186),
.C(n_5083),
.Y(n_5440)
);

AO21x2_ASAP7_75t_L g5441 ( 
.A1(n_5367),
.A2(n_5379),
.B(n_5368),
.Y(n_5441)
);

NAND3xp33_ASAP7_75t_L g5442 ( 
.A(n_5317),
.B(n_5035),
.C(n_5036),
.Y(n_5442)
);

INVx1_ASAP7_75t_L g5443 ( 
.A(n_5213),
.Y(n_5443)
);

AND2x2_ASAP7_75t_L g5444 ( 
.A(n_5199),
.B(n_5139),
.Y(n_5444)
);

O2A1O1Ixp5_ASAP7_75t_L g5445 ( 
.A1(n_5246),
.A2(n_5281),
.B(n_5400),
.C(n_5393),
.Y(n_5445)
);

A2O1A1Ixp33_ASAP7_75t_SL g5446 ( 
.A1(n_5372),
.A2(n_5016),
.B(n_5015),
.C(n_4967),
.Y(n_5446)
);

AOI221xp5_ASAP7_75t_L g5447 ( 
.A1(n_5380),
.A2(n_5161),
.B1(n_5150),
.B2(n_5166),
.C(n_4971),
.Y(n_5447)
);

AND2x4_ASAP7_75t_L g5448 ( 
.A(n_5280),
.B(n_5139),
.Y(n_5448)
);

AO31x2_ASAP7_75t_L g5449 ( 
.A1(n_5400),
.A2(n_5092),
.A3(n_5153),
.B(n_5180),
.Y(n_5449)
);

BUFx12f_ASAP7_75t_L g5450 ( 
.A(n_5192),
.Y(n_5450)
);

NAND2xp5_ASAP7_75t_L g5451 ( 
.A(n_5246),
.B(n_5281),
.Y(n_5451)
);

AND2x4_ASAP7_75t_L g5452 ( 
.A(n_5280),
.B(n_5139),
.Y(n_5452)
);

INVx1_ASAP7_75t_L g5453 ( 
.A(n_5214),
.Y(n_5453)
);

OAI21xp5_ASAP7_75t_L g5454 ( 
.A1(n_5232),
.A2(n_5043),
.B(n_5175),
.Y(n_5454)
);

INVx2_ASAP7_75t_L g5455 ( 
.A(n_5220),
.Y(n_5455)
);

AO31x2_ASAP7_75t_L g5456 ( 
.A1(n_5374),
.A2(n_5119),
.A3(n_5140),
.B(n_4965),
.Y(n_5456)
);

BUFx2_ASAP7_75t_L g5457 ( 
.A(n_5276),
.Y(n_5457)
);

INVx2_ASAP7_75t_L g5458 ( 
.A(n_5206),
.Y(n_5458)
);

AOI21xp33_ASAP7_75t_L g5459 ( 
.A1(n_5211),
.A2(n_5003),
.B(n_5087),
.Y(n_5459)
);

INVx3_ASAP7_75t_L g5460 ( 
.A(n_5254),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5229),
.Y(n_5461)
);

AOI22xp33_ASAP7_75t_SL g5462 ( 
.A1(n_5200),
.A2(n_5066),
.B1(n_5084),
.B2(n_5089),
.Y(n_5462)
);

OA21x2_ASAP7_75t_L g5463 ( 
.A1(n_5233),
.A2(n_4996),
.B(n_5026),
.Y(n_5463)
);

OAI21x1_ASAP7_75t_L g5464 ( 
.A1(n_5233),
.A2(n_5032),
.B(n_5177),
.Y(n_5464)
);

BUFx12f_ASAP7_75t_L g5465 ( 
.A(n_5265),
.Y(n_5465)
);

OA21x2_ASAP7_75t_L g5466 ( 
.A1(n_5355),
.A2(n_5218),
.B(n_5269),
.Y(n_5466)
);

NAND2xp5_ASAP7_75t_L g5467 ( 
.A(n_5282),
.B(n_5084),
.Y(n_5467)
);

INVx2_ASAP7_75t_L g5468 ( 
.A(n_5210),
.Y(n_5468)
);

AO21x2_ASAP7_75t_L g5469 ( 
.A1(n_5218),
.A2(n_5096),
.B(n_4999),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_5210),
.Y(n_5470)
);

NAND2xp5_ASAP7_75t_L g5471 ( 
.A(n_5211),
.B(n_5084),
.Y(n_5471)
);

OA21x2_ASAP7_75t_L g5472 ( 
.A1(n_5239),
.A2(n_5067),
.B(n_5042),
.Y(n_5472)
);

AOI22xp5_ASAP7_75t_L g5473 ( 
.A1(n_5370),
.A2(n_5066),
.B1(n_2193),
.B2(n_2205),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_5234),
.Y(n_5474)
);

OAI21x1_ASAP7_75t_L g5475 ( 
.A1(n_5302),
.A2(n_5120),
.B(n_5019),
.Y(n_5475)
);

OA21x2_ASAP7_75t_L g5476 ( 
.A1(n_5238),
.A2(n_5249),
.B(n_5350),
.Y(n_5476)
);

OAI21x1_ASAP7_75t_L g5477 ( 
.A1(n_5339),
.A2(n_5120),
.B(n_5019),
.Y(n_5477)
);

AOI22x1_ASAP7_75t_L g5478 ( 
.A1(n_5224),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_5478)
);

AOI21xp5_ASAP7_75t_L g5479 ( 
.A1(n_5197),
.A2(n_5019),
.B(n_5014),
.Y(n_5479)
);

OAI21x1_ASAP7_75t_L g5480 ( 
.A1(n_5339),
.A2(n_5120),
.B(n_5014),
.Y(n_5480)
);

AO31x2_ASAP7_75t_L g5481 ( 
.A1(n_5295),
.A2(n_5296),
.A3(n_5262),
.B(n_5364),
.Y(n_5481)
);

BUFx12f_ASAP7_75t_L g5482 ( 
.A(n_5396),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_5202),
.Y(n_5483)
);

OAI21x1_ASAP7_75t_L g5484 ( 
.A1(n_5190),
.A2(n_5248),
.B(n_5219),
.Y(n_5484)
);

NOR2xp33_ASAP7_75t_L g5485 ( 
.A(n_5191),
.B(n_85),
.Y(n_5485)
);

NAND2xp5_ASAP7_75t_L g5486 ( 
.A(n_5289),
.B(n_5076),
.Y(n_5486)
);

INVx3_ASAP7_75t_L g5487 ( 
.A(n_5254),
.Y(n_5487)
);

CKINVDCx20_ASAP7_75t_R g5488 ( 
.A(n_5216),
.Y(n_5488)
);

OAI21x1_ASAP7_75t_L g5489 ( 
.A1(n_5264),
.A2(n_5076),
.B(n_4954),
.Y(n_5489)
);

INVx1_ASAP7_75t_L g5490 ( 
.A(n_5256),
.Y(n_5490)
);

INVx2_ASAP7_75t_L g5491 ( 
.A(n_5189),
.Y(n_5491)
);

OAI22xp33_ASAP7_75t_L g5492 ( 
.A1(n_5370),
.A2(n_4954),
.B1(n_743),
.B2(n_763),
.Y(n_5492)
);

OAI21x1_ASAP7_75t_L g5493 ( 
.A1(n_5264),
.A2(n_2097),
.B(n_2060),
.Y(n_5493)
);

AOI21xp5_ASAP7_75t_L g5494 ( 
.A1(n_5197),
.A2(n_1512),
.B(n_1510),
.Y(n_5494)
);

AND2x4_ASAP7_75t_L g5495 ( 
.A(n_5294),
.B(n_86),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5257),
.Y(n_5496)
);

AOI21x1_ASAP7_75t_L g5497 ( 
.A1(n_5225),
.A2(n_2027),
.B(n_1988),
.Y(n_5497)
);

AOI22xp5_ASAP7_75t_L g5498 ( 
.A1(n_5241),
.A2(n_5386),
.B1(n_5267),
.B2(n_5288),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5258),
.Y(n_5499)
);

OA21x2_ASAP7_75t_L g5500 ( 
.A1(n_5394),
.A2(n_998),
.B(n_988),
.Y(n_5500)
);

AND2x4_ASAP7_75t_L g5501 ( 
.A(n_5294),
.B(n_88),
.Y(n_5501)
);

AO221x2_ASAP7_75t_L g5502 ( 
.A1(n_5241),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.C(n_92),
.Y(n_5502)
);

OAI21x1_ASAP7_75t_L g5503 ( 
.A1(n_5266),
.A2(n_2097),
.B(n_2060),
.Y(n_5503)
);

OAI21x1_ASAP7_75t_L g5504 ( 
.A1(n_5266),
.A2(n_2097),
.B(n_2060),
.Y(n_5504)
);

OA21x2_ASAP7_75t_L g5505 ( 
.A1(n_5394),
.A2(n_5402),
.B(n_5395),
.Y(n_5505)
);

OAI21x1_ASAP7_75t_SL g5506 ( 
.A1(n_5309),
.A2(n_93),
.B(n_94),
.Y(n_5506)
);

INVx2_ASAP7_75t_L g5507 ( 
.A(n_5273),
.Y(n_5507)
);

BUFx10_ASAP7_75t_L g5508 ( 
.A(n_5237),
.Y(n_5508)
);

OA21x2_ASAP7_75t_L g5509 ( 
.A1(n_5193),
.A2(n_1060),
.B(n_1003),
.Y(n_5509)
);

NOR2xp33_ASAP7_75t_L g5510 ( 
.A(n_5283),
.B(n_93),
.Y(n_5510)
);

NOR2xp33_ASAP7_75t_L g5511 ( 
.A(n_5201),
.B(n_96),
.Y(n_5511)
);

BUFx2_ASAP7_75t_L g5512 ( 
.A(n_5244),
.Y(n_5512)
);

OAI21x1_ASAP7_75t_L g5513 ( 
.A1(n_5259),
.A2(n_2087),
.B(n_2036),
.Y(n_5513)
);

OR2x2_ASAP7_75t_L g5514 ( 
.A(n_5231),
.B(n_97),
.Y(n_5514)
);

AO31x2_ASAP7_75t_L g5515 ( 
.A1(n_5245),
.A2(n_101),
.A3(n_98),
.B(n_99),
.Y(n_5515)
);

AND2x2_ASAP7_75t_L g5516 ( 
.A(n_5221),
.B(n_98),
.Y(n_5516)
);

CKINVDCx20_ASAP7_75t_R g5517 ( 
.A(n_5343),
.Y(n_5517)
);

O2A1O1Ixp33_ASAP7_75t_SL g5518 ( 
.A1(n_5215),
.A2(n_103),
.B(n_99),
.C(n_101),
.Y(n_5518)
);

OR2x6_ASAP7_75t_L g5519 ( 
.A(n_5292),
.B(n_1510),
.Y(n_5519)
);

AND2x2_ASAP7_75t_L g5520 ( 
.A(n_5250),
.B(n_105),
.Y(n_5520)
);

INVx1_ASAP7_75t_L g5521 ( 
.A(n_5321),
.Y(n_5521)
);

OR2x2_ASAP7_75t_SL g5522 ( 
.A(n_5404),
.B(n_1512),
.Y(n_5522)
);

INVx1_ASAP7_75t_SL g5523 ( 
.A(n_5287),
.Y(n_5523)
);

AOI221xp5_ASAP7_75t_L g5524 ( 
.A1(n_5410),
.A2(n_1091),
.B1(n_1512),
.B2(n_2210),
.C(n_2205),
.Y(n_5524)
);

AOI22xp33_ASAP7_75t_L g5525 ( 
.A1(n_5388),
.A2(n_2210),
.B1(n_2213),
.B2(n_2212),
.Y(n_5525)
);

OA21x2_ASAP7_75t_L g5526 ( 
.A1(n_5371),
.A2(n_2222),
.B(n_2199),
.Y(n_5526)
);

INVxp67_ASAP7_75t_SL g5527 ( 
.A(n_5297),
.Y(n_5527)
);

OAI21x1_ASAP7_75t_L g5528 ( 
.A1(n_5382),
.A2(n_106),
.B(n_107),
.Y(n_5528)
);

AND2x6_ASAP7_75t_L g5529 ( 
.A(n_5198),
.B(n_2212),
.Y(n_5529)
);

BUFx6f_ASAP7_75t_L g5530 ( 
.A(n_5344),
.Y(n_5530)
);

O2A1O1Ixp5_ASAP7_75t_L g5531 ( 
.A1(n_5195),
.A2(n_111),
.B(n_108),
.C(n_109),
.Y(n_5531)
);

OAI21xp5_ASAP7_75t_L g5532 ( 
.A1(n_5230),
.A2(n_1955),
.B(n_1952),
.Y(n_5532)
);

OAI22xp33_ASAP7_75t_L g5533 ( 
.A1(n_5332),
.A2(n_2213),
.B1(n_2219),
.B2(n_2212),
.Y(n_5533)
);

INVx1_ASAP7_75t_SL g5534 ( 
.A(n_5406),
.Y(n_5534)
);

AND2x4_ASAP7_75t_L g5535 ( 
.A(n_5243),
.B(n_111),
.Y(n_5535)
);

OA21x2_ASAP7_75t_L g5536 ( 
.A1(n_5195),
.A2(n_112),
.B(n_114),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5326),
.Y(n_5537)
);

BUFx4_ASAP7_75t_SL g5538 ( 
.A(n_5305),
.Y(n_5538)
);

OA21x2_ASAP7_75t_L g5539 ( 
.A1(n_5336),
.A2(n_114),
.B(n_116),
.Y(n_5539)
);

OAI21x1_ASAP7_75t_L g5540 ( 
.A1(n_5315),
.A2(n_117),
.B(n_118),
.Y(n_5540)
);

BUFx10_ASAP7_75t_L g5541 ( 
.A(n_5365),
.Y(n_5541)
);

CKINVDCx16_ASAP7_75t_R g5542 ( 
.A(n_5357),
.Y(n_5542)
);

INVx2_ASAP7_75t_L g5543 ( 
.A(n_5285),
.Y(n_5543)
);

NAND2x1p5_ASAP7_75t_L g5544 ( 
.A(n_5342),
.B(n_2595),
.Y(n_5544)
);

AO31x2_ASAP7_75t_L g5545 ( 
.A1(n_5251),
.A2(n_120),
.A3(n_117),
.B(n_119),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5247),
.Y(n_5546)
);

OA21x2_ASAP7_75t_L g5547 ( 
.A1(n_5311),
.A2(n_121),
.B(n_122),
.Y(n_5547)
);

INVx1_ASAP7_75t_SL g5548 ( 
.A(n_5252),
.Y(n_5548)
);

OA21x2_ASAP7_75t_L g5549 ( 
.A1(n_5316),
.A2(n_122),
.B(n_123),
.Y(n_5549)
);

CKINVDCx20_ASAP7_75t_R g5550 ( 
.A(n_5263),
.Y(n_5550)
);

NOR2xp33_ASAP7_75t_L g5551 ( 
.A(n_5268),
.B(n_128),
.Y(n_5551)
);

OAI21x1_ASAP7_75t_L g5552 ( 
.A1(n_5304),
.A2(n_130),
.B(n_132),
.Y(n_5552)
);

OAI21xp5_ASAP7_75t_L g5553 ( 
.A1(n_5270),
.A2(n_1955),
.B(n_1952),
.Y(n_5553)
);

CKINVDCx6p67_ASAP7_75t_R g5554 ( 
.A(n_5348),
.Y(n_5554)
);

OAI21x1_ASAP7_75t_L g5555 ( 
.A1(n_5306),
.A2(n_133),
.B(n_134),
.Y(n_5555)
);

BUFx6f_ASAP7_75t_L g5556 ( 
.A(n_5344),
.Y(n_5556)
);

AOI22xp33_ASAP7_75t_L g5557 ( 
.A1(n_5369),
.A2(n_2219),
.B1(n_2232),
.B2(n_2227),
.Y(n_5557)
);

AO31x2_ASAP7_75t_L g5558 ( 
.A1(n_5383),
.A2(n_136),
.A3(n_134),
.B(n_135),
.Y(n_5558)
);

OAI21x1_ASAP7_75t_L g5559 ( 
.A1(n_5314),
.A2(n_5284),
.B(n_5322),
.Y(n_5559)
);

AO31x2_ASAP7_75t_L g5560 ( 
.A1(n_5327),
.A2(n_140),
.A3(n_138),
.B(n_139),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_5274),
.Y(n_5561)
);

OAI21x1_ASAP7_75t_L g5562 ( 
.A1(n_5314),
.A2(n_138),
.B(n_139),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_5274),
.Y(n_5563)
);

OAI21x1_ASAP7_75t_L g5564 ( 
.A1(n_5284),
.A2(n_141),
.B(n_142),
.Y(n_5564)
);

OA21x2_ASAP7_75t_L g5565 ( 
.A1(n_5347),
.A2(n_142),
.B(n_143),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_5369),
.A2(n_2227),
.B1(n_2232),
.B2(n_2157),
.Y(n_5566)
);

OAI21x1_ASAP7_75t_L g5567 ( 
.A1(n_5385),
.A2(n_5313),
.B(n_5312),
.Y(n_5567)
);

OAI21x1_ASAP7_75t_L g5568 ( 
.A1(n_5334),
.A2(n_145),
.B(n_147),
.Y(n_5568)
);

OAI21x1_ASAP7_75t_L g5569 ( 
.A1(n_5337),
.A2(n_148),
.B(n_149),
.Y(n_5569)
);

BUFx6f_ASAP7_75t_L g5570 ( 
.A(n_5365),
.Y(n_5570)
);

NOR2xp33_ASAP7_75t_L g5571 ( 
.A(n_5325),
.B(n_151),
.Y(n_5571)
);

AO21x2_ASAP7_75t_L g5572 ( 
.A1(n_5247),
.A2(n_151),
.B(n_152),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_5222),
.Y(n_5573)
);

AND2x2_ASAP7_75t_L g5574 ( 
.A(n_5318),
.B(n_153),
.Y(n_5574)
);

AOI21xp5_ASAP7_75t_L g5575 ( 
.A1(n_5332),
.A2(n_2232),
.B(n_2227),
.Y(n_5575)
);

OAI22xp5_ASAP7_75t_L g5576 ( 
.A1(n_5432),
.A2(n_5242),
.B1(n_5378),
.B2(n_5362),
.Y(n_5576)
);

AO21x2_ASAP7_75t_L g5577 ( 
.A1(n_5546),
.A2(n_5381),
.B(n_5377),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_5490),
.Y(n_5578)
);

AO31x2_ASAP7_75t_L g5579 ( 
.A1(n_5430),
.A2(n_5353),
.A3(n_5278),
.B(n_5366),
.Y(n_5579)
);

BUFx2_ASAP7_75t_L g5580 ( 
.A(n_5517),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5461),
.Y(n_5581)
);

AOI21xp5_ASAP7_75t_L g5582 ( 
.A1(n_5414),
.A2(n_5353),
.B(n_5261),
.Y(n_5582)
);

OAI21x1_ASAP7_75t_L g5583 ( 
.A1(n_5445),
.A2(n_5223),
.B(n_5331),
.Y(n_5583)
);

OAI21x1_ASAP7_75t_L g5584 ( 
.A1(n_5484),
.A2(n_5389),
.B(n_5384),
.Y(n_5584)
);

OAI21xp5_ASAP7_75t_L g5585 ( 
.A1(n_5498),
.A2(n_5261),
.B(n_5387),
.Y(n_5585)
);

OAI21xp5_ASAP7_75t_L g5586 ( 
.A1(n_5426),
.A2(n_5399),
.B(n_5338),
.Y(n_5586)
);

AO21x2_ASAP7_75t_L g5587 ( 
.A1(n_5546),
.A2(n_5381),
.B(n_5377),
.Y(n_5587)
);

AOI221xp5_ASAP7_75t_L g5588 ( 
.A1(n_5418),
.A2(n_5356),
.B1(n_5253),
.B2(n_5235),
.C(n_5286),
.Y(n_5588)
);

AOI22xp33_ASAP7_75t_L g5589 ( 
.A1(n_5502),
.A2(n_5472),
.B1(n_5509),
.B2(n_5470),
.Y(n_5589)
);

AO22x2_ASAP7_75t_L g5590 ( 
.A1(n_5468),
.A2(n_5523),
.B1(n_5458),
.B2(n_5483),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5496),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5499),
.Y(n_5592)
);

AOI221x1_ASAP7_75t_L g5593 ( 
.A1(n_5573),
.A2(n_5291),
.B1(n_5260),
.B2(n_5278),
.C(n_5341),
.Y(n_5593)
);

CKINVDCx5p33_ASAP7_75t_R g5594 ( 
.A(n_5488),
.Y(n_5594)
);

OAI21x1_ASAP7_75t_L g5595 ( 
.A1(n_5460),
.A2(n_5375),
.B(n_5303),
.Y(n_5595)
);

NOR2xp33_ASAP7_75t_L g5596 ( 
.A(n_5450),
.B(n_5279),
.Y(n_5596)
);

AO21x2_ASAP7_75t_L g5597 ( 
.A1(n_5573),
.A2(n_5205),
.B(n_5277),
.Y(n_5597)
);

OA21x2_ASAP7_75t_L g5598 ( 
.A1(n_5439),
.A2(n_5340),
.B(n_5358),
.Y(n_5598)
);

OA21x2_ASAP7_75t_L g5599 ( 
.A1(n_5427),
.A2(n_5352),
.B(n_5349),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5536),
.Y(n_5600)
);

BUFx2_ASAP7_75t_L g5601 ( 
.A(n_5550),
.Y(n_5601)
);

AOI21xp5_ASAP7_75t_L g5602 ( 
.A1(n_5446),
.A2(n_5442),
.B(n_5411),
.Y(n_5602)
);

INVx1_ASAP7_75t_SL g5603 ( 
.A(n_5538),
.Y(n_5603)
);

BUFx3_ASAP7_75t_L g5604 ( 
.A(n_5465),
.Y(n_5604)
);

OAI21x1_ASAP7_75t_L g5605 ( 
.A1(n_5487),
.A2(n_5303),
.B(n_5363),
.Y(n_5605)
);

CKINVDCx20_ASAP7_75t_R g5606 ( 
.A(n_5423),
.Y(n_5606)
);

NAND2xp5_ASAP7_75t_L g5607 ( 
.A(n_5535),
.B(n_5217),
.Y(n_5607)
);

BUFx8_ASAP7_75t_L g5608 ( 
.A(n_5437),
.Y(n_5608)
);

OAI21x1_ASAP7_75t_L g5609 ( 
.A1(n_5451),
.A2(n_5363),
.B(n_5308),
.Y(n_5609)
);

OA21x2_ASAP7_75t_L g5610 ( 
.A1(n_5467),
.A2(n_5328),
.B(n_5401),
.Y(n_5610)
);

AND2x4_ASAP7_75t_L g5611 ( 
.A(n_5512),
.B(n_5320),
.Y(n_5611)
);

OA21x2_ASAP7_75t_L g5612 ( 
.A1(n_5486),
.A2(n_5361),
.B(n_5335),
.Y(n_5612)
);

INVx2_ASAP7_75t_L g5613 ( 
.A(n_5476),
.Y(n_5613)
);

NAND2xp5_ASAP7_75t_SL g5614 ( 
.A(n_5495),
.B(n_5217),
.Y(n_5614)
);

INVx1_ASAP7_75t_L g5615 ( 
.A(n_5474),
.Y(n_5615)
);

OAI21x1_ASAP7_75t_L g5616 ( 
.A1(n_5428),
.A2(n_5308),
.B(n_5373),
.Y(n_5616)
);

NAND2xp5_ASAP7_75t_L g5617 ( 
.A(n_5561),
.B(n_5291),
.Y(n_5617)
);

OAI22xp5_ASAP7_75t_L g5618 ( 
.A1(n_5501),
.A2(n_5242),
.B1(n_5378),
.B2(n_5362),
.Y(n_5618)
);

NAND2xp5_ASAP7_75t_L g5619 ( 
.A(n_5563),
.B(n_5291),
.Y(n_5619)
);

AOI21x1_ASAP7_75t_L g5620 ( 
.A1(n_5457),
.A2(n_5271),
.B(n_5398),
.Y(n_5620)
);

AOI22x1_ASAP7_75t_L g5621 ( 
.A1(n_5542),
.A2(n_5341),
.B1(n_5359),
.B2(n_5373),
.Y(n_5621)
);

OAI21x1_ASAP7_75t_L g5622 ( 
.A1(n_5466),
.A2(n_5376),
.B(n_5408),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5572),
.B(n_5301),
.Y(n_5623)
);

OAI21x1_ASAP7_75t_L g5624 ( 
.A1(n_5466),
.A2(n_5376),
.B(n_5403),
.Y(n_5624)
);

NOR2xp67_ASAP7_75t_L g5625 ( 
.A(n_5482),
.B(n_5301),
.Y(n_5625)
);

A2O1A1Ixp33_ASAP7_75t_L g5626 ( 
.A1(n_5440),
.A2(n_5422),
.B(n_5425),
.C(n_5571),
.Y(n_5626)
);

OA21x2_ASAP7_75t_L g5627 ( 
.A1(n_5471),
.A2(n_5271),
.B(n_5409),
.Y(n_5627)
);

A2O1A1Ixp33_ASAP7_75t_L g5628 ( 
.A1(n_5415),
.A2(n_5319),
.B(n_5405),
.C(n_5293),
.Y(n_5628)
);

OAI21x1_ASAP7_75t_L g5629 ( 
.A1(n_5567),
.A2(n_5346),
.B(n_5307),
.Y(n_5629)
);

AOI21xp5_ASAP7_75t_L g5630 ( 
.A1(n_5534),
.A2(n_5405),
.B(n_5351),
.Y(n_5630)
);

AO31x2_ASAP7_75t_L g5631 ( 
.A1(n_5551),
.A2(n_5346),
.A3(n_5300),
.B(n_5299),
.Y(n_5631)
);

AO31x2_ASAP7_75t_L g5632 ( 
.A1(n_5419),
.A2(n_5346),
.A3(n_5333),
.B(n_5324),
.Y(n_5632)
);

NAND2x1p5_ASAP7_75t_L g5633 ( 
.A(n_5501),
.B(n_5227),
.Y(n_5633)
);

AOI21xp5_ASAP7_75t_L g5634 ( 
.A1(n_5518),
.A2(n_5397),
.B(n_5333),
.Y(n_5634)
);

AND2x2_ASAP7_75t_L g5635 ( 
.A(n_5433),
.B(n_5275),
.Y(n_5635)
);

BUFx2_ASAP7_75t_R g5636 ( 
.A(n_5436),
.Y(n_5636)
);

OAI21x1_ASAP7_75t_L g5637 ( 
.A1(n_5433),
.A2(n_5346),
.B(n_5407),
.Y(n_5637)
);

AO21x2_ASAP7_75t_L g5638 ( 
.A1(n_5516),
.A2(n_154),
.B(n_156),
.Y(n_5638)
);

BUFx6f_ASAP7_75t_L g5639 ( 
.A(n_5570),
.Y(n_5639)
);

AO21x2_ASAP7_75t_L g5640 ( 
.A1(n_5494),
.A2(n_157),
.B(n_158),
.Y(n_5640)
);

OR2x6_ASAP7_75t_L g5641 ( 
.A(n_5519),
.B(n_2227),
.Y(n_5641)
);

OAI21x1_ASAP7_75t_SL g5642 ( 
.A1(n_5506),
.A2(n_158),
.B(n_159),
.Y(n_5642)
);

INVx1_ASAP7_75t_SL g5643 ( 
.A(n_5554),
.Y(n_5643)
);

HB1xp67_ASAP7_75t_L g5644 ( 
.A(n_5539),
.Y(n_5644)
);

NOR2xp33_ASAP7_75t_L g5645 ( 
.A(n_5416),
.B(n_159),
.Y(n_5645)
);

NOR2xp67_ASAP7_75t_L g5646 ( 
.A(n_5412),
.B(n_161),
.Y(n_5646)
);

AOI21xp5_ASAP7_75t_L g5647 ( 
.A1(n_5500),
.A2(n_162),
.B(n_163),
.Y(n_5647)
);

NOR2xp67_ASAP7_75t_SL g5648 ( 
.A(n_5570),
.B(n_2595),
.Y(n_5648)
);

INVxp67_ASAP7_75t_L g5649 ( 
.A(n_5570),
.Y(n_5649)
);

OAI22xp33_ASAP7_75t_L g5650 ( 
.A1(n_5500),
.A2(n_2232),
.B1(n_2157),
.B2(n_2070),
.Y(n_5650)
);

OA21x2_ASAP7_75t_L g5651 ( 
.A1(n_5435),
.A2(n_162),
.B(n_164),
.Y(n_5651)
);

AOI21xp5_ASAP7_75t_SL g5652 ( 
.A1(n_5547),
.A2(n_164),
.B(n_165),
.Y(n_5652)
);

AOI21xp5_ASAP7_75t_L g5653 ( 
.A1(n_5420),
.A2(n_165),
.B(n_166),
.Y(n_5653)
);

INVx1_ASAP7_75t_L g5654 ( 
.A(n_5549),
.Y(n_5654)
);

INVx1_ASAP7_75t_L g5655 ( 
.A(n_5549),
.Y(n_5655)
);

AO21x2_ASAP7_75t_L g5656 ( 
.A1(n_5521),
.A2(n_166),
.B(n_168),
.Y(n_5656)
);

INVx6_ASAP7_75t_L g5657 ( 
.A(n_5416),
.Y(n_5657)
);

NAND2xp5_ASAP7_75t_SL g5658 ( 
.A(n_5508),
.B(n_2611),
.Y(n_5658)
);

A2O1A1Ixp33_ASAP7_75t_L g5659 ( 
.A1(n_5531),
.A2(n_176),
.B(n_173),
.C(n_174),
.Y(n_5659)
);

AOI21xp5_ASAP7_75t_L g5660 ( 
.A1(n_5434),
.A2(n_174),
.B(n_177),
.Y(n_5660)
);

AOI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_5510),
.A2(n_177),
.B(n_179),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5565),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_5565),
.Y(n_5663)
);

AOI22xp33_ASAP7_75t_L g5664 ( 
.A1(n_5472),
.A2(n_2157),
.B1(n_2070),
.B2(n_2083),
.Y(n_5664)
);

OAI21x1_ASAP7_75t_L g5665 ( 
.A1(n_5464),
.A2(n_180),
.B(n_181),
.Y(n_5665)
);

AOI22xp5_ASAP7_75t_L g5666 ( 
.A1(n_5447),
.A2(n_2070),
.B1(n_2083),
.B2(n_2067),
.Y(n_5666)
);

A2O1A1Ixp33_ASAP7_75t_L g5667 ( 
.A1(n_5454),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_5667)
);

OA21x2_ASAP7_75t_L g5668 ( 
.A1(n_5438),
.A2(n_184),
.B(n_185),
.Y(n_5668)
);

AND2x4_ASAP7_75t_L g5669 ( 
.A(n_5548),
.B(n_186),
.Y(n_5669)
);

HB1xp67_ASAP7_75t_L g5670 ( 
.A(n_5505),
.Y(n_5670)
);

HB1xp67_ASAP7_75t_L g5671 ( 
.A(n_5505),
.Y(n_5671)
);

INVx6_ASAP7_75t_L g5672 ( 
.A(n_5541),
.Y(n_5672)
);

BUFx6f_ASAP7_75t_L g5673 ( 
.A(n_5564),
.Y(n_5673)
);

BUFx6f_ASAP7_75t_SL g5674 ( 
.A(n_5541),
.Y(n_5674)
);

NAND2xp5_ASAP7_75t_L g5675 ( 
.A(n_5514),
.B(n_188),
.Y(n_5675)
);

INVx2_ASAP7_75t_L g5676 ( 
.A(n_5481),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5560),
.Y(n_5677)
);

OAI21x1_ASAP7_75t_L g5678 ( 
.A1(n_5479),
.A2(n_5455),
.B(n_5431),
.Y(n_5678)
);

HB1xp67_ASAP7_75t_L g5679 ( 
.A(n_5469),
.Y(n_5679)
);

NAND2xp5_ASAP7_75t_L g5680 ( 
.A(n_5545),
.B(n_189),
.Y(n_5680)
);

BUFx6f_ASAP7_75t_L g5681 ( 
.A(n_5528),
.Y(n_5681)
);

AO21x2_ASAP7_75t_L g5682 ( 
.A1(n_5537),
.A2(n_5441),
.B(n_5497),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5537),
.Y(n_5683)
);

OAI21x1_ASAP7_75t_L g5684 ( 
.A1(n_5438),
.A2(n_191),
.B(n_192),
.Y(n_5684)
);

AOI21xp5_ASAP7_75t_L g5685 ( 
.A1(n_5429),
.A2(n_192),
.B(n_193),
.Y(n_5685)
);

INVx2_ASAP7_75t_L g5686 ( 
.A(n_5481),
.Y(n_5686)
);

AO31x2_ASAP7_75t_L g5687 ( 
.A1(n_5485),
.A2(n_197),
.A3(n_195),
.B(n_196),
.Y(n_5687)
);

AO21x2_ASAP7_75t_L g5688 ( 
.A1(n_5574),
.A2(n_195),
.B(n_196),
.Y(n_5688)
);

AOI21xp33_ASAP7_75t_SL g5689 ( 
.A1(n_5511),
.A2(n_197),
.B(n_198),
.Y(n_5689)
);

NAND2xp5_ASAP7_75t_L g5690 ( 
.A(n_5515),
.B(n_5558),
.Y(n_5690)
);

AO31x2_ASAP7_75t_L g5691 ( 
.A1(n_5443),
.A2(n_202),
.A3(n_199),
.B(n_200),
.Y(n_5691)
);

INVx1_ASAP7_75t_L g5692 ( 
.A(n_5443),
.Y(n_5692)
);

OAI21x1_ASAP7_75t_L g5693 ( 
.A1(n_5453),
.A2(n_200),
.B(n_204),
.Y(n_5693)
);

A2O1A1Ixp33_ASAP7_75t_L g5694 ( 
.A1(n_5413),
.A2(n_207),
.B(n_205),
.C(n_206),
.Y(n_5694)
);

INVx5_ASAP7_75t_L g5695 ( 
.A(n_5529),
.Y(n_5695)
);

AOI21xp5_ASAP7_75t_L g5696 ( 
.A1(n_5459),
.A2(n_208),
.B(n_209),
.Y(n_5696)
);

AND2x2_ASAP7_75t_L g5697 ( 
.A(n_5520),
.B(n_210),
.Y(n_5697)
);

INVx1_ASAP7_75t_L g5698 ( 
.A(n_5453),
.Y(n_5698)
);

NAND2xp5_ASAP7_75t_L g5699 ( 
.A(n_5463),
.B(n_210),
.Y(n_5699)
);

INVx2_ASAP7_75t_L g5700 ( 
.A(n_5507),
.Y(n_5700)
);

AOI22xp33_ASAP7_75t_L g5701 ( 
.A1(n_5444),
.A2(n_5524),
.B1(n_5525),
.B2(n_5462),
.Y(n_5701)
);

AND2x4_ASAP7_75t_L g5702 ( 
.A(n_5448),
.B(n_211),
.Y(n_5702)
);

OA21x2_ASAP7_75t_L g5703 ( 
.A1(n_5475),
.A2(n_5480),
.B(n_5477),
.Y(n_5703)
);

OAI222xp33_ASAP7_75t_L g5704 ( 
.A1(n_5473),
.A2(n_5527),
.B1(n_5491),
.B2(n_5452),
.C1(n_5543),
.C2(n_5492),
.Y(n_5704)
);

OR2x2_ASAP7_75t_L g5705 ( 
.A(n_5463),
.B(n_213),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_L g5706 ( 
.A(n_5456),
.B(n_214),
.Y(n_5706)
);

OAI21xp5_ASAP7_75t_L g5707 ( 
.A1(n_5478),
.A2(n_1955),
.B(n_1952),
.Y(n_5707)
);

AO21x2_ASAP7_75t_L g5708 ( 
.A1(n_5575),
.A2(n_215),
.B(n_218),
.Y(n_5708)
);

OAI21xp5_ASAP7_75t_L g5709 ( 
.A1(n_5478),
.A2(n_1955),
.B(n_1952),
.Y(n_5709)
);

BUFx2_ASAP7_75t_L g5710 ( 
.A(n_5417),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_5568),
.Y(n_5711)
);

INVx3_ASAP7_75t_L g5712 ( 
.A(n_5452),
.Y(n_5712)
);

INVx3_ASAP7_75t_L g5713 ( 
.A(n_5530),
.Y(n_5713)
);

AND2x2_ASAP7_75t_L g5714 ( 
.A(n_5530),
.B(n_223),
.Y(n_5714)
);

INVx1_ASAP7_75t_L g5715 ( 
.A(n_5569),
.Y(n_5715)
);

INVx1_ASAP7_75t_L g5716 ( 
.A(n_5578),
.Y(n_5716)
);

HB1xp67_ASAP7_75t_L g5717 ( 
.A(n_5670),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5651),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_5651),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_5591),
.Y(n_5720)
);

NOR2xp33_ASAP7_75t_L g5721 ( 
.A(n_5636),
.B(n_5530),
.Y(n_5721)
);

INVx4_ASAP7_75t_SL g5722 ( 
.A(n_5657),
.Y(n_5722)
);

INVx2_ASAP7_75t_SL g5723 ( 
.A(n_5580),
.Y(n_5723)
);

OR2x6_ASAP7_75t_L g5724 ( 
.A(n_5625),
.B(n_5562),
.Y(n_5724)
);

INVx1_ASAP7_75t_L g5725 ( 
.A(n_5592),
.Y(n_5725)
);

NAND2xp5_ASAP7_75t_L g5726 ( 
.A(n_5644),
.B(n_5456),
.Y(n_5726)
);

INVxp67_ASAP7_75t_SL g5727 ( 
.A(n_5699),
.Y(n_5727)
);

NOR2xp33_ASAP7_75t_L g5728 ( 
.A(n_5603),
.B(n_5556),
.Y(n_5728)
);

AOI22xp33_ASAP7_75t_L g5729 ( 
.A1(n_5589),
.A2(n_5421),
.B1(n_5553),
.B2(n_5532),
.Y(n_5729)
);

INVx2_ASAP7_75t_L g5730 ( 
.A(n_5673),
.Y(n_5730)
);

OR2x6_ASAP7_75t_L g5731 ( 
.A(n_5639),
.B(n_5540),
.Y(n_5731)
);

OA21x2_ASAP7_75t_L g5732 ( 
.A1(n_5613),
.A2(n_5489),
.B(n_5513),
.Y(n_5732)
);

OR2x6_ASAP7_75t_L g5733 ( 
.A(n_5639),
.B(n_5552),
.Y(n_5733)
);

INVx2_ASAP7_75t_L g5734 ( 
.A(n_5668),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5581),
.Y(n_5735)
);

HB1xp67_ASAP7_75t_L g5736 ( 
.A(n_5671),
.Y(n_5736)
);

CKINVDCx20_ASAP7_75t_R g5737 ( 
.A(n_5606),
.Y(n_5737)
);

AO21x2_ASAP7_75t_L g5738 ( 
.A1(n_5706),
.A2(n_5533),
.B(n_5555),
.Y(n_5738)
);

OA21x2_ASAP7_75t_L g5739 ( 
.A1(n_5602),
.A2(n_5588),
.B(n_5593),
.Y(n_5739)
);

OAI21x1_ASAP7_75t_L g5740 ( 
.A1(n_5678),
.A2(n_5559),
.B(n_5424),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5615),
.Y(n_5741)
);

INVx2_ASAP7_75t_L g5742 ( 
.A(n_5668),
.Y(n_5742)
);

HB1xp67_ASAP7_75t_L g5743 ( 
.A(n_5679),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5665),
.Y(n_5744)
);

INVx2_ASAP7_75t_L g5745 ( 
.A(n_5601),
.Y(n_5745)
);

AND2x2_ASAP7_75t_L g5746 ( 
.A(n_5635),
.B(n_5544),
.Y(n_5746)
);

INVx2_ASAP7_75t_L g5747 ( 
.A(n_5681),
.Y(n_5747)
);

NAND2x1p5_ASAP7_75t_L g5748 ( 
.A(n_5695),
.B(n_5493),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5705),
.Y(n_5749)
);

INVx2_ASAP7_75t_L g5750 ( 
.A(n_5702),
.Y(n_5750)
);

INVx3_ASAP7_75t_L g5751 ( 
.A(n_5672),
.Y(n_5751)
);

INVx1_ASAP7_75t_L g5752 ( 
.A(n_5691),
.Y(n_5752)
);

INVx1_ASAP7_75t_L g5753 ( 
.A(n_5680),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_5586),
.A2(n_5566),
.B(n_5557),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5677),
.Y(n_5755)
);

BUFx2_ASAP7_75t_L g5756 ( 
.A(n_5608),
.Y(n_5756)
);

INVx1_ASAP7_75t_L g5757 ( 
.A(n_5654),
.Y(n_5757)
);

INVx1_ASAP7_75t_L g5758 ( 
.A(n_5655),
.Y(n_5758)
);

BUFx2_ASAP7_75t_L g5759 ( 
.A(n_5608),
.Y(n_5759)
);

NAND2xp5_ASAP7_75t_L g5760 ( 
.A(n_5662),
.B(n_5449),
.Y(n_5760)
);

OAI21x1_ASAP7_75t_L g5761 ( 
.A1(n_5712),
.A2(n_5526),
.B(n_5504),
.Y(n_5761)
);

INVx1_ASAP7_75t_SL g5762 ( 
.A(n_5643),
.Y(n_5762)
);

OAI22xp33_ASAP7_75t_L g5763 ( 
.A1(n_5585),
.A2(n_5522),
.B1(n_5529),
.B2(n_5503),
.Y(n_5763)
);

AND2x4_ASAP7_75t_L g5764 ( 
.A(n_5649),
.B(n_5529),
.Y(n_5764)
);

OR2x6_ASAP7_75t_L g5765 ( 
.A(n_5685),
.B(n_5529),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5683),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_5597),
.Y(n_5767)
);

BUFx6f_ASAP7_75t_L g5768 ( 
.A(n_5604),
.Y(n_5768)
);

BUFx3_ASAP7_75t_L g5769 ( 
.A(n_5669),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5663),
.Y(n_5770)
);

BUFx2_ASAP7_75t_L g5771 ( 
.A(n_5633),
.Y(n_5771)
);

BUFx6f_ASAP7_75t_L g5772 ( 
.A(n_5714),
.Y(n_5772)
);

AOI22xp5_ASAP7_75t_L g5773 ( 
.A1(n_5653),
.A2(n_1955),
.B1(n_1952),
.B2(n_2067),
.Y(n_5773)
);

INVx3_ASAP7_75t_L g5774 ( 
.A(n_5674),
.Y(n_5774)
);

BUFx3_ASAP7_75t_L g5775 ( 
.A(n_5594),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5656),
.Y(n_5776)
);

AOI21xp5_ASAP7_75t_L g5777 ( 
.A1(n_5652),
.A2(n_224),
.B(n_225),
.Y(n_5777)
);

INVx2_ASAP7_75t_L g5778 ( 
.A(n_5627),
.Y(n_5778)
);

INVx2_ASAP7_75t_L g5779 ( 
.A(n_5703),
.Y(n_5779)
);

OAI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_5582),
.A2(n_228),
.B1(n_225),
.B2(n_226),
.Y(n_5780)
);

BUFx6f_ASAP7_75t_L g5781 ( 
.A(n_5645),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5692),
.Y(n_5782)
);

INVx1_ASAP7_75t_L g5783 ( 
.A(n_5698),
.Y(n_5783)
);

HB1xp67_ASAP7_75t_L g5784 ( 
.A(n_5682),
.Y(n_5784)
);

BUFx6f_ASAP7_75t_L g5785 ( 
.A(n_5684),
.Y(n_5785)
);

INVx2_ASAP7_75t_L g5786 ( 
.A(n_5600),
.Y(n_5786)
);

AO21x2_ASAP7_75t_L g5787 ( 
.A1(n_5676),
.A2(n_226),
.B(n_228),
.Y(n_5787)
);

NAND2xp5_ASAP7_75t_L g5788 ( 
.A(n_5590),
.B(n_229),
.Y(n_5788)
);

INVx2_ASAP7_75t_L g5789 ( 
.A(n_5686),
.Y(n_5789)
);

CKINVDCx8_ASAP7_75t_R g5790 ( 
.A(n_5596),
.Y(n_5790)
);

INVx2_ASAP7_75t_L g5791 ( 
.A(n_5687),
.Y(n_5791)
);

AOI22xp33_ASAP7_75t_L g5792 ( 
.A1(n_5690),
.A2(n_5660),
.B1(n_5638),
.B2(n_5647),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5715),
.Y(n_5793)
);

INVx2_ASAP7_75t_L g5794 ( 
.A(n_5703),
.Y(n_5794)
);

INVx1_ASAP7_75t_L g5795 ( 
.A(n_5711),
.Y(n_5795)
);

BUFx6f_ASAP7_75t_L g5796 ( 
.A(n_5693),
.Y(n_5796)
);

AND2x2_ASAP7_75t_L g5797 ( 
.A(n_5611),
.B(n_231),
.Y(n_5797)
);

AND2x2_ASAP7_75t_L g5798 ( 
.A(n_5710),
.B(n_232),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5675),
.Y(n_5799)
);

NAND2xp5_ASAP7_75t_L g5800 ( 
.A(n_5590),
.B(n_233),
.Y(n_5800)
);

INVx2_ASAP7_75t_L g5801 ( 
.A(n_5629),
.Y(n_5801)
);

INVx2_ASAP7_75t_L g5802 ( 
.A(n_5624),
.Y(n_5802)
);

INVx2_ASAP7_75t_L g5803 ( 
.A(n_5622),
.Y(n_5803)
);

INVx2_ASAP7_75t_L g5804 ( 
.A(n_5579),
.Y(n_5804)
);

INVx2_ASAP7_75t_L g5805 ( 
.A(n_5579),
.Y(n_5805)
);

CKINVDCx5p33_ASAP7_75t_R g5806 ( 
.A(n_5697),
.Y(n_5806)
);

NAND2xp5_ASAP7_75t_L g5807 ( 
.A(n_5688),
.B(n_234),
.Y(n_5807)
);

CKINVDCx20_ASAP7_75t_R g5808 ( 
.A(n_5618),
.Y(n_5808)
);

AOI22xp33_ASAP7_75t_L g5809 ( 
.A1(n_5696),
.A2(n_2108),
.B1(n_2109),
.B2(n_2096),
.Y(n_5809)
);

INVx1_ASAP7_75t_L g5810 ( 
.A(n_5623),
.Y(n_5810)
);

HB1xp67_ASAP7_75t_L g5811 ( 
.A(n_5583),
.Y(n_5811)
);

HB1xp67_ASAP7_75t_L g5812 ( 
.A(n_5598),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5617),
.Y(n_5813)
);

INVx2_ASAP7_75t_L g5814 ( 
.A(n_5632),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5619),
.Y(n_5815)
);

AOI21xp5_ASAP7_75t_L g5816 ( 
.A1(n_5667),
.A2(n_5576),
.B(n_5626),
.Y(n_5816)
);

OAI21xp5_ASAP7_75t_L g5817 ( 
.A1(n_5661),
.A2(n_235),
.B(n_236),
.Y(n_5817)
);

AOI22xp33_ASAP7_75t_SL g5818 ( 
.A1(n_5642),
.A2(n_1955),
.B1(n_1952),
.B2(n_241),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5620),
.Y(n_5819)
);

INVx1_ASAP7_75t_L g5820 ( 
.A(n_5607),
.Y(n_5820)
);

INVx1_ASAP7_75t_L g5821 ( 
.A(n_5708),
.Y(n_5821)
);

INVx2_ASAP7_75t_L g5822 ( 
.A(n_5612),
.Y(n_5822)
);

OA21x2_ASAP7_75t_L g5823 ( 
.A1(n_5704),
.A2(n_243),
.B(n_244),
.Y(n_5823)
);

OAI211xp5_ASAP7_75t_L g5824 ( 
.A1(n_5739),
.A2(n_5689),
.B(n_5694),
.C(n_5630),
.Y(n_5824)
);

AOI221xp5_ASAP7_75t_L g5825 ( 
.A1(n_5727),
.A2(n_5659),
.B1(n_5701),
.B2(n_5664),
.C(n_5666),
.Y(n_5825)
);

OAI22xp5_ASAP7_75t_L g5826 ( 
.A1(n_5808),
.A2(n_5816),
.B1(n_5806),
.B2(n_5729),
.Y(n_5826)
);

INVx2_ASAP7_75t_L g5827 ( 
.A(n_5769),
.Y(n_5827)
);

AOI22xp33_ASAP7_75t_L g5828 ( 
.A1(n_5823),
.A2(n_5640),
.B1(n_5650),
.B2(n_5700),
.Y(n_5828)
);

NAND2xp5_ASAP7_75t_L g5829 ( 
.A(n_5723),
.B(n_5646),
.Y(n_5829)
);

AOI22xp33_ASAP7_75t_L g5830 ( 
.A1(n_5718),
.A2(n_5634),
.B1(n_5587),
.B2(n_5577),
.Y(n_5830)
);

AOI21x1_ASAP7_75t_L g5831 ( 
.A1(n_5788),
.A2(n_5614),
.B(n_5658),
.Y(n_5831)
);

OR2x6_ASAP7_75t_L g5832 ( 
.A(n_5781),
.B(n_5628),
.Y(n_5832)
);

AND2x2_ASAP7_75t_L g5833 ( 
.A(n_5762),
.B(n_5745),
.Y(n_5833)
);

OAI22xp5_ASAP7_75t_SL g5834 ( 
.A1(n_5721),
.A2(n_5713),
.B1(n_5641),
.B2(n_5621),
.Y(n_5834)
);

AOI221xp5_ASAP7_75t_L g5835 ( 
.A1(n_5788),
.A2(n_5631),
.B1(n_5709),
.B2(n_5707),
.C(n_5648),
.Y(n_5835)
);

INVx3_ASAP7_75t_L g5836 ( 
.A(n_5775),
.Y(n_5836)
);

AOI22xp33_ASAP7_75t_SL g5837 ( 
.A1(n_5719),
.A2(n_5599),
.B1(n_5609),
.B2(n_5616),
.Y(n_5837)
);

AOI222xp33_ASAP7_75t_L g5838 ( 
.A1(n_5800),
.A2(n_5631),
.B1(n_5605),
.B2(n_5637),
.C1(n_5595),
.C2(n_5584),
.Y(n_5838)
);

OAI22xp5_ASAP7_75t_L g5839 ( 
.A1(n_5806),
.A2(n_5729),
.B1(n_5771),
.B2(n_5765),
.Y(n_5839)
);

OAI33xp33_ASAP7_75t_L g5840 ( 
.A1(n_5780),
.A2(n_5610),
.A3(n_5612),
.B1(n_5599),
.B2(n_249),
.B3(n_251),
.Y(n_5840)
);

OAI33xp33_ASAP7_75t_L g5841 ( 
.A1(n_5780),
.A2(n_5610),
.A3(n_249),
.B1(n_252),
.B2(n_247),
.B3(n_248),
.Y(n_5841)
);

CKINVDCx5p33_ASAP7_75t_R g5842 ( 
.A(n_5737),
.Y(n_5842)
);

OAI221xp5_ASAP7_75t_SL g5843 ( 
.A1(n_5792),
.A2(n_253),
.B1(n_250),
.B2(n_252),
.C(n_255),
.Y(n_5843)
);

INVx1_ASAP7_75t_L g5844 ( 
.A(n_5786),
.Y(n_5844)
);

OAI22xp33_ASAP7_75t_L g5845 ( 
.A1(n_5765),
.A2(n_5719),
.B1(n_5742),
.B2(n_5812),
.Y(n_5845)
);

INVx1_ASAP7_75t_L g5846 ( 
.A(n_5786),
.Y(n_5846)
);

NAND2xp5_ASAP7_75t_L g5847 ( 
.A(n_5749),
.B(n_255),
.Y(n_5847)
);

OAI21x1_ASAP7_75t_L g5848 ( 
.A1(n_5740),
.A2(n_256),
.B(n_257),
.Y(n_5848)
);

AOI221xp5_ASAP7_75t_L g5849 ( 
.A1(n_5821),
.A2(n_2112),
.B1(n_2118),
.B2(n_2110),
.C(n_2109),
.Y(n_5849)
);

NAND2xp5_ASAP7_75t_L g5850 ( 
.A(n_5799),
.B(n_256),
.Y(n_5850)
);

AOI22xp33_ASAP7_75t_SL g5851 ( 
.A1(n_5812),
.A2(n_5734),
.B1(n_5784),
.B2(n_5776),
.Y(n_5851)
);

AND2x6_ASAP7_75t_SL g5852 ( 
.A(n_5728),
.B(n_258),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5770),
.Y(n_5853)
);

INVx4_ASAP7_75t_SL g5854 ( 
.A(n_5768),
.Y(n_5854)
);

AND2x4_ASAP7_75t_L g5855 ( 
.A(n_5751),
.B(n_259),
.Y(n_5855)
);

OAI211xp5_ASAP7_75t_L g5856 ( 
.A1(n_5717),
.A2(n_265),
.B(n_261),
.C(n_264),
.Y(n_5856)
);

OAI211xp5_ASAP7_75t_L g5857 ( 
.A1(n_5717),
.A2(n_266),
.B(n_261),
.C(n_265),
.Y(n_5857)
);

INVx1_ASAP7_75t_L g5858 ( 
.A(n_5757),
.Y(n_5858)
);

OAI211xp5_ASAP7_75t_SL g5859 ( 
.A1(n_5726),
.A2(n_274),
.B(n_268),
.C(n_271),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5758),
.Y(n_5860)
);

AOI22xp5_ASAP7_75t_L g5861 ( 
.A1(n_5817),
.A2(n_2127),
.B1(n_2131),
.B2(n_2120),
.Y(n_5861)
);

INVx2_ASAP7_75t_SL g5862 ( 
.A(n_5756),
.Y(n_5862)
);

OA21x2_ASAP7_75t_L g5863 ( 
.A1(n_5767),
.A2(n_275),
.B(n_276),
.Y(n_5863)
);

OAI22xp33_ASAP7_75t_L g5864 ( 
.A1(n_5778),
.A2(n_2137),
.B1(n_2131),
.B2(n_280),
.Y(n_5864)
);

INVx2_ASAP7_75t_SL g5865 ( 
.A(n_5759),
.Y(n_5865)
);

AOI21xp5_ASAP7_75t_L g5866 ( 
.A1(n_5777),
.A2(n_278),
.B(n_279),
.Y(n_5866)
);

AOI221xp5_ASAP7_75t_L g5867 ( 
.A1(n_5753),
.A2(n_2137),
.B1(n_284),
.B2(n_282),
.C(n_283),
.Y(n_5867)
);

NOR2x1_ASAP7_75t_L g5868 ( 
.A(n_5774),
.B(n_282),
.Y(n_5868)
);

AOI21xp5_ASAP7_75t_L g5869 ( 
.A1(n_5777),
.A2(n_284),
.B(n_285),
.Y(n_5869)
);

AND2x4_ASAP7_75t_SL g5870 ( 
.A(n_5768),
.B(n_287),
.Y(n_5870)
);

INVx1_ASAP7_75t_L g5871 ( 
.A(n_5735),
.Y(n_5871)
);

OAI211xp5_ASAP7_75t_SL g5872 ( 
.A1(n_5726),
.A2(n_295),
.B(n_290),
.C(n_294),
.Y(n_5872)
);

AO21x2_ASAP7_75t_L g5873 ( 
.A1(n_5743),
.A2(n_294),
.B(n_295),
.Y(n_5873)
);

OAI211xp5_ASAP7_75t_L g5874 ( 
.A1(n_5736),
.A2(n_298),
.B(n_296),
.C(n_297),
.Y(n_5874)
);

NAND2xp5_ASAP7_75t_SL g5875 ( 
.A(n_5772),
.B(n_2611),
.Y(n_5875)
);

INVx1_ASAP7_75t_L g5876 ( 
.A(n_5741),
.Y(n_5876)
);

AOI22xp33_ASAP7_75t_L g5877 ( 
.A1(n_5791),
.A2(n_2007),
.B1(n_2025),
.B2(n_2023),
.Y(n_5877)
);

AND2x2_ASAP7_75t_L g5878 ( 
.A(n_5746),
.B(n_300),
.Y(n_5878)
);

NAND2xp5_ASAP7_75t_L g5879 ( 
.A(n_5744),
.B(n_303),
.Y(n_5879)
);

AOI22xp33_ASAP7_75t_SL g5880 ( 
.A1(n_5779),
.A2(n_307),
.B1(n_304),
.B2(n_305),
.Y(n_5880)
);

INVx1_ASAP7_75t_L g5881 ( 
.A(n_5755),
.Y(n_5881)
);

OAI21xp33_ASAP7_75t_SL g5882 ( 
.A1(n_5736),
.A2(n_305),
.B(n_308),
.Y(n_5882)
);

INVx5_ASAP7_75t_SL g5883 ( 
.A(n_5722),
.Y(n_5883)
);

OAI221xp5_ASAP7_75t_L g5884 ( 
.A1(n_5754),
.A2(n_312),
.B1(n_309),
.B2(n_310),
.C(n_313),
.Y(n_5884)
);

A2O1A1Ixp33_ASAP7_75t_L g5885 ( 
.A1(n_5817),
.A2(n_321),
.B(n_317),
.C(n_318),
.Y(n_5885)
);

INVx3_ASAP7_75t_L g5886 ( 
.A(n_5790),
.Y(n_5886)
);

OR2x2_ASAP7_75t_L g5887 ( 
.A(n_5795),
.B(n_323),
.Y(n_5887)
);

AOI22xp33_ASAP7_75t_L g5888 ( 
.A1(n_5752),
.A2(n_2030),
.B1(n_2044),
.B2(n_2035),
.Y(n_5888)
);

AOI21xp33_ASAP7_75t_L g5889 ( 
.A1(n_5801),
.A2(n_325),
.B(n_326),
.Y(n_5889)
);

OA21x2_ASAP7_75t_L g5890 ( 
.A1(n_5794),
.A2(n_5760),
.B(n_5814),
.Y(n_5890)
);

AOI221xp5_ASAP7_75t_L g5891 ( 
.A1(n_5760),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_5891)
);

OAI22xp5_ASAP7_75t_SL g5892 ( 
.A1(n_5724),
.A2(n_337),
.B1(n_332),
.B2(n_335),
.Y(n_5892)
);

INVx2_ASAP7_75t_L g5893 ( 
.A(n_5787),
.Y(n_5893)
);

OAI22xp33_ASAP7_75t_L g5894 ( 
.A1(n_5819),
.A2(n_5807),
.B1(n_5785),
.B2(n_5796),
.Y(n_5894)
);

OAI33xp33_ASAP7_75t_L g5895 ( 
.A1(n_5810),
.A2(n_337),
.A3(n_338),
.B1(n_339),
.B2(n_340),
.B3(n_342),
.Y(n_5895)
);

AND2x4_ASAP7_75t_L g5896 ( 
.A(n_5722),
.B(n_338),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5793),
.Y(n_5897)
);

AND2x2_ASAP7_75t_L g5898 ( 
.A(n_5833),
.B(n_5813),
.Y(n_5898)
);

AND2x4_ASAP7_75t_L g5899 ( 
.A(n_5862),
.B(n_5750),
.Y(n_5899)
);

BUFx3_ASAP7_75t_L g5900 ( 
.A(n_5842),
.Y(n_5900)
);

HB1xp67_ASAP7_75t_L g5901 ( 
.A(n_5873),
.Y(n_5901)
);

INVx1_ASAP7_75t_L g5902 ( 
.A(n_5844),
.Y(n_5902)
);

NAND2xp33_ASAP7_75t_R g5903 ( 
.A(n_5886),
.B(n_5807),
.Y(n_5903)
);

INVx2_ASAP7_75t_L g5904 ( 
.A(n_5863),
.Y(n_5904)
);

OR2x2_ASAP7_75t_L g5905 ( 
.A(n_5827),
.B(n_5820),
.Y(n_5905)
);

AOI22xp33_ASAP7_75t_L g5906 ( 
.A1(n_5840),
.A2(n_5796),
.B1(n_5738),
.B2(n_5822),
.Y(n_5906)
);

AND2x2_ASAP7_75t_L g5907 ( 
.A(n_5836),
.B(n_5815),
.Y(n_5907)
);

HB1xp67_ASAP7_75t_L g5908 ( 
.A(n_5882),
.Y(n_5908)
);

AND2x2_ASAP7_75t_L g5909 ( 
.A(n_5883),
.B(n_5797),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5846),
.Y(n_5910)
);

INVx2_ASAP7_75t_L g5911 ( 
.A(n_5868),
.Y(n_5911)
);

AND2x4_ASAP7_75t_L g5912 ( 
.A(n_5865),
.B(n_5854),
.Y(n_5912)
);

INVx2_ASAP7_75t_L g5913 ( 
.A(n_5852),
.Y(n_5913)
);

HB1xp67_ASAP7_75t_L g5914 ( 
.A(n_5882),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5890),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5890),
.Y(n_5916)
);

INVx2_ASAP7_75t_L g5917 ( 
.A(n_5892),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5896),
.Y(n_5918)
);

INVx3_ASAP7_75t_L g5919 ( 
.A(n_5848),
.Y(n_5919)
);

AO21x2_ASAP7_75t_L g5920 ( 
.A1(n_5894),
.A2(n_5811),
.B(n_5730),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5893),
.Y(n_5921)
);

BUFx2_ASAP7_75t_L g5922 ( 
.A(n_5829),
.Y(n_5922)
);

INVx1_ASAP7_75t_L g5923 ( 
.A(n_5879),
.Y(n_5923)
);

NAND2xp5_ASAP7_75t_L g5924 ( 
.A(n_5866),
.B(n_5869),
.Y(n_5924)
);

INVx1_ASAP7_75t_L g5925 ( 
.A(n_5847),
.Y(n_5925)
);

INVx3_ASAP7_75t_L g5926 ( 
.A(n_5831),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5897),
.Y(n_5927)
);

BUFx3_ASAP7_75t_L g5928 ( 
.A(n_5855),
.Y(n_5928)
);

INVxp67_ASAP7_75t_SL g5929 ( 
.A(n_5843),
.Y(n_5929)
);

AND2x2_ASAP7_75t_L g5930 ( 
.A(n_5878),
.B(n_5798),
.Y(n_5930)
);

INVx2_ASAP7_75t_L g5931 ( 
.A(n_5887),
.Y(n_5931)
);

AO31x2_ASAP7_75t_L g5932 ( 
.A1(n_5826),
.A2(n_5839),
.A3(n_5860),
.B(n_5858),
.Y(n_5932)
);

HB1xp67_ASAP7_75t_L g5933 ( 
.A(n_5853),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5871),
.Y(n_5934)
);

INVx2_ASAP7_75t_L g5935 ( 
.A(n_5832),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5876),
.Y(n_5936)
);

INVx2_ASAP7_75t_SL g5937 ( 
.A(n_5870),
.Y(n_5937)
);

INVx2_ASAP7_75t_L g5938 ( 
.A(n_5850),
.Y(n_5938)
);

HB1xp67_ASAP7_75t_L g5939 ( 
.A(n_5881),
.Y(n_5939)
);

AND2x2_ASAP7_75t_L g5940 ( 
.A(n_5851),
.B(n_5766),
.Y(n_5940)
);

INVx3_ASAP7_75t_L g5941 ( 
.A(n_5845),
.Y(n_5941)
);

BUFx2_ASAP7_75t_L g5942 ( 
.A(n_5834),
.Y(n_5942)
);

INVx2_ASAP7_75t_L g5943 ( 
.A(n_5884),
.Y(n_5943)
);

INVx3_ASAP7_75t_L g5944 ( 
.A(n_5824),
.Y(n_5944)
);

INVx2_ASAP7_75t_L g5945 ( 
.A(n_5875),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5838),
.B(n_5716),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5885),
.Y(n_5947)
);

AND2x4_ASAP7_75t_L g5948 ( 
.A(n_5912),
.B(n_5764),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_5944),
.B(n_5720),
.Y(n_5949)
);

INVx2_ASAP7_75t_L g5950 ( 
.A(n_5900),
.Y(n_5950)
);

OAI22xp5_ASAP7_75t_SL g5951 ( 
.A1(n_5944),
.A2(n_5880),
.B1(n_5837),
.B2(n_5828),
.Y(n_5951)
);

AND2x2_ASAP7_75t_L g5952 ( 
.A(n_5909),
.B(n_5725),
.Y(n_5952)
);

AOI22xp33_ASAP7_75t_L g5953 ( 
.A1(n_5908),
.A2(n_5825),
.B1(n_5841),
.B2(n_5830),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5901),
.Y(n_5954)
);

AOI22xp33_ASAP7_75t_SL g5955 ( 
.A1(n_5914),
.A2(n_5857),
.B1(n_5874),
.B2(n_5856),
.Y(n_5955)
);

AND2x4_ASAP7_75t_L g5956 ( 
.A(n_5928),
.B(n_5747),
.Y(n_5956)
);

NAND2xp5_ASAP7_75t_L g5957 ( 
.A(n_5915),
.B(n_5782),
.Y(n_5957)
);

INVx2_ASAP7_75t_L g5958 ( 
.A(n_5930),
.Y(n_5958)
);

NAND2xp5_ASAP7_75t_L g5959 ( 
.A(n_5916),
.B(n_5783),
.Y(n_5959)
);

AND2x2_ASAP7_75t_SL g5960 ( 
.A(n_5942),
.B(n_5835),
.Y(n_5960)
);

AOI22xp33_ASAP7_75t_L g5961 ( 
.A1(n_5924),
.A2(n_5872),
.B1(n_5859),
.B2(n_5802),
.Y(n_5961)
);

NOR2xp33_ASAP7_75t_L g5962 ( 
.A(n_5913),
.B(n_5895),
.Y(n_5962)
);

BUFx3_ASAP7_75t_L g5963 ( 
.A(n_5899),
.Y(n_5963)
);

AND2x2_ASAP7_75t_L g5964 ( 
.A(n_5898),
.B(n_5731),
.Y(n_5964)
);

HB1xp67_ASAP7_75t_L g5965 ( 
.A(n_5920),
.Y(n_5965)
);

AOI221xp5_ASAP7_75t_L g5966 ( 
.A1(n_5906),
.A2(n_5891),
.B1(n_5889),
.B2(n_5867),
.C(n_5864),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5933),
.Y(n_5967)
);

INVx1_ASAP7_75t_L g5968 ( 
.A(n_5939),
.Y(n_5968)
);

AND2x4_ASAP7_75t_L g5969 ( 
.A(n_5918),
.B(n_5733),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5939),
.Y(n_5970)
);

AND2x2_ASAP7_75t_L g5971 ( 
.A(n_5907),
.B(n_5803),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_L g5972 ( 
.A(n_5940),
.B(n_5941),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5941),
.B(n_5789),
.Y(n_5973)
);

AND2x2_ASAP7_75t_L g5974 ( 
.A(n_5922),
.B(n_5748),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_5926),
.B(n_5861),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_5926),
.B(n_5732),
.Y(n_5976)
);

NAND2x1p5_ASAP7_75t_SL g5977 ( 
.A(n_5917),
.B(n_5804),
.Y(n_5977)
);

NAND2xp5_ASAP7_75t_L g5978 ( 
.A(n_5926),
.B(n_5732),
.Y(n_5978)
);

NAND3xp33_ASAP7_75t_L g5979 ( 
.A(n_5903),
.B(n_5849),
.C(n_5809),
.Y(n_5979)
);

OR2x2_ASAP7_75t_L g5980 ( 
.A(n_5932),
.B(n_5761),
.Y(n_5980)
);

AND2x4_ASAP7_75t_L g5981 ( 
.A(n_5937),
.B(n_5805),
.Y(n_5981)
);

CKINVDCx20_ASAP7_75t_R g5982 ( 
.A(n_5937),
.Y(n_5982)
);

OAI22xp5_ASAP7_75t_L g5983 ( 
.A1(n_5906),
.A2(n_5763),
.B1(n_5818),
.B2(n_5773),
.Y(n_5983)
);

AOI22xp33_ASAP7_75t_L g5984 ( 
.A1(n_5946),
.A2(n_5904),
.B1(n_5943),
.B2(n_5929),
.Y(n_5984)
);

INVx1_ASAP7_75t_L g5985 ( 
.A(n_5931),
.Y(n_5985)
);

INVx1_ASAP7_75t_L g5986 ( 
.A(n_5965),
.Y(n_5986)
);

INVx2_ASAP7_75t_L g5987 ( 
.A(n_5963),
.Y(n_5987)
);

AND2x2_ASAP7_75t_L g5988 ( 
.A(n_5948),
.B(n_5905),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5982),
.Y(n_5989)
);

NAND2xp5_ASAP7_75t_L g5990 ( 
.A(n_5972),
.B(n_5955),
.Y(n_5990)
);

NAND4xp25_ASAP7_75t_L g5991 ( 
.A(n_5949),
.B(n_5984),
.C(n_5953),
.D(n_5950),
.Y(n_5991)
);

INVxp67_ASAP7_75t_SL g5992 ( 
.A(n_5954),
.Y(n_5992)
);

INVx2_ASAP7_75t_L g5993 ( 
.A(n_5964),
.Y(n_5993)
);

AOI22xp33_ASAP7_75t_L g5994 ( 
.A1(n_5951),
.A2(n_5911),
.B1(n_5917),
.B2(n_5947),
.Y(n_5994)
);

NAND2xp5_ASAP7_75t_L g5995 ( 
.A(n_5955),
.B(n_5925),
.Y(n_5995)
);

AND2x2_ASAP7_75t_L g5996 ( 
.A(n_5958),
.B(n_5927),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5977),
.Y(n_5997)
);

HB1xp67_ASAP7_75t_L g5998 ( 
.A(n_5949),
.Y(n_5998)
);

INVx2_ASAP7_75t_L g5999 ( 
.A(n_5980),
.Y(n_5999)
);

AND2x2_ASAP7_75t_L g6000 ( 
.A(n_5952),
.B(n_5934),
.Y(n_6000)
);

NAND2xp5_ASAP7_75t_L g6001 ( 
.A(n_5962),
.B(n_5919),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5974),
.B(n_5936),
.Y(n_6002)
);

INVx2_ASAP7_75t_L g6003 ( 
.A(n_5969),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5961),
.B(n_5919),
.Y(n_6004)
);

OAI22xp5_ASAP7_75t_L g6005 ( 
.A1(n_5951),
.A2(n_5902),
.B1(n_5910),
.B2(n_5938),
.Y(n_6005)
);

INVxp67_ASAP7_75t_L g6006 ( 
.A(n_5985),
.Y(n_6006)
);

AND2x4_ASAP7_75t_L g6007 ( 
.A(n_5956),
.B(n_5935),
.Y(n_6007)
);

INVx2_ASAP7_75t_L g6008 ( 
.A(n_5960),
.Y(n_6008)
);

OAI33xp33_ASAP7_75t_L g6009 ( 
.A1(n_6005),
.A2(n_5967),
.A3(n_5970),
.B1(n_5968),
.B2(n_5959),
.B3(n_5957),
.Y(n_6009)
);

AO21x2_ASAP7_75t_L g6010 ( 
.A1(n_5986),
.A2(n_5978),
.B(n_5976),
.Y(n_6010)
);

HB1xp67_ASAP7_75t_L g6011 ( 
.A(n_5990),
.Y(n_6011)
);

AND2x4_ASAP7_75t_L g6012 ( 
.A(n_5989),
.B(n_5981),
.Y(n_6012)
);

AOI22xp33_ASAP7_75t_L g6013 ( 
.A1(n_6008),
.A2(n_5979),
.B1(n_5966),
.B2(n_5983),
.Y(n_6013)
);

AND2x2_ASAP7_75t_L g6014 ( 
.A(n_5988),
.B(n_5971),
.Y(n_6014)
);

AOI321xp33_ASAP7_75t_L g6015 ( 
.A1(n_5994),
.A2(n_6001),
.A3(n_6008),
.B1(n_6004),
.B2(n_5997),
.C(n_5995),
.Y(n_6015)
);

HB1xp67_ASAP7_75t_L g6016 ( 
.A(n_5998),
.Y(n_6016)
);

AOI22xp33_ASAP7_75t_L g6017 ( 
.A1(n_5997),
.A2(n_5975),
.B1(n_5973),
.B2(n_5923),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_6000),
.B(n_5945),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_6007),
.Y(n_6019)
);

HB1xp67_ASAP7_75t_L g6020 ( 
.A(n_5999),
.Y(n_6020)
);

OR2x2_ASAP7_75t_L g6021 ( 
.A(n_5991),
.B(n_5921),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_6016),
.Y(n_6022)
);

INVx1_ASAP7_75t_L g6023 ( 
.A(n_6020),
.Y(n_6023)
);

AND2x4_ASAP7_75t_L g6024 ( 
.A(n_6012),
.B(n_5987),
.Y(n_6024)
);

AND2x2_ASAP7_75t_L g6025 ( 
.A(n_6014),
.B(n_6002),
.Y(n_6025)
);

INVxp67_ASAP7_75t_SL g6026 ( 
.A(n_6011),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_6019),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_6018),
.B(n_5996),
.Y(n_6028)
);

NAND2xp5_ASAP7_75t_SL g6029 ( 
.A(n_6015),
.B(n_5993),
.Y(n_6029)
);

INVx1_ASAP7_75t_L g6030 ( 
.A(n_6010),
.Y(n_6030)
);

AND2x2_ASAP7_75t_L g6031 ( 
.A(n_6028),
.B(n_6025),
.Y(n_6031)
);

INVxp67_ASAP7_75t_L g6032 ( 
.A(n_6026),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_6024),
.Y(n_6033)
);

AOI21xp5_ASAP7_75t_L g6034 ( 
.A1(n_6029),
.A2(n_5992),
.B(n_6009),
.Y(n_6034)
);

OAI22xp5_ASAP7_75t_L g6035 ( 
.A1(n_6030),
.A2(n_6013),
.B1(n_6021),
.B2(n_6017),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_6023),
.Y(n_6036)
);

INVxp67_ASAP7_75t_L g6037 ( 
.A(n_6031),
.Y(n_6037)
);

NAND2xp5_ASAP7_75t_L g6038 ( 
.A(n_6034),
.B(n_6022),
.Y(n_6038)
);

OR2x6_ASAP7_75t_L g6039 ( 
.A(n_6033),
.B(n_6027),
.Y(n_6039)
);

NAND2xp5_ASAP7_75t_L g6040 ( 
.A(n_6034),
.B(n_6006),
.Y(n_6040)
);

NAND2xp5_ASAP7_75t_L g6041 ( 
.A(n_6035),
.B(n_6017),
.Y(n_6041)
);

NOR2xp67_ASAP7_75t_L g6042 ( 
.A(n_6037),
.B(n_6032),
.Y(n_6042)
);

NOR4xp25_ASAP7_75t_L g6043 ( 
.A(n_6041),
.B(n_6015),
.C(n_6040),
.D(n_6038),
.Y(n_6043)
);

OR2x2_ASAP7_75t_L g6044 ( 
.A(n_6043),
.B(n_6039),
.Y(n_6044)
);

NAND2x1_ASAP7_75t_L g6045 ( 
.A(n_6042),
.B(n_6036),
.Y(n_6045)
);

INVx1_ASAP7_75t_SL g6046 ( 
.A(n_6044),
.Y(n_6046)
);

NOR2xp33_ASAP7_75t_L g6047 ( 
.A(n_6045),
.B(n_6003),
.Y(n_6047)
);

AOI21xp33_ASAP7_75t_L g6048 ( 
.A1(n_6044),
.A2(n_5888),
.B(n_5877),
.Y(n_6048)
);

AND2x2_ASAP7_75t_L g6049 ( 
.A(n_6047),
.B(n_349),
.Y(n_6049)
);

INVx1_ASAP7_75t_L g6050 ( 
.A(n_6048),
.Y(n_6050)
);

OAI21xp5_ASAP7_75t_L g6051 ( 
.A1(n_6046),
.A2(n_352),
.B(n_353),
.Y(n_6051)
);

OAI21xp5_ASAP7_75t_SL g6052 ( 
.A1(n_6046),
.A2(n_353),
.B(n_354),
.Y(n_6052)
);

NOR2xp33_ASAP7_75t_SL g6053 ( 
.A(n_6049),
.B(n_375),
.Y(n_6053)
);

NAND2xp5_ASAP7_75t_SL g6054 ( 
.A(n_6051),
.B(n_376),
.Y(n_6054)
);

NOR4xp25_ASAP7_75t_SL g6055 ( 
.A(n_6052),
.B(n_387),
.C(n_379),
.D(n_383),
.Y(n_6055)
);

AOI221xp5_ASAP7_75t_L g6056 ( 
.A1(n_6050),
.A2(n_394),
.B1(n_396),
.B2(n_397),
.C(n_398),
.Y(n_6056)
);

AOI22xp5_ASAP7_75t_L g6057 ( 
.A1(n_6053),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_6057)
);

AOI222xp33_ASAP7_75t_L g6058 ( 
.A1(n_6054),
.A2(n_423),
.B1(n_426),
.B2(n_430),
.C1(n_432),
.C2(n_433),
.Y(n_6058)
);

AND2x2_ASAP7_75t_L g6059 ( 
.A(n_6055),
.B(n_430),
.Y(n_6059)
);

OAI221xp5_ASAP7_75t_L g6060 ( 
.A1(n_6056),
.A2(n_438),
.B1(n_440),
.B2(n_443),
.C(n_444),
.Y(n_6060)
);

NAND2xp5_ASAP7_75t_L g6061 ( 
.A(n_6059),
.B(n_446),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_SL g6062 ( 
.A(n_6058),
.B(n_2031),
.Y(n_6062)
);

INVx1_ASAP7_75t_SL g6063 ( 
.A(n_6057),
.Y(n_6063)
);

OR2x2_ASAP7_75t_L g6064 ( 
.A(n_6061),
.B(n_6060),
.Y(n_6064)
);

OAI211xp5_ASAP7_75t_SL g6065 ( 
.A1(n_6063),
.A2(n_460),
.B(n_461),
.C(n_462),
.Y(n_6065)
);

O2A1O1Ixp5_ASAP7_75t_L g6066 ( 
.A1(n_6062),
.A2(n_465),
.B(n_466),
.C(n_467),
.Y(n_6066)
);

NOR4xp25_ASAP7_75t_L g6067 ( 
.A(n_6064),
.B(n_478),
.C(n_479),
.D(n_480),
.Y(n_6067)
);

NOR3xp33_ASAP7_75t_L g6068 ( 
.A(n_6065),
.B(n_481),
.C(n_482),
.Y(n_6068)
);

NOR3xp33_ASAP7_75t_L g6069 ( 
.A(n_6066),
.B(n_485),
.C(n_486),
.Y(n_6069)
);

NAND3xp33_ASAP7_75t_SL g6070 ( 
.A(n_6067),
.B(n_6069),
.C(n_6068),
.Y(n_6070)
);

AOI221x1_ASAP7_75t_L g6071 ( 
.A1(n_6070),
.A2(n_502),
.B1(n_503),
.B2(n_504),
.C(n_505),
.Y(n_6071)
);

INVx2_ASAP7_75t_SL g6072 ( 
.A(n_6071),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_6072),
.Y(n_6073)
);

INVx2_ASAP7_75t_L g6074 ( 
.A(n_6072),
.Y(n_6074)
);

INVx2_ASAP7_75t_L g6075 ( 
.A(n_6073),
.Y(n_6075)
);

HB1xp67_ASAP7_75t_L g6076 ( 
.A(n_6074),
.Y(n_6076)
);

AO22x2_ASAP7_75t_L g6077 ( 
.A1(n_6075),
.A2(n_511),
.B1(n_512),
.B2(n_514),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_6076),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_6078),
.Y(n_6079)
);

INVx2_ASAP7_75t_L g6080 ( 
.A(n_6079),
.Y(n_6080)
);

INVx2_ASAP7_75t_L g6081 ( 
.A(n_6079),
.Y(n_6081)
);

NAND2x1_ASAP7_75t_L g6082 ( 
.A(n_6079),
.B(n_6077),
.Y(n_6082)
);

INVx3_ASAP7_75t_L g6083 ( 
.A(n_6080),
.Y(n_6083)
);

INVx1_ASAP7_75t_L g6084 ( 
.A(n_6081),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_6083),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_6084),
.B(n_6082),
.Y(n_6086)
);

HB1xp67_ASAP7_75t_L g6087 ( 
.A(n_6085),
.Y(n_6087)
);

AOI22xp5_ASAP7_75t_L g6088 ( 
.A1(n_6086),
.A2(n_2175),
.B1(n_533),
.B2(n_534),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_6087),
.Y(n_6089)
);

OAI22xp5_ASAP7_75t_L g6090 ( 
.A1(n_6089),
.A2(n_6088),
.B1(n_536),
.B2(n_540),
.Y(n_6090)
);

INVx2_ASAP7_75t_L g6091 ( 
.A(n_6089),
.Y(n_6091)
);

O2A1O1Ixp33_ASAP7_75t_L g6092 ( 
.A1(n_6089),
.A2(n_535),
.B(n_540),
.C(n_541),
.Y(n_6092)
);

AOI221xp5_ASAP7_75t_L g6093 ( 
.A1(n_6091),
.A2(n_545),
.B1(n_546),
.B2(n_548),
.C(n_549),
.Y(n_6093)
);

AOI221xp5_ASAP7_75t_L g6094 ( 
.A1(n_6092),
.A2(n_549),
.B1(n_550),
.B2(n_551),
.C(n_552),
.Y(n_6094)
);

OAI21xp5_ASAP7_75t_L g6095 ( 
.A1(n_6090),
.A2(n_550),
.B(n_552),
.Y(n_6095)
);

NAND2xp5_ASAP7_75t_SL g6096 ( 
.A(n_6094),
.B(n_2035),
.Y(n_6096)
);

OAI22xp33_ASAP7_75t_L g6097 ( 
.A1(n_6096),
.A2(n_6095),
.B1(n_6093),
.B2(n_556),
.Y(n_6097)
);

OA21x2_ASAP7_75t_L g6098 ( 
.A1(n_6097),
.A2(n_557),
.B(n_561),
.Y(n_6098)
);

OAI22xp5_ASAP7_75t_L g6099 ( 
.A1(n_6097),
.A2(n_2044),
.B1(n_2046),
.B2(n_1997),
.Y(n_6099)
);

INVx1_ASAP7_75t_L g6100 ( 
.A(n_6098),
.Y(n_6100)
);

AOI22xp5_ASAP7_75t_SL g6101 ( 
.A1(n_6099),
.A2(n_562),
.B1(n_563),
.B2(n_564),
.Y(n_6101)
);

AOI22xp33_ASAP7_75t_L g6102 ( 
.A1(n_6098),
.A2(n_2046),
.B1(n_1999),
.B2(n_566),
.Y(n_6102)
);

OR2x2_ASAP7_75t_L g6103 ( 
.A(n_6100),
.B(n_564),
.Y(n_6103)
);

AO21x1_ASAP7_75t_L g6104 ( 
.A1(n_6102),
.A2(n_6101),
.B(n_568),
.Y(n_6104)
);

OAI21xp5_ASAP7_75t_L g6105 ( 
.A1(n_6100),
.A2(n_567),
.B(n_571),
.Y(n_6105)
);

AOI22xp5_ASAP7_75t_L g6106 ( 
.A1(n_6104),
.A2(n_1999),
.B1(n_2719),
.B2(n_2672),
.Y(n_6106)
);

AOI22xp33_ASAP7_75t_SL g6107 ( 
.A1(n_6103),
.A2(n_572),
.B1(n_575),
.B2(n_578),
.Y(n_6107)
);

AOI22xp33_ASAP7_75t_L g6108 ( 
.A1(n_6106),
.A2(n_6105),
.B1(n_583),
.B2(n_584),
.Y(n_6108)
);

AOI211xp5_ASAP7_75t_L g6109 ( 
.A1(n_6108),
.A2(n_6107),
.B(n_590),
.C(n_592),
.Y(n_6109)
);


endmodule