module fake_jpeg_17511_n_331 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_13),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_16),
.Y(n_86)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_11),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_16),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_23),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_88),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_70),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_32),
.B1(n_26),
.B2(n_15),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_75),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_31),
.Y(n_82)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_29),
.B(n_24),
.C(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_25),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_29),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_86),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_15),
.B1(n_19),
.B2(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_97),
.B1(n_105),
.B2(n_20),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_18),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_28),
.B1(n_19),
.B2(n_21),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_28),
.B1(n_19),
.B2(n_23),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_72),
.B1(n_103),
.B2(n_112),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_41),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_23),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_17),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_101),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_41),
.B(n_21),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_45),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_37),
.B(n_17),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_37),
.B(n_17),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_114),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_37),
.B(n_11),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_41),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_126),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_118),
.A2(n_133),
.B1(n_150),
.B2(n_106),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_119),
.B(n_165),
.Y(n_183)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_20),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_128),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_67),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_132),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_140),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_135),
.A2(n_161),
.B1(n_136),
.B2(n_144),
.Y(n_203)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_25),
.B1(n_9),
.B2(n_3),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_175)
);

OAI211xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_92),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_94),
.Y(n_180)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

AO22x1_ASAP7_75t_SL g147 ( 
.A1(n_83),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_100),
.B(n_5),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_94),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_162),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_70),
.A2(n_6),
.B1(n_8),
.B2(n_115),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_90),
.A2(n_6),
.B1(n_103),
.B2(n_110),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_93),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_155),
.B(n_163),
.Y(n_196)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_67),
.B1(n_84),
.B2(n_77),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_164),
.B1(n_131),
.B2(n_112),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_70),
.B(n_69),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_116),
.B1(n_87),
.B2(n_97),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_95),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_77),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_84),
.A2(n_76),
.B1(n_106),
.B2(n_110),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_109),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_167),
.B(n_190),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_142),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_168),
.B(n_172),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_146),
.Y(n_170)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_123),
.B(n_76),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_176),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_148),
.B(n_135),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_201),
.B1(n_148),
.B2(n_161),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_199),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_122),
.B(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_188),
.B(n_185),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_125),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_142),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_187),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_124),
.B(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_195),
.B(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_127),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_126),
.B(n_117),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g201 ( 
.A1(n_118),
.A2(n_119),
.B1(n_161),
.B2(n_135),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_156),
.B1(n_154),
.B2(n_139),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_184),
.B1(n_173),
.B2(n_203),
.Y(n_229)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_203),
.A2(n_192),
.B(n_175),
.Y(n_233)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_142),
.C(n_129),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_151),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_208),
.A2(n_212),
.B1(n_218),
.B2(n_221),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_201),
.A2(n_183),
.B(n_172),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_208),
.B(n_239),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_201),
.A2(n_133),
.B1(n_147),
.B2(n_141),
.Y(n_212)
);

AO21x1_ASAP7_75t_L g265 ( 
.A1(n_213),
.A2(n_233),
.B(n_214),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_217),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_147),
.B1(n_149),
.B2(n_135),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_128),
.B1(n_145),
.B2(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_193),
.B1(n_168),
.B2(n_171),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_230),
.Y(n_247)
);

AND2x6_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_180),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_226),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_170),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_229),
.A2(n_221),
.B(n_236),
.C(n_219),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_191),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_179),
.A2(n_197),
.B1(n_204),
.B2(n_170),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_166),
.B(n_177),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_171),
.A2(n_175),
.B1(n_197),
.B2(n_194),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_177),
.B(n_186),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_178),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_228),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_242),
.B(n_240),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_233),
.A2(n_176),
.B1(n_185),
.B2(n_194),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_213),
.A2(n_227),
.B(n_239),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_251),
.A2(n_256),
.B(n_258),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_211),
.A2(n_220),
.B(n_218),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_224),
.C(n_219),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_210),
.A2(n_223),
.B(n_222),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_245),
.B1(n_244),
.B2(n_243),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_209),
.A2(n_216),
.B(n_241),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_262),
.A2(n_253),
.B(n_260),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_242),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_258),
.B1(n_261),
.B2(n_265),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_262),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_265),
.A2(n_246),
.B1(n_245),
.B2(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_266),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_269),
.B(n_286),
.Y(n_292)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_248),
.Y(n_273)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_248),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_276),
.B(n_277),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_264),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_280),
.A2(n_282),
.B1(n_271),
.B2(n_279),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_259),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_281),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_261),
.B1(n_249),
.B2(n_257),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_284),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_267),
.B1(n_244),
.B2(n_243),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_289),
.Y(n_302)
);

OA21x2_ASAP7_75t_SL g290 ( 
.A1(n_269),
.A2(n_285),
.B(n_279),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_SL g304 ( 
.A(n_290),
.B(n_270),
.C(n_275),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_300),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_272),
.B(n_276),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_296),
.B1(n_298),
.B2(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_274),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_300),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g312 ( 
.A(n_306),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_308),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_291),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_288),
.A2(n_301),
.B1(n_292),
.B2(n_289),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_311),
.B1(n_309),
.B2(n_302),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_297),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_291),
.B1(n_294),
.B2(n_298),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_307),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_293),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_305),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_317),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_309),
.C(n_314),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_324),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_325),
.A2(n_321),
.B(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_327),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_312),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_313),
.Y(n_331)
);


endmodule