module fake_jpeg_6774_n_17 (n_3, n_2, n_1, n_0, n_4, n_17);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_17;

wire n_13;
wire n_11;
wire n_14;
wire n_16;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_5;
wire n_7;

AND2x2_ASAP7_75t_L g5 ( 
.A(n_2),
.B(n_1),
.Y(n_5)
);

AOI22xp33_ASAP7_75t_L g6 ( 
.A1(n_3),
.A2(n_1),
.B1(n_0),
.B2(n_4),
.Y(n_6)
);

CKINVDCx9p33_ASAP7_75t_R g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

MAJx2_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_4),
.C(n_2),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_9),
.B(n_10),
.C(n_8),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_3),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g11 ( 
.A1(n_5),
.A2(n_0),
.B(n_2),
.Y(n_11)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_11),
.A2(n_12),
.B(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_7),
.B(n_0),
.Y(n_12)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_14),
.C(n_15),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_8),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_14),
.B(n_8),
.Y(n_17)
);


endmodule