module real_jpeg_20092_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_0),
.A2(n_41),
.B1(n_49),
.B2(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_0),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_1),
.B(n_38),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_1),
.A2(n_14),
.B(n_28),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_1),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_1),
.A2(n_30),
.B1(n_128),
.B2(n_129),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_1),
.B(n_144),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_38),
.B(n_100),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_59),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_147)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_4),
.A2(n_26),
.B(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_4),
.A2(n_104),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_85),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_8),
.A2(n_55),
.B1(n_56),
.B2(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_55),
.B1(n_56),
.B2(n_76),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_76),
.Y(n_116)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_14),
.A2(n_55),
.B(n_80),
.C(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_14),
.B(n_55),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_14),
.Y(n_82)
);

INVx11_ASAP7_75t_SL g57 ( 
.A(n_15),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_107),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_106),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_90),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_20),
.B(n_90),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_68),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_29),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_30),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_30),
.A2(n_114),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_30),
.A2(n_116),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_31),
.B(n_66),
.Y(n_105)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_31),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_31),
.B(n_43),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_41),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_41),
.B(n_44),
.C(n_62),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_51),
.Y(n_53)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI32xp33_ASAP7_75t_L g99 ( 
.A1(n_39),
.A2(n_52),
.A3(n_55),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_62),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_43),
.CON(n_40),
.SN(n_40)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_61),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_43),
.A2(n_56),
.B(n_82),
.C(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_43),
.B(n_81),
.Y(n_131)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_60),
.C(n_63),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_47),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_58),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_48),
.A2(n_50),
.B1(n_54),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_54),
.B1(n_58),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_51),
.B(n_56),
.Y(n_101)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_54),
.Y(n_144)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_89),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_83),
.B(n_86),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_79),
.A2(n_81),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_79),
.A2(n_81),
.B1(n_124),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_79),
.A2(n_81),
.B1(n_96),
.B2(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_98),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_91),
.A2(n_92),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_95),
.B(n_98),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_102),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_130),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_164),
.B(n_169),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_151),
.B(n_163),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_138),
.B(n_150),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_125),
.B(n_137),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_117),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_117),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_132),
.B(n_136),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_131),
.Y(n_136)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_146),
.C(n_148),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_153),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_161),
.B2(n_162),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_154),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_156),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);


endmodule