module fake_jpeg_27130_n_192 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_1),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_49),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g50 ( 
.A1(n_17),
.A2(n_1),
.B(n_2),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_19),
.B(n_18),
.C(n_4),
.Y(n_68)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_34),
.B1(n_31),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_23),
.B1(n_27),
.B2(n_26),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_6),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_23),
.B(n_27),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_68),
.B(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_26),
.B1(n_25),
.B2(n_20),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_24),
.B1(n_32),
.B2(n_25),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_65),
.B1(n_73),
.B2(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_46),
.A2(n_20),
.B1(n_19),
.B2(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_10),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_37),
.A2(n_24),
.B1(n_32),
.B2(n_22),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_71),
.B1(n_69),
.B2(n_66),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_37),
.A2(n_22),
.B1(n_32),
.B2(n_4),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_37),
.A2(n_22),
.B1(n_3),
.B2(n_5),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_6),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_9),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_53),
.Y(n_106)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_85),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_83),
.A2(n_92),
.B1(n_82),
.B2(n_85),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_7),
.C(n_8),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_87),
.C(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_76),
.B(n_13),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_10),
.B1(n_11),
.B2(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_100),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_75),
.B(n_54),
.C(n_60),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_98),
.A2(n_101),
.B1(n_55),
.B2(n_77),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_75),
.B(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_72),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_55),
.B(n_59),
.C(n_72),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_112),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_77),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_122),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_77),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_118),
.B1(n_80),
.B2(n_91),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_102),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_95),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_123),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_122),
.B1(n_105),
.B2(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_134),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_95),
.B(n_86),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

NOR4xp25_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_90),
.C(n_92),
.D(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_131),
.C(n_133),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_120),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_101),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_78),
.C(n_79),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_96),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_114),
.B1(n_115),
.B2(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_113),
.B1(n_116),
.B2(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_138),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_154),
.B1(n_139),
.B2(n_140),
.Y(n_164)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_153),
.B(n_155),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_118),
.B1(n_107),
.B2(n_122),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_155),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_131),
.B(n_134),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_161),
.B(n_110),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_163),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_128),
.C(n_135),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_166),
.C(n_149),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_133),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_164),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_129),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_139),
.B1(n_125),
.B2(n_137),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_117),
.C(n_110),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_170),
.B(n_172),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_162),
.A2(n_146),
.B(n_141),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_143),
.B(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_143),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_180),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_161),
.B(n_164),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_171),
.C(n_157),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_142),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_159),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_166),
.C(n_142),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_183),
.A2(n_175),
.A3(n_145),
.B1(n_156),
.B2(n_172),
.C1(n_158),
.C2(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_182),
.C(n_184),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_188),
.B(n_160),
.Y(n_191)
);

FAx1_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_189),
.CI(n_148),
.CON(n_192),
.SN(n_192)
);


endmodule