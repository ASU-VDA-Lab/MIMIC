module fake_jpeg_1284_n_122 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_48),
.Y(n_56)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_49),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_37),
.B1(n_36),
.B2(n_40),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_41),
.B1(n_38),
.B2(n_33),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_45),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_36),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_40),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_77),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_59),
.B1(n_58),
.B2(n_32),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_79),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_8),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_2),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_62),
.B(n_4),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_4),
.B(n_5),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_85),
.B(n_15),
.Y(n_105)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_89),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_5),
.B(n_6),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

NOR3xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_92),
.C(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_6),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_94),
.Y(n_95)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_9),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_97),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_9),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_10),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_102),
.B(n_105),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_12),
.B(n_13),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_14),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_95),
.C(n_104),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_103),
.Y(n_112)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_91),
.A3(n_17),
.B1(n_18),
.B2(n_19),
.C1(n_20),
.C2(n_22),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_101),
.B(n_29),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_30),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_113),
.Y(n_116)
);

NOR2xp67_ASAP7_75t_SL g115 ( 
.A(n_114),
.B(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_116),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_107),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_110),
.C(n_26),
.Y(n_122)
);


endmodule