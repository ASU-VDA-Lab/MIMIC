module fake_jpeg_4504_n_141 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_141);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_0),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_29),
.B(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_15),
.Y(n_39)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_27),
.B1(n_28),
.B2(n_21),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_25),
.Y(n_60)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_31),
.B(n_23),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_29),
.B(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_19),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_28),
.B1(n_27),
.B2(n_37),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_15),
.B1(n_19),
.B2(n_24),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_21),
.B1(n_37),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_13),
.B1(n_20),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_13),
.B1(n_17),
.B2(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_61),
.B1(n_11),
.B2(n_3),
.Y(n_84)
);

OR2x4_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_36),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_63),
.Y(n_88)
);

OA22x2_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_36),
.B1(n_33),
.B2(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_65),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_64),
.B1(n_72),
.B2(n_45),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_33),
.B1(n_38),
.B2(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_33),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_22),
.B1(n_24),
.B2(n_16),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_84),
.B1(n_61),
.B2(n_53),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_38),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_32),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_32),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_86),
.Y(n_93)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_89),
.B(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_102),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_59),
.B1(n_58),
.B2(n_52),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_59),
.B1(n_62),
.B2(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_99),
.B(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_66),
.B1(n_32),
.B2(n_18),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_99),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_16),
.B(n_3),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_16),
.B1(n_63),
.B2(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_105),
.B(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_111),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_98),
.A2(n_77),
.B1(n_85),
.B2(n_86),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_110),
.A2(n_85),
.B(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_110),
.B(n_93),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_112),
.C(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_118),
.C(n_119),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_2),
.Y(n_125)
);

OAI322xp33_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_100),
.A3(n_97),
.B1(n_77),
.B2(n_93),
.C1(n_74),
.C2(n_8),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_77),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_104),
.B1(n_4),
.B2(n_5),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_126),
.Y(n_128)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_114),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_113),
.B(n_116),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_9),
.B(n_131),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_113),
.C(n_119),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_8),
.Y(n_133)
);

OAI321xp33_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_122),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_6),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_134),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_135),
.C(n_127),
.Y(n_136)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_128),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_138),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_137),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_134),
.Y(n_141)
);


endmodule