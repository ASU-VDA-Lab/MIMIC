module fake_jpeg_16585_n_138 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_138);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_1),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_68),
.B(n_48),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_55),
.CON(n_69),
.SN(n_69)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_73),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_60),
.A2(n_55),
.B1(n_45),
.B2(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_74),
.B1(n_78),
.B2(n_80),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_46),
.B1(n_58),
.B2(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_52),
.B1(n_42),
.B2(n_51),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_58),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_2),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_56),
.B1(n_54),
.B2(n_44),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_54),
.B1(n_43),
.B2(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_60),
.A2(n_57),
.B1(n_48),
.B2(n_3),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_82),
.B(n_83),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_1),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_90),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_67),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_7),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_6),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_67),
.B1(n_76),
.B2(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_98),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_106),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_27),
.B1(n_40),
.B2(n_39),
.Y(n_105)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_87),
.B1(n_98),
.B2(n_97),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_115),
.B1(n_116),
.B2(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_114),
.B1(n_107),
.B2(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g115 ( 
.A1(n_103),
.A2(n_93),
.B1(n_88),
.B2(n_86),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_89),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_100),
.C(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_119),
.B(n_112),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_120),
.B(n_121),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_125),
.B1(n_118),
.B2(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_122),
.A2(n_115),
.B1(n_119),
.B2(n_110),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_127),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_93),
.C(n_28),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_128),
.C(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_128),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_25),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_24),
.B(n_38),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_18),
.A3(n_37),
.B1(n_36),
.B2(n_34),
.C1(n_12),
.C2(n_13),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_17),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_29),
.C(n_33),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_16),
.A3(n_31),
.B1(n_30),
.B2(n_41),
.C(n_11),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_8),
.Y(n_138)
);


endmodule