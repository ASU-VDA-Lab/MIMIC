module real_aes_7614_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_635;
wire n_357;
wire n_792;
wire n_673;
wire n_386;
wire n_503;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_1014;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_742;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_948;
wire n_399;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_816;
wire n_539;
wire n_400;
wire n_626;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_994;
wire n_372;
wire n_495;
wire n_892;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_940;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_999;
wire n_913;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_1003;
wire n_533;
wire n_1000;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_749;
wire n_385;
wire n_358;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_691;
wire n_481;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_0), .A2(n_148), .B1(n_581), .B2(n_999), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_1), .B(n_569), .Y(n_655) );
XOR2x2_ASAP7_75t_L g623 ( .A(n_2), .B(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_3), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_4), .A2(n_258), .B1(n_721), .B2(n_757), .Y(n_756) );
OA22x2_ASAP7_75t_L g791 ( .A1(n_5), .A2(n_792), .B1(n_793), .B2(n_816), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_5), .Y(n_792) );
OA22x2_ASAP7_75t_L g739 ( .A1(n_6), .A2(n_740), .B1(n_741), .B2(n_764), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_6), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_7), .A2(n_76), .B1(n_473), .B2(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_8), .A2(n_246), .B1(n_450), .B2(n_534), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_9), .A2(n_305), .B1(n_461), .B2(n_475), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_10), .Y(n_391) );
AO22x2_ASAP7_75t_L g358 ( .A1(n_11), .A2(n_183), .B1(n_359), .B2(n_360), .Y(n_358) );
INVx1_ASAP7_75t_L g978 ( .A(n_11), .Y(n_978) );
AOI22xp5_ASAP7_75t_SL g580 ( .A1(n_12), .A2(n_332), .B1(n_420), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_13), .A2(n_173), .B1(n_628), .B2(n_887), .Y(n_886) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_14), .A2(n_260), .B1(n_381), .B2(n_599), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_15), .A2(n_54), .B1(n_751), .B2(n_948), .Y(n_947) );
AOI22xp5_ASAP7_75t_SL g575 ( .A1(n_16), .A2(n_206), .B1(n_406), .B2(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_17), .A2(n_93), .B1(n_402), .B2(n_773), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_18), .A2(n_23), .B1(n_534), .B2(n_778), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_19), .A2(n_334), .B1(n_422), .B2(n_479), .Y(n_893) );
CKINVDCx20_ASAP7_75t_R g833 ( .A(n_20), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_21), .Y(n_872) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_22), .A2(n_324), .B1(n_426), .B2(n_509), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_24), .A2(n_225), .B1(n_462), .B2(n_613), .Y(n_832) );
INVx1_ASAP7_75t_L g639 ( .A(n_25), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_26), .A2(n_318), .B1(n_509), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_27), .A2(n_149), .B1(n_572), .B2(n_573), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_28), .A2(n_295), .B1(n_510), .B2(n_665), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_29), .A2(n_87), .B1(n_382), .B2(n_444), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g959 ( .A1(n_30), .A2(n_48), .B1(n_512), .B2(n_538), .Y(n_959) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_31), .Y(n_753) );
AO22x2_ASAP7_75t_L g362 ( .A1(n_32), .A2(n_98), .B1(n_359), .B2(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_33), .A2(n_220), .B1(n_684), .B2(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_34), .A2(n_167), .B1(n_686), .B2(n_724), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_35), .A2(n_237), .B1(n_605), .B2(n_773), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_36), .A2(n_214), .B1(n_528), .B2(n_601), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_37), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g597 ( .A1(n_38), .A2(n_290), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g1000 ( .A1(n_39), .A2(n_283), .B1(n_468), .B2(n_689), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_40), .A2(n_188), .B1(n_519), .B2(n_520), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_41), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g820 ( .A1(n_42), .A2(n_232), .B1(n_431), .B2(n_467), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_43), .B(n_601), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_44), .B(n_449), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_45), .A2(n_227), .B1(n_375), .B2(n_449), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g989 ( .A1(n_46), .A2(n_164), .B1(n_449), .B2(n_563), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_47), .A2(n_125), .B1(n_406), .B2(n_413), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_49), .B(n_385), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g844 ( .A(n_50), .Y(n_844) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_51), .A2(n_288), .B1(n_473), .B2(n_502), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_52), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_53), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_55), .A2(n_319), .B1(n_462), .B2(n_471), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_56), .A2(n_255), .B1(n_523), .B2(n_613), .Y(n_659) );
AOI22xp5_ASAP7_75t_SL g482 ( .A1(n_57), .A2(n_483), .B1(n_513), .B2(n_514), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_57), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_58), .A2(n_174), .B1(n_478), .B2(n_583), .Y(n_864) );
INVx1_ASAP7_75t_L g585 ( .A(n_59), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_60), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_61), .Y(n_498) );
AOI222xp33_ASAP7_75t_L g541 ( .A1(n_62), .A2(n_170), .B1(n_199), .B2(n_542), .C1(n_543), .C2(n_544), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_63), .A2(n_66), .B1(n_607), .B2(n_609), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_64), .A2(n_229), .B1(n_426), .B2(n_584), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_65), .A2(n_91), .B1(n_584), .B2(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_67), .A2(n_127), .B1(n_505), .B2(n_523), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_68), .A2(n_215), .B1(n_376), .B2(n_532), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_69), .A2(n_195), .B1(n_402), .B2(n_519), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_70), .A2(n_201), .B1(n_430), .B2(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_SL g577 ( .A1(n_71), .A2(n_212), .B1(n_413), .B2(n_578), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g952 ( .A1(n_72), .A2(n_189), .B1(n_444), .B2(n_953), .Y(n_952) );
OA22x2_ASAP7_75t_L g586 ( .A1(n_73), .A2(n_587), .B1(n_588), .B2(n_617), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_73), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_74), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_75), .A2(n_210), .B1(n_426), .B2(n_463), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g511 ( .A1(n_77), .A2(n_111), .B1(n_413), .B2(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_78), .A2(n_239), .B1(n_523), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_79), .A2(n_262), .B1(n_422), .B2(n_522), .Y(n_884) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_80), .A2(n_181), .B1(n_689), .B2(n_691), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_81), .A2(n_101), .B1(n_406), .B2(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g824 ( .A(n_82), .Y(n_824) );
AO22x2_ASAP7_75t_L g366 ( .A1(n_83), .A2(n_219), .B1(n_359), .B2(n_360), .Y(n_366) );
INVx1_ASAP7_75t_L g975 ( .A(n_83), .Y(n_975) );
CKINVDCx20_ASAP7_75t_R g811 ( .A(n_84), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_85), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_86), .A2(n_88), .B1(n_684), .B2(n_686), .Y(n_683) );
AOI22xp5_ASAP7_75t_SL g582 ( .A1(n_89), .A2(n_177), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_90), .A2(n_256), .B1(n_512), .B2(n_540), .Y(n_539) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_92), .A2(n_336), .B(n_344), .C(n_980), .Y(n_335) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_94), .Y(n_933) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_95), .A2(n_168), .B1(n_776), .B2(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_96), .A2(n_100), .B1(n_543), .B2(n_544), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_97), .A2(n_150), .B1(n_532), .B2(n_808), .Y(n_901) );
INVx1_ASAP7_75t_L g979 ( .A(n_98), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_99), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_102), .A2(n_291), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_103), .A2(n_166), .B1(n_502), .B2(n_1003), .Y(n_1002) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_104), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_105), .B(n_528), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_106), .A2(n_176), .B1(n_994), .B2(n_995), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_107), .A2(n_202), .B1(n_583), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g611 ( .A1(n_108), .A2(n_230), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_109), .A2(n_122), .B1(n_375), .B2(n_381), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g956 ( .A1(n_110), .A2(n_156), .B1(n_605), .B2(n_860), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_112), .A2(n_292), .B1(n_512), .B2(n_721), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_113), .A2(n_203), .B1(n_444), .B2(n_532), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_114), .A2(n_209), .B1(n_598), .B2(n_599), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_115), .A2(n_321), .B1(n_726), .B2(n_728), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_116), .A2(n_300), .B1(n_381), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_SL g802 ( .A1(n_117), .A2(n_172), .B1(n_465), .B2(n_691), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g614 ( .A1(n_118), .A2(n_133), .B1(n_402), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_119), .A2(n_158), .B1(n_528), .B2(n_776), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_120), .A2(n_316), .B1(n_475), .B2(n_478), .Y(n_474) );
XNOR2x2_ASAP7_75t_L g765 ( .A(n_121), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g666 ( .A(n_123), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_124), .B(n_569), .Y(n_828) );
AND2x6_ASAP7_75t_L g338 ( .A(n_126), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g972 ( .A(n_126), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_128), .A2(n_323), .B1(n_420), .B2(n_422), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_129), .A2(n_157), .B1(n_502), .B2(n_663), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_130), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g992 ( .A(n_131), .B(n_527), .Y(n_992) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_132), .A2(n_306), .B1(n_426), .B2(n_430), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_134), .A2(n_160), .B1(n_505), .B2(n_605), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g991 ( .A(n_135), .B(n_601), .Y(n_991) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_136), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_137), .A2(n_151), .B1(n_663), .B2(n_904), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_138), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_139), .B(n_654), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_140), .Y(n_879) );
AOI222xp33_ASAP7_75t_L g780 ( .A1(n_141), .A2(n_175), .B1(n_296), .B2(n_385), .C1(n_781), .C2(n_782), .Y(n_780) );
AO22x2_ASAP7_75t_L g368 ( .A1(n_142), .A2(n_211), .B1(n_359), .B2(n_363), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g976 ( .A(n_142), .B(n_977), .Y(n_976) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_143), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_144), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_145), .A2(n_250), .B1(n_428), .B2(n_477), .Y(n_831) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_146), .A2(n_153), .B1(n_461), .B2(n_463), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_147), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_152), .A2(n_221), .B1(n_462), .B2(n_512), .Y(n_905) );
AOI22xp33_ASAP7_75t_SL g464 ( .A1(n_154), .A2(n_281), .B1(n_465), .B2(n_468), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_155), .A2(n_274), .B1(n_478), .B2(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_159), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_161), .Y(n_874) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_162), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_163), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_165), .A2(n_261), .B1(n_540), .B2(n_616), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_169), .A2(n_259), .B1(n_720), .B2(n_721), .Y(n_719) );
XOR2xp5_ASAP7_75t_L g981 ( .A(n_171), .B(n_982), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_178), .A2(n_200), .B1(n_402), .B2(n_406), .Y(n_401) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_179), .A2(n_194), .B1(n_409), .B2(n_413), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_180), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_182), .A2(n_198), .B1(n_422), .B2(n_616), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_184), .B(n_527), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_185), .A2(n_311), .B1(n_381), .B2(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_186), .A2(n_224), .B1(n_510), .B2(n_665), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_187), .A2(n_231), .B1(n_493), .B2(n_749), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g861 ( .A1(n_190), .A2(n_263), .B1(n_721), .B2(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_191), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_192), .A2(n_315), .B1(n_504), .B2(n_505), .Y(n_503) );
OA22x2_ASAP7_75t_L g347 ( .A1(n_193), .A2(n_348), .B1(n_349), .B2(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_193), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_196), .A2(n_213), .B1(n_522), .B2(n_523), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_197), .A2(n_285), .B1(n_520), .B2(n_686), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_204), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_205), .Y(n_561) );
INVx2_ASAP7_75t_L g343 ( .A(n_207), .Y(n_343) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_208), .A2(n_254), .B1(n_523), .B2(n_665), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_216), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_217), .Y(n_708) );
XNOR2x1_ASAP7_75t_L g942 ( .A(n_218), .B(n_943), .Y(n_942) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_222), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g871 ( .A(n_223), .Y(n_871) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_226), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_228), .Y(n_745) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_233), .A2(n_252), .B1(n_471), .B2(n_473), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_234), .Y(n_940) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_235), .Y(n_918) );
AOI22x1_ASAP7_75t_L g700 ( .A1(n_236), .A2(n_701), .B1(n_729), .B2(n_730), .Y(n_700) );
INVx1_ASAP7_75t_L g729 ( .A(n_236), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_238), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_240), .Y(n_854) );
OA22x2_ASAP7_75t_L g910 ( .A1(n_241), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
CKINVDCx16_ASAP7_75t_R g911 ( .A(n_241), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_242), .B(n_527), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_243), .A2(n_308), .B1(n_413), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g359 ( .A(n_244), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_244), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_245), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_247), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_248), .A2(n_294), .B1(n_540), .B2(n_862), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_249), .Y(n_592) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_251), .A2(n_286), .B1(n_409), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g796 ( .A1(n_253), .A2(n_322), .B1(n_502), .B2(n_694), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g938 ( .A(n_257), .Y(n_938) );
CKINVDCx20_ASAP7_75t_R g921 ( .A(n_264), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g924 ( .A(n_265), .Y(n_924) );
INVx1_ASAP7_75t_L g1014 ( .A(n_266), .Y(n_1014) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_266), .A2(n_984), .B1(n_1014), .B2(n_1018), .Y(n_1017) );
XNOR2x1_ASAP7_75t_L g867 ( .A(n_267), .B(n_868), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_268), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_269), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_270), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_271), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_272), .A2(n_313), .B1(n_535), .B2(n_572), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_273), .Y(n_906) );
AND2x2_ASAP7_75t_L g342 ( .A(n_275), .B(n_343), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_276), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_277), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_278), .Y(n_848) );
INVx1_ASAP7_75t_L g339 ( .A(n_279), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_280), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_282), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_284), .A2(n_320), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_287), .A2(n_330), .B1(n_382), .B2(n_599), .Y(n_875) );
XOR2x2_ASAP7_75t_L g837 ( .A(n_289), .B(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_293), .B(n_634), .Y(n_899) );
CKINVDCx20_ASAP7_75t_R g709 ( .A(n_297), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_298), .A2(n_328), .B1(n_450), .B2(n_534), .Y(n_897) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_299), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_301), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_302), .B(n_654), .Y(n_653) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_303), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_304), .A2(n_333), .B1(n_634), .B2(n_635), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_307), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_309), .A2(n_317), .B1(n_584), .B2(n_773), .Y(n_772) );
XNOR2x1_ASAP7_75t_L g667 ( .A(n_310), .B(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_312), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_314), .B(n_569), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_325), .B(n_375), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g988 ( .A(n_326), .Y(n_988) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_327), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_329), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_331), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_339), .Y(n_971) );
OAI21xp5_ASAP7_75t_L g1012 ( .A1(n_340), .A2(n_970), .B(n_1013), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_737), .B1(n_965), .B2(n_966), .C(n_967), .Y(n_344) );
INVx1_ASAP7_75t_L g965 ( .A(n_345), .Y(n_965) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_552), .B1(n_735), .B2(n_736), .Y(n_345) );
INVx1_ASAP7_75t_L g735 ( .A(n_346), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_432), .B1(n_550), .B2(n_551), .Y(n_346) );
INVx2_ASAP7_75t_SL g550 ( .A(n_347), .Y(n_550) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND3x1_ASAP7_75t_L g350 ( .A(n_351), .B(n_400), .C(n_418), .Y(n_350) );
NOR3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_373), .C(n_390), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_369), .B2(n_370), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_354), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_354), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_707) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_355), .Y(n_438) );
INVx2_ASAP7_75t_L g843 ( .A(n_355), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_355), .A2(n_710), .B1(n_871), .B2(n_872), .Y(n_870) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_364), .Y(n_355) );
INVx2_ASAP7_75t_L g429 ( .A(n_356), .Y(n_429) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_362), .Y(n_356) );
AND2x2_ASAP7_75t_L g372 ( .A(n_357), .B(n_362), .Y(n_372) );
AND2x2_ASAP7_75t_L g405 ( .A(n_357), .B(n_379), .Y(n_405) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g380 ( .A(n_358), .B(n_368), .Y(n_380) );
AND2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_362), .Y(n_387) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_361), .Y(n_363) );
INVx2_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
INVx1_ASAP7_75t_L g416 ( .A(n_362), .Y(n_416) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2x1p5_ASAP7_75t_L g371 ( .A(n_365), .B(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g407 ( .A(n_365), .B(n_405), .Y(n_407) );
AND2x4_ASAP7_75t_L g530 ( .A(n_365), .B(n_429), .Y(n_530) );
AND2x6_ASAP7_75t_L g569 ( .A(n_365), .B(n_372), .Y(n_569) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g378 ( .A(n_366), .Y(n_378) );
INVx1_ASAP7_75t_L g389 ( .A(n_366), .Y(n_389) );
INVx1_ASAP7_75t_L g399 ( .A(n_366), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_366), .B(n_368), .Y(n_417) );
AND2x2_ASAP7_75t_L g388 ( .A(n_367), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g412 ( .A(n_368), .B(n_399), .Y(n_412) );
OAI22xp5_ASAP7_75t_SL g437 ( .A1(n_370), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_437) );
BUFx3_ASAP7_75t_L g673 ( .A(n_370), .Y(n_673) );
INVx2_ASAP7_75t_L g846 ( .A(n_370), .Y(n_846) );
BUFx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g489 ( .A(n_371), .Y(n_489) );
AND2x2_ASAP7_75t_L g411 ( .A(n_372), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g431 ( .A(n_372), .B(n_388), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_384), .Y(n_373) );
BUFx2_ASAP7_75t_L g543 ( .A(n_375), .Y(n_543) );
INVx4_ASAP7_75t_L g564 ( .A(n_375), .Y(n_564) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_376), .Y(n_444) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_376), .Y(n_493) );
BUFx2_ASAP7_75t_L g781 ( .A(n_376), .Y(n_781) );
BUFx4f_ASAP7_75t_SL g808 ( .A(n_376), .Y(n_808) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g383 ( .A(n_378), .Y(n_383) );
INVx1_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
AND2x4_ASAP7_75t_L g382 ( .A(n_380), .B(n_383), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_380), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g532 ( .A(n_380), .B(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g545 ( .A(n_381), .Y(n_545) );
BUFx4f_ASAP7_75t_SL g782 ( .A(n_381), .Y(n_782) );
BUFx12f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_382), .Y(n_450) );
BUFx6f_ASAP7_75t_L g751 ( .A(n_382), .Y(n_751) );
INVx1_ASAP7_75t_L g810 ( .A(n_382), .Y(n_810) );
INVx3_ASAP7_75t_L g638 ( .A(n_385), .Y(n_638) );
BUFx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g446 ( .A(n_386), .Y(n_446) );
BUFx6f_ASAP7_75t_L g542 ( .A(n_386), .Y(n_542) );
INVx4_ASAP7_75t_L g560 ( .A(n_386), .Y(n_560) );
INVx2_ASAP7_75t_L g650 ( .A(n_386), .Y(n_650) );
AND2x6_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_L g396 ( .A(n_387), .Y(n_396) );
AND2x4_ASAP7_75t_L g535 ( .A(n_387), .B(n_398), .Y(n_535) );
AND2x2_ASAP7_75t_L g404 ( .A(n_388), .B(n_405), .Y(n_404) );
AND2x6_ASAP7_75t_L g428 ( .A(n_388), .B(n_429), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_394), .B2(n_395), .Y(n_390) );
BUFx3_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
INVx4_ASAP7_75t_L g497 ( .A(n_392), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_392), .A2(n_680), .B1(n_744), .B2(n_745), .Y(n_743) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_392), .Y(n_855) );
OAI22xp33_ASAP7_75t_SL g923 ( .A1(n_392), .A2(n_455), .B1(n_924), .B2(n_925), .Y(n_923) );
AND2x2_ASAP7_75t_L g665 ( .A(n_393), .B(n_424), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g456 ( .A(n_395), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_395), .A2(n_495), .B1(n_496), .B2(n_498), .Y(n_494) );
OR2x6_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_408), .Y(n_400) );
INVx3_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx3_ASAP7_75t_L g522 ( .A(n_403), .Y(n_522) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_404), .Y(n_462) );
BUFx2_ASAP7_75t_SL g509 ( .A(n_404), .Y(n_509) );
BUFx2_ASAP7_75t_SL g576 ( .A(n_404), .Y(n_576) );
AND2x2_ASAP7_75t_L g421 ( .A(n_405), .B(n_412), .Y(n_421) );
AND2x4_ASAP7_75t_L g423 ( .A(n_405), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_405), .B(n_412), .Y(n_936) );
INVx1_ASAP7_75t_L g939 ( .A(n_406), .Y(n_939) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx3_ASAP7_75t_L g479 ( .A(n_407), .Y(n_479) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_407), .Y(n_510) );
BUFx3_ASAP7_75t_L g616 ( .A(n_407), .Y(n_616) );
INVx2_ASAP7_75t_L g763 ( .A(n_407), .Y(n_763) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_409), .Y(n_720) );
BUFx2_ASAP7_75t_L g757 ( .A(n_409), .Y(n_757) );
INVx5_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx4_ASAP7_75t_L g467 ( .A(n_410), .Y(n_467) );
INVx3_ASAP7_75t_L g512 ( .A(n_410), .Y(n_512) );
INVx1_ASAP7_75t_L g608 ( .A(n_410), .Y(n_608) );
INVx2_ASAP7_75t_L g628 ( .A(n_410), .Y(n_628) );
BUFx3_ASAP7_75t_L g690 ( .A(n_410), .Y(n_690) );
INVx8_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g540 ( .A(n_414), .Y(n_540) );
BUFx2_ASAP7_75t_L g609 ( .A(n_414), .Y(n_609) );
INVx6_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g468 ( .A(n_415), .Y(n_468) );
INVx1_ASAP7_75t_SL g691 ( .A(n_415), .Y(n_691) );
INVx1_ASAP7_75t_L g721 ( .A(n_415), .Y(n_721) );
OR2x6_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g533 ( .A(n_416), .Y(n_533) );
INVx1_ASAP7_75t_L g424 ( .A(n_417), .Y(n_424) );
AND2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_425), .Y(n_418) );
BUFx2_ASAP7_75t_L g728 ( .A(n_420), .Y(n_728) );
BUFx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx3_ASAP7_75t_L g477 ( .A(n_421), .Y(n_477) );
BUFx3_ASAP7_75t_L g523 ( .A(n_421), .Y(n_523) );
BUFx3_ASAP7_75t_L g605 ( .A(n_421), .Y(n_605) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_SL g473 ( .A(n_423), .Y(n_473) );
BUFx3_ASAP7_75t_L g520 ( .A(n_423), .Y(n_520) );
BUFx2_ASAP7_75t_L g581 ( .A(n_423), .Y(n_581) );
BUFx3_ASAP7_75t_L g613 ( .A(n_423), .Y(n_613) );
INVx1_ASAP7_75t_L g695 ( .A(n_423), .Y(n_695) );
BUFx2_ASAP7_75t_SL g860 ( .A(n_423), .Y(n_860) );
INVx4_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g504 ( .A(n_427), .Y(n_504) );
INVx2_ASAP7_75t_SL g583 ( .A(n_427), .Y(n_583) );
INVx4_ASAP7_75t_L g760 ( .A(n_427), .Y(n_760) );
INVx11_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx11_ASAP7_75t_L g472 ( .A(n_428), .Y(n_472) );
BUFx3_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx3_ASAP7_75t_L g463 ( .A(n_431), .Y(n_463) );
INVx6_ASAP7_75t_L g506 ( .A(n_431), .Y(n_506) );
BUFx3_ASAP7_75t_L g663 ( .A(n_431), .Y(n_663) );
INVx1_ASAP7_75t_L g551 ( .A(n_432), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_480), .B1(n_481), .B2(n_549), .Y(n_432) );
INVx2_ASAP7_75t_L g549 ( .A(n_433), .Y(n_549) );
XNOR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_458), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_441), .C(n_452), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_438), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_438), .A2(n_488), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g917 ( .A(n_438), .Y(n_917) );
OAI222xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_445), .B1(n_446), .B2(n_447), .C1(n_448), .C2(n_451), .Y(n_441) );
INVx2_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g490 ( .A1(n_446), .A2(n_491), .B(n_492), .Y(n_490) );
OAI222xp33_ASAP7_75t_L g590 ( .A1(n_448), .A2(n_591), .B1(n_592), .B2(n_593), .C1(n_594), .C2(n_595), .Y(n_590) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx4f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B1(n_455), .B2(n_457), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_455), .A2(n_854), .B1(n_855), .B2(n_856), .Y(n_853) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g680 ( .A(n_456), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_469), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
BUFx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g685 ( .A(n_462), .Y(n_685) );
BUFx3_ASAP7_75t_L g724 ( .A(n_462), .Y(n_724) );
BUFx6f_ASAP7_75t_L g1003 ( .A(n_462), .Y(n_1003) );
INVx1_ASAP7_75t_L g727 ( .A(n_463), .Y(n_727) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g578 ( .A(n_467), .Y(n_578) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_467), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_474), .Y(n_469) );
INVx1_ASAP7_75t_L g799 ( .A(n_471), .Y(n_799) );
INVx5_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g519 ( .A(n_472), .Y(n_519) );
INVx1_ASAP7_75t_L g612 ( .A(n_472), .Y(n_612) );
INVx4_ASAP7_75t_L g773 ( .A(n_472), .Y(n_773) );
INVx2_ASAP7_75t_SL g904 ( .A(n_472), .Y(n_904) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx4f_ASAP7_75t_SL g502 ( .A(n_477), .Y(n_502) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AO22x1_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_515), .B1(n_547), .B2(n_548), .Y(n_481) );
INVx1_ASAP7_75t_L g547 ( .A(n_482), .Y(n_547) );
INVx2_ASAP7_75t_L g513 ( .A(n_483), .Y(n_513) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_499), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_490), .C(n_494), .Y(n_484) );
OA211x2_ASAP7_75t_L g524 ( .A1(n_488), .A2(n_525), .B(n_526), .C(n_531), .Y(n_524) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g710 ( .A(n_489), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_493), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_496), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_496), .A2(n_680), .B1(n_712), .B2(n_713), .Y(n_711) );
INVx3_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g880 ( .A(n_497), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_500), .B(n_507), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_503), .Y(n_500) );
INVx2_ASAP7_75t_L g932 ( .A(n_505), .Y(n_932) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g538 ( .A(n_506), .Y(n_538) );
INVx2_ASAP7_75t_L g584 ( .A(n_506), .Y(n_584) );
INVx2_ASAP7_75t_L g887 ( .A(n_506), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx4_ASAP7_75t_L g687 ( .A(n_510), .Y(n_687) );
INVx1_ASAP7_75t_L g548 ( .A(n_515), .Y(n_548) );
XOR2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_546), .Y(n_515) );
NAND4xp75_ASAP7_75t_L g516 ( .A(n_517), .B(n_524), .C(n_536), .D(n_541), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx5_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g634 ( .A(n_529), .Y(n_634) );
INVx2_ASAP7_75t_L g654 ( .A(n_529), .Y(n_654) );
INVx2_ASAP7_75t_L g815 ( .A(n_529), .Y(n_815) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx3_ASAP7_75t_L g572 ( .A(n_532), .Y(n_572) );
BUFx2_ASAP7_75t_L g598 ( .A(n_532), .Y(n_598) );
INVx1_ASAP7_75t_L g779 ( .A(n_532), .Y(n_779) );
BUFx2_ASAP7_75t_L g953 ( .A(n_532), .Y(n_953) );
INVx1_ASAP7_75t_SL g996 ( .A(n_534), .Y(n_996) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_SL g573 ( .A(n_535), .Y(n_573) );
BUFx3_ASAP7_75t_L g599 ( .A(n_535), .Y(n_599) );
BUFx2_ASAP7_75t_SL g948 ( .A(n_535), .Y(n_948) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
INVx2_ASAP7_75t_SL g805 ( .A(n_542), .Y(n_805) );
INVx2_ASAP7_75t_L g987 ( .A(n_542), .Y(n_987) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g736 ( .A(n_552), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_619), .B1(n_620), .B2(n_734), .Y(n_552) );
INVx1_ASAP7_75t_L g734 ( .A(n_553), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_586), .B2(n_618), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
XOR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_585), .Y(n_556) );
NAND3x1_ASAP7_75t_L g557 ( .A(n_558), .B(n_574), .C(n_579), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_559), .B(n_565), .Y(n_558) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_561), .B(n_562), .Y(n_559) );
BUFx2_ASAP7_75t_L g591 ( .A(n_560), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_560), .A2(n_824), .B(n_825), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g895 ( .A1(n_560), .A2(n_896), .B(n_897), .Y(n_895) );
OAI21xp5_ASAP7_75t_SL g945 ( .A1(n_560), .A2(n_946), .B(n_947), .Y(n_945) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g565 ( .A(n_566), .B(n_570), .C(n_571), .Y(n_565) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_SL g776 ( .A(n_568), .Y(n_776) );
INVx1_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
BUFx4f_ASAP7_75t_L g635 ( .A(n_569), .Y(n_635) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
INVx1_ASAP7_75t_L g618 ( .A(n_586), .Y(n_618) );
INVx1_ASAP7_75t_L g617 ( .A(n_588), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_602), .C(n_610), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_596), .Y(n_589) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_593), .A2(n_650), .B1(n_704), .B2(n_705), .C(n_706), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_606), .Y(n_602) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx2_ASAP7_75t_L g718 ( .A(n_613), .Y(n_718) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI22xp5_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_697), .B1(n_698), .B2(n_733), .Y(n_620) );
INVx1_ASAP7_75t_L g733 ( .A(n_621), .Y(n_733) );
AO22x1_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_641), .B2(n_642), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
NOR4xp75_ASAP7_75t_L g624 ( .A(n_625), .B(n_629), .C(n_632), .D(n_637), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_633), .B(n_636), .Y(n_632) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_639), .B(n_640), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g873 ( .A1(n_638), .A2(n_874), .B(n_875), .Y(n_873) );
OAI21xp33_ASAP7_75t_SL g920 ( .A1(n_638), .A2(n_921), .B(n_922), .Y(n_920) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
XNOR2x1_ASAP7_75t_SL g642 ( .A(n_643), .B(n_667), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_643), .A2(n_700), .B1(n_731), .B2(n_732), .Y(n_699) );
INVx1_ASAP7_75t_L g731 ( .A(n_643), .Y(n_731) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
XOR2x2_ASAP7_75t_L g645 ( .A(n_646), .B(n_666), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_647), .B(n_657), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_652), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B(n_651), .Y(n_648) );
OAI21xp33_ASAP7_75t_SL g674 ( .A1(n_650), .A2(n_675), .B(n_676), .Y(n_674) );
OAI21xp33_ASAP7_75t_L g746 ( .A1(n_650), .A2(n_747), .B(n_748), .Y(n_746) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_650), .A2(n_848), .B1(n_849), .B2(n_851), .C(n_852), .Y(n_847) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .C(n_656), .Y(n_652) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_681), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .C(n_677), .Y(n_669) );
OAI22xp5_ASAP7_75t_SL g915 ( .A1(n_673), .A2(n_916), .B1(n_918), .B2(n_919), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_692), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_688), .Y(n_682) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx4_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx3_ASAP7_75t_L g999 ( .A(n_687), .Y(n_999) );
INVx3_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_695), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_937) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g732 ( .A(n_700), .Y(n_732) );
INVx2_ASAP7_75t_SL g730 ( .A(n_701), .Y(n_730) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_714), .Y(n_701) );
NOR3xp33_ASAP7_75t_SL g702 ( .A(n_703), .B(n_707), .C(n_711), .Y(n_702) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_722), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g966 ( .A(n_737), .Y(n_966) );
XOR2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_785), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_765), .B1(n_783), .B2(n_784), .Y(n_738) );
INVx1_ASAP7_75t_L g783 ( .A(n_739), .Y(n_783) );
INVx2_ASAP7_75t_L g764 ( .A(n_741), .Y(n_764) );
NAND2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_755), .Y(n_741) );
NOR3xp33_ASAP7_75t_SL g742 ( .A(n_743), .B(n_746), .C(n_752), .Y(n_742) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
BUFx3_ASAP7_75t_L g850 ( .A(n_751), .Y(n_850) );
AND4x1_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .C(n_759), .D(n_761), .Y(n_755) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g784 ( .A(n_765), .Y(n_784) );
NAND4xp75_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .C(n_774), .D(n_780), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
AND2x2_ASAP7_75t_SL g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g994 ( .A(n_779), .Y(n_994) );
INVx1_ASAP7_75t_L g878 ( .A(n_781), .Y(n_878) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_788), .B1(n_835), .B2(n_964), .Y(n_786) );
INVx1_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B1(n_817), .B2(n_834), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g816 ( .A(n_793), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_794), .B(n_803), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_800), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx2_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_804), .B(n_812), .Y(n_803) );
OAI222xp33_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_807), .B2(n_809), .C1(n_810), .C2(n_811), .Y(n_804) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
INVx3_ASAP7_75t_L g834 ( .A(n_817), .Y(n_834) );
OAI22x1_ASAP7_75t_L g941 ( .A1(n_817), .A2(n_834), .B1(n_942), .B2(n_961), .Y(n_941) );
XOR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_833), .Y(n_817) );
NAND3x1_ASAP7_75t_SL g818 ( .A(n_819), .B(n_822), .C(n_830), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_823), .B(n_826), .Y(n_822) );
NAND3xp33_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .C(n_829), .Y(n_826) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
INVx1_ASAP7_75t_L g964 ( .A(n_835), .Y(n_964) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_909), .B1(n_962), .B2(n_963), .Y(n_835) );
INVx2_ASAP7_75t_L g962 ( .A(n_836), .Y(n_962) );
OA22x2_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_866), .B1(n_907), .B2(n_908), .Y(n_836) );
INVx2_ASAP7_75t_L g907 ( .A(n_837), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_857), .Y(n_838) );
NOR3xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_847), .C(n_853), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_841), .A2(n_842), .B1(n_844), .B2(n_845), .Y(n_840) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_863), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_861), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_865), .Y(n_863) );
INVx2_ASAP7_75t_L g908 ( .A(n_866), .Y(n_908) );
XOR2x2_ASAP7_75t_L g866 ( .A(n_867), .B(n_889), .Y(n_866) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_881), .Y(n_868) );
NOR3xp33_ASAP7_75t_L g869 ( .A(n_870), .B(n_873), .C(n_876), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_885), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_884), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_888), .Y(n_885) );
XOR2x2_ASAP7_75t_L g889 ( .A(n_890), .B(n_906), .Y(n_889) );
NAND3x1_ASAP7_75t_L g890 ( .A(n_891), .B(n_894), .C(n_902), .Y(n_890) );
AND2x2_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
NOR2x1_ASAP7_75t_L g894 ( .A(n_895), .B(n_898), .Y(n_894) );
NAND3xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_900), .C(n_901), .Y(n_898) );
AND2x2_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx1_ASAP7_75t_L g963 ( .A(n_909), .Y(n_963) );
XNOR2x2_ASAP7_75t_L g909 ( .A(n_910), .B(n_941), .Y(n_909) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_914), .B(n_926), .Y(n_913) );
NOR3xp33_ASAP7_75t_L g914 ( .A(n_915), .B(n_920), .C(n_923), .Y(n_914) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g926 ( .A(n_927), .B(n_930), .C(n_937), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_932), .B1(n_933), .B2(n_934), .Y(n_930) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx2_ASAP7_75t_L g961 ( .A(n_942), .Y(n_961) );
AND2x4_ASAP7_75t_L g943 ( .A(n_944), .B(n_954), .Y(n_943) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_945), .B(n_949), .Y(n_944) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .C(n_952), .Y(n_949) );
NOR2x1_ASAP7_75t_L g954 ( .A(n_955), .B(n_958), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
INVx1_ASAP7_75t_SL g967 ( .A(n_968), .Y(n_967) );
NOR2x1_ASAP7_75t_L g968 ( .A(n_969), .B(n_973), .Y(n_968) );
OR2x2_ASAP7_75t_SL g1021 ( .A(n_969), .B(n_974), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_972), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g1006 ( .A(n_970), .Y(n_1006) );
INVx1_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_971), .B(n_1010), .Y(n_1013) );
CKINVDCx16_ASAP7_75t_R g1010 ( .A(n_972), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g973 ( .A(n_974), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_979), .Y(n_977) );
OAI322xp33_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_1005), .A3(n_1007), .B1(n_1011), .B2(n_1014), .C1(n_1015), .C2(n_1019), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g982 ( .A(n_983), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g1018 ( .A(n_984), .Y(n_1018) );
NAND3x1_ASAP7_75t_L g984 ( .A(n_985), .B(n_997), .C(n_1001), .Y(n_984) );
NOR2x1_ASAP7_75t_L g985 ( .A(n_986), .B(n_990), .Y(n_985) );
OAI21xp5_ASAP7_75t_SL g986 ( .A1(n_987), .A2(n_988), .B(n_989), .Y(n_986) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_991), .B(n_992), .C(n_993), .Y(n_990) );
INVx2_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
AND2x2_ASAP7_75t_L g997 ( .A(n_998), .B(n_1000), .Y(n_997) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1004), .Y(n_1001) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
BUFx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
CKINVDCx16_ASAP7_75t_R g1011 ( .A(n_1012), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_1020), .Y(n_1019) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_1021), .Y(n_1020) );
endmodule