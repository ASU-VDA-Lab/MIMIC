module fake_netlist_1_6738_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
BUFx8_ASAP7_75t_SL g3 ( .A(n_2), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_0), .B(n_2), .Y(n_4) );
NAND2x1p5_ASAP7_75t_L g5 ( .A(n_4), .B(n_0), .Y(n_5) );
OAI22xp5_ASAP7_75t_SL g6 ( .A1(n_3), .A2(n_2), .B1(n_1), .B2(n_0), .Y(n_6) );
NAND2x1_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
INVx1_ASAP7_75t_SL g8 ( .A(n_5), .Y(n_8) );
INVxp67_ASAP7_75t_SL g9 ( .A(n_8), .Y(n_9) );
AOI221xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_6), .B1(n_7), .B2(n_4), .C(n_3), .Y(n_10) );
OAI22xp33_ASAP7_75t_SL g11 ( .A1(n_9), .A2(n_0), .B1(n_1), .B2(n_8), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
AOI22xp33_ASAP7_75t_SL g13 ( .A1(n_12), .A2(n_1), .B1(n_10), .B2(n_9), .Y(n_13) );
endmodule