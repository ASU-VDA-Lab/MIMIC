module real_jpeg_33704_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_0),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_0),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_0),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_0),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_1),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_2),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_3),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_4),
.Y(n_88)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_4),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_192),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_5),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_5),
.A2(n_195),
.B1(n_282),
.B2(n_287),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_5),
.A2(n_195),
.B1(n_339),
.B2(n_343),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_5),
.A2(n_195),
.B1(n_361),
.B2(n_367),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_6),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_6),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_6),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_8),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_147),
.B1(n_159),
.B2(n_162),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g437 ( 
.A1(n_8),
.A2(n_105),
.B1(n_147),
.B2(n_438),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_8),
.A2(n_147),
.B1(n_511),
.B2(n_513),
.Y(n_510)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

OAI22x1_ASAP7_75t_SL g62 ( 
.A1(n_10),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_10),
.Y(n_66)
);

AO22x2_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_66),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_10),
.A2(n_66),
.B1(n_208),
.B2(n_211),
.Y(n_207)
);

OAI22x1_ASAP7_75t_L g240 ( 
.A1(n_10),
.A2(n_66),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_11),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_11),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_12),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_12),
.A2(n_51),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AO22x1_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_51),
.B1(n_220),
.B2(n_223),
.Y(n_219)
);

AOI22x1_ASAP7_75t_SL g259 ( 
.A1(n_12),
.A2(n_51),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_SL g452 ( 
.A(n_12),
.B(n_453),
.Y(n_452)
);

OAI32xp33_ASAP7_75t_L g477 ( 
.A1(n_12),
.A2(n_478),
.A3(n_484),
.B1(n_486),
.B2(n_490),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_12),
.B(n_154),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_15),
.B(n_18),
.Y(n_14)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_SL g16 ( 
.A(n_17),
.Y(n_16)
);

AOI21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_70),
.B(n_550),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_54),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_20),
.A2(n_313),
.B(n_351),
.Y(n_404)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_21),
.A2(n_395),
.B(n_425),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_22),
.A2(n_314),
.B1(n_317),
.B2(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_22),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_45),
.B(n_46),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_23),
.B(n_46),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_23),
.B(n_158),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_23),
.Y(n_370)
);

NOR2x1p5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_35),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_26),
.Y(n_164)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_29),
.Y(n_182)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_32),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_32),
.Y(n_177)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_35),
.B(n_158),
.Y(n_157)
);

AO22x2_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_38),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g342 ( 
.A(n_38),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_41),
.Y(n_184)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_57),
.Y(n_56)
);

OAI21x1_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_51),
.B(n_52),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_50),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_51),
.B(n_58),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g442 ( 
.A1(n_51),
.A2(n_443),
.A3(n_446),
.B1(n_451),
.B2(n_452),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_51),
.B(n_487),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_51),
.B(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_51),
.B(n_201),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_52),
.Y(n_185)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_54),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_56),
.B(n_255),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_57),
.B(n_62),
.Y(n_254)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_58),
.Y(n_375)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OA21x2_ASAP7_75t_SL g374 ( 
.A1(n_60),
.A2(n_360),
.B(n_375),
.Y(n_374)
);

OA21x2_ASAP7_75t_SL g383 ( 
.A1(n_60),
.A2(n_360),
.B(n_375),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_61),
.B(n_157),
.Y(n_298)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_419),
.C(n_426),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_356),
.C(n_397),
.Y(n_71)
);

INVxp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_325),
.B(n_327),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_300),
.B(n_303),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_266),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_232),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_77),
.B(n_232),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_165),
.C(n_213),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_78),
.B(n_456),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_155),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_109),
.Y(n_79)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_80),
.B(n_109),
.C(n_155),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_80),
.B(n_374),
.C(n_376),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_80),
.A2(n_377),
.B(n_385),
.Y(n_384)
);

NOR3xp33_ASAP7_75t_L g385 ( 
.A(n_80),
.B(n_345),
.C(n_379),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_80),
.Y(n_392)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_80),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_92),
.B(n_102),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_81),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_81),
.B(n_281),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g316 ( 
.A1(n_81),
.A2(n_92),
.B1(n_240),
.B2(n_281),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_81),
.B(n_102),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_81),
.B(n_437),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_81),
.Y(n_526)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_93),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_91),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_85),
.Y(n_498)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_87),
.Y(n_198)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_87),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_87),
.Y(n_489)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_88),
.Y(n_206)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_92),
.B(n_102),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_92),
.B(n_240),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_92),
.B(n_437),
.Y(n_436)
);

OAI22xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_96),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_96),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_101),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_104),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_107),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_108),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_145),
.Y(n_109)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_110),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_111),
.B(n_154),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_L g391 ( 
.A(n_111),
.B(n_154),
.Y(n_391)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_119),
.B(n_146),
.Y(n_228)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_120),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g323 ( 
.A(n_120),
.B(n_259),
.Y(n_323)
);

AO21x2_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_129),
.B(n_137),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g451 ( 
.A(n_121),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_133),
.A2(n_138),
.B1(n_140),
.B2(n_142),
.Y(n_137)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_138),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_145),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_154),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_154),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_154),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_154),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_156),
.B(n_254),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_165),
.B(n_214),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_186),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_166),
.B(n_186),
.Y(n_250)
);

OAI31xp33_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_170),
.A3(n_174),
.B(n_178),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_183),
.B(n_185),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_183),
.Y(n_343)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_191),
.B(n_199),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_207),
.Y(n_226)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_191),
.A2(n_226),
.B(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_193),
.Y(n_512)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_199),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_199),
.B(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_200),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_200),
.B(n_510),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_227),
.B(n_231),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_215),
.A2(n_216),
.B(n_217),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_217),
.Y(n_231)
);

NOR2x1p5_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_225),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_218),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_219),
.Y(n_315)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_222),
.Y(n_224)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g527 ( 
.A(n_226),
.B(n_509),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_227),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

NOR2x1p5_ASAP7_75t_SL g322 ( 
.A(n_230),
.B(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_248),
.Y(n_232)
);

XOR2x1_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_247),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_247),
.C(n_248),
.Y(n_267)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_235),
.B(n_237),
.Y(n_299)
);

AO21x2_ASAP7_75t_L g314 ( 
.A1(n_236),
.A2(n_277),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_238),
.B(n_471),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_239),
.B(n_436),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_246),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_265),
.C(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_265),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_254),
.A2(n_360),
.B(n_370),
.Y(n_359)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_257),
.Y(n_379)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_259),
.A2(n_296),
.B(n_297),
.Y(n_295)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_266),
.B(n_548),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_267),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_268),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_292),
.B2(n_293),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_273),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_271),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_274),
.A2(n_280),
.B(n_291),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_275),
.B(n_509),
.Y(n_508)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_291),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_291),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_305),
.C(n_307),
.Y(n_304)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_299),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_297),
.A2(n_338),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_299),
.C(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR3xp33_ASAP7_75t_L g546 ( 
.A(n_303),
.B(n_328),
.C(n_547),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_304),
.B(n_308),
.Y(n_326)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_310),
.A2(n_359),
.B1(n_371),
.B2(n_372),
.Y(n_358)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_319),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_330),
.C(n_331),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_SL g441 ( 
.A(n_314),
.B(n_442),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_314),
.A2(n_317),
.B1(n_442),
.B2(n_465),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_317),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_319),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_320),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_323),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_324),
.Y(n_353)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_329),
.B(n_332),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_352),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_348),
.Y(n_333)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_346),
.Y(n_334)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_335),
.B(n_346),
.Y(n_412)
);

NAND2x1_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_344),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_347),
.B(n_436),
.Y(n_435)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_348),
.Y(n_400)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_351),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_352),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.C(n_355),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_356),
.A2(n_420),
.B(n_423),
.Y(n_419)
);

NAND3xp33_ASAP7_75t_L g426 ( 
.A(n_356),
.B(n_397),
.C(n_427),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_380),
.B(n_394),
.Y(n_356)
);

OAI31xp33_ASAP7_75t_SL g423 ( 
.A1(n_357),
.A2(n_380),
.A3(n_394),
.B(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_373),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_359),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_371),
.C(n_373),
.Y(n_396)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx6_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.C(n_387),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_386),
.B1(n_393),
.B2(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_382),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_386),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_386),
.A2(n_393),
.B1(n_408),
.B2(n_410),
.Y(n_407)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.C(n_393),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_396),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_413),
.Y(n_397)
);

NOR2xp67_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.C(n_402),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_404),
.B(n_411),
.C(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_406),
.A2(n_407),
.B1(n_411),
.B2(n_412),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_408),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_413),
.A2(n_421),
.B(n_422),
.Y(n_420)
);

NOR2x1_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_414),
.B(n_416),
.Y(n_422)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_546),
.B(n_549),
.Y(n_428)
);

AO21x1_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_457),
.B(n_545),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_455),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_431),
.B(n_455),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.C(n_441),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_433),
.B1(n_460),
.B2(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_435),
.B(n_441),
.Y(n_461)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx8_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_SL g453 ( 
.A(n_454),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_472),
.B(n_544),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_459),
.B(n_462),
.Y(n_544)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_466),
.C(n_469),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g463 ( 
.A(n_464),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_464),
.B(n_540),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_466),
.A2(n_467),
.B1(n_469),
.B2(n_470),
.Y(n_540)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_538),
.B(n_543),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_516),
.B(n_537),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_501),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_475),
.B(n_501),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_499),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_476),
.A2(n_477),
.B1(n_499),
.B2(n_500),
.Y(n_522)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_483),
.Y(n_515)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_494),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_507),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_508),
.C(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_510),
.B(n_520),
.Y(n_519)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_513),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_523),
.B(n_536),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_522),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_522),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_530),
.Y(n_529)
);

BUFx4f_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_524),
.A2(n_528),
.B(n_535),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_527),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_525),
.B(n_527),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_534),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_541),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_539),
.B(n_541),
.Y(n_543)
);


endmodule