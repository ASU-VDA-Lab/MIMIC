module fake_jpeg_26457_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_30),
.B(n_32),
.Y(n_59)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_30),
.B(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_44),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_24),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_48),
.B(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_19),
.B1(n_25),
.B2(n_23),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_14),
.B1(n_39),
.B2(n_29),
.Y(n_78)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_24),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_26),
.C(n_23),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_19),
.B1(n_25),
.B2(n_15),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_39),
.B1(n_29),
.B2(n_27),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_37),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_20),
.C(n_15),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_73),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_72),
.B1(n_43),
.B2(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_20),
.B1(n_14),
.B2(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_78),
.B1(n_43),
.B2(n_52),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_44),
.C(n_57),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_83),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_60),
.B1(n_61),
.B2(n_75),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_91),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_48),
.B(n_41),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_48),
.C(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_64),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_58),
.C(n_59),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_80),
.A2(n_78),
.B1(n_68),
.B2(n_43),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_101),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_79),
.C(n_87),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_111),
.C(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_89),
.C(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_114),
.B1(n_67),
.B2(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_106),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_99),
.B1(n_98),
.B2(n_96),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_109),
.A2(n_96),
.B1(n_81),
.B2(n_84),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_42),
.B1(n_97),
.B2(n_65),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_125),
.B1(n_120),
.B2(n_117),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_65),
.B1(n_69),
.B2(n_27),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_126),
.B(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_116),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_115),
.C(n_118),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_7),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_4),
.B(n_5),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_129),
.B(n_6),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_136),
.Y(n_137)
);


endmodule