module real_jpeg_5256_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g128 ( 
.A(n_0),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_1),
.A2(n_64),
.B1(n_182),
.B2(n_186),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_3),
.A2(n_83),
.B1(n_139),
.B2(n_216),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_3),
.A2(n_83),
.B1(n_293),
.B2(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_3),
.A2(n_70),
.B1(n_83),
.B2(n_311),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_4),
.A2(n_156),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_4),
.A2(n_177),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_4),
.A2(n_56),
.B1(n_177),
.B2(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_5),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_5),
.Y(n_251)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_7),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_7),
.Y(n_249)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_8),
.A2(n_73),
.B1(n_241),
.B2(n_244),
.Y(n_240)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_9),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_11),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_12),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_12),
.A2(n_100),
.B1(n_101),
.B2(n_137),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_12),
.A2(n_137),
.B1(n_274),
.B2(n_311),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_12),
.A2(n_137),
.B1(n_293),
.B2(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_13),
.Y(n_164)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_13),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_14),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_15),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_99),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_15),
.A2(n_99),
.B1(n_203),
.B2(n_206),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_15),
.A2(n_56),
.B1(n_70),
.B2(n_99),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_16),
.A2(n_40),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_16),
.B(n_302),
.C(n_305),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_16),
.B(n_125),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_16),
.B(n_249),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_16),
.B(n_179),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_16),
.B(n_360),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_259),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_258),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_220),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_21),
.B(n_220),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_150),
.C(n_199),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_22),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_23),
.B(n_77),
.C(n_111),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_24),
.A2(n_44),
.B1(n_45),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_24),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.A3(n_30),
.B1(n_34),
.B2(n_39),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_26),
.Y(n_145)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_27),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_27),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_28),
.A2(n_31),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_36),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_114)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_37),
.A2(n_40),
.B(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_38),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g210 ( 
.A1(n_39),
.A2(n_40),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_40),
.B(n_89),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_40),
.A2(n_46),
.B(n_312),
.Y(n_331)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_53),
.B1(n_65),
.B2(n_68),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_46),
.A2(n_191),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_46),
.A2(n_310),
.B(n_312),
.Y(n_309)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_47),
.A2(n_69),
.B1(n_190),
.B2(n_197),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_47),
.A2(n_54),
.B1(n_273),
.B2(n_278),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_47),
.B(n_314),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_47),
.A2(n_66),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_52),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_57),
.Y(n_307)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_58),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_63),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_65),
.A2(n_336),
.B(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_72),
.Y(n_254)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_110),
.B2(n_111),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_87),
.B(n_97),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_79),
.A2(n_89),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_88),
.B(n_98),
.Y(n_213)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_89)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g367 ( 
.A(n_94),
.Y(n_367)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_105),
.Y(n_97)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_105),
.A2(n_210),
.B(n_212),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_105),
.Y(n_234)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_133),
.B(n_141),
.Y(n_111)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_112),
.A2(n_125),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_112),
.B(n_227),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_112),
.A2(n_141),
.B(n_357),
.Y(n_356)
);

INVx3_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_113),
.A2(n_134),
.B1(n_149),
.B2(n_215),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_125),
.Y(n_113)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_125),
.Y(n_149)
);

AO22x2_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_129),
.B2(n_131),
.Y(n_125)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_128),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_128),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_130),
.Y(n_297)
);

AOI32xp33_ASAP7_75t_L g366 ( 
.A1(n_131),
.A2(n_293),
.A3(n_359),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_132),
.Y(n_369)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_149),
.Y(n_141)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_142),
.Y(n_227)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_149),
.A2(n_215),
.B(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_150),
.A2(n_151),
.B1(n_199),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_189),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_152),
.B(n_189),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_175),
.B1(n_178),
.B2(n_180),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_153),
.A2(n_292),
.B(n_298),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_153),
.A2(n_178),
.B1(n_318),
.B2(n_353),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_153),
.A2(n_298),
.B(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_154),
.A2(n_179),
.B1(n_181),
.B2(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_167),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_165),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_167),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_167),
.A2(n_201),
.B(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_169),
.Y(n_304)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_172),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_175),
.A2(n_178),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_179),
.B(n_202),
.Y(n_298)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_199),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_208),
.C(n_214),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_200),
.B(n_214),
.Y(n_264)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_204),
.Y(n_354)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_206),
.Y(n_245)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_208),
.A2(n_209),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_219),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_238),
.B1(n_256),
.B2(n_257),
.Y(n_222)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_246),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_244),
.Y(n_319)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_249),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_285),
.B(n_388),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_282),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_262),
.B(n_282),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.C(n_269),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_263),
.B(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_269),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.C(n_281),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_270),
.B(n_379),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_272),
.B(n_281),
.Y(n_379)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_273),
.Y(n_365)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_382),
.B(n_387),
.Y(n_285)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_371),
.B(n_381),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_347),
.B(n_370),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_322),
.B(n_346),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_308),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_290),
.B(n_308),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_299),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_291),
.A2(n_299),
.B1(n_300),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_315),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_316),
.C(n_321),
.Y(n_348)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_310),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_313),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_320),
.B2(n_321),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_319),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_339),
.B(n_345),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_332),
.B(n_338),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_331),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_337),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_337),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_335),
.B(n_336),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_334),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_343),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_349),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_363),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_355),
.B2(n_356),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_355),
.C(n_363),
.Y(n_372)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_366),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_372),
.B(n_373),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_378),
.B2(n_380),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_377),
.C(n_380),
.Y(n_383)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_378),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_383),
.B(n_384),
.Y(n_387)
);


endmodule