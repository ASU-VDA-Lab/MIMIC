module real_jpeg_16663_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_L g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

AND2x4_ASAP7_75t_SL g68 ( 
.A(n_0),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_0),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_0),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_0),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_0),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_1),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_1),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_1),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_1),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_1),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_2),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_3),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_3),
.Y(n_327)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_3),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_4),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_4),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_4),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_4),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_4),
.B(n_422),
.Y(n_421)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_5),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_6),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_7),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_7),
.Y(n_146)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_7),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_7),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_8),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_8),
.B(n_168),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_8),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_8),
.B(n_193),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_8),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_8),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_9),
.A2(n_15),
.B1(n_36),
.B2(n_39),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_9),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_9),
.B(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_9),
.B(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_10),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_10),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_10),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_11),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_11),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_11),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_11),
.B(n_50),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_11),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_11),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_11),
.B(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_12),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_13),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_13),
.B(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_13),
.B(n_433),
.Y(n_432)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

BUFx4f_ASAP7_75t_L g362 ( 
.A(n_14),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_15),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_15),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_15),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_15),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_15),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_15),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_15),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_15),
.B(n_339),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_16),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_394),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_213),
.B(n_393),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_171),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_20),
.B(n_171),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_92),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_21),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_57),
.C(n_78),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_23),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.C(n_43),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_24),
.B(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_25),
.B(n_28),
.C(n_32),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_25),
.B(n_163),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_30),
.B(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_31),
.Y(n_190)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_31),
.Y(n_309)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_33),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_34),
.A2(n_35),
.B1(n_43),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_35),
.A2(n_236),
.B(n_242),
.Y(n_235)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_42),
.Y(n_165)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_42),
.Y(n_267)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_43),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.C(n_55),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_44),
.A2(n_45),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_44),
.A2(n_45),
.B1(n_55),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g439 ( 
.A(n_45),
.B(n_103),
.C(n_119),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_49),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_54),
.Y(n_142)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_55),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_58),
.A2(n_79),
.B1(n_80),
.B2(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_58),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.C(n_72),
.Y(n_58)
);

XOR2x2_ASAP7_75t_SL g207 ( 
.A(n_59),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.C(n_65),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_60),
.A2(n_65),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_60),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_60),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_62),
.B(n_249),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_64),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_65),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_69),
.Y(n_353)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_76),
.Y(n_241)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_81),
.B(n_89),
.C(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_88),
.B2(n_89),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_84),
.B(n_221),
.C(n_231),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_84),
.A2(n_231),
.B1(n_232),
.B2(n_379),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_84),
.Y(n_379)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_91),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_123),
.B1(n_169),
.B2(n_170),
.Y(n_92)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_93),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_93),
.B(n_398),
.C(n_399),
.Y(n_397)
);

XOR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_116),
.Y(n_93)
);

XNOR2x1_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_95),
.B(n_104),
.C(n_116),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_103),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_103),
.B1(n_121),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_103),
.Y(n_121)
);

XNOR2x2_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_105),
.B(n_112),
.C(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_107),
.Y(n_419)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_111),
.Y(n_155)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_114),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_115),
.Y(n_263)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_119),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g410 ( 
.A1(n_119),
.A2(n_122),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_120),
.B(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_156),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_124),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_143),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_128),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_134),
.C(n_139),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_129),
.A2(n_139),
.B1(n_140),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_132),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_134),
.B(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_139),
.B(n_260),
.C(n_264),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_139),
.A2(n_140),
.B1(n_264),
.B2(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2x2_ASAP7_75t_SL g176 ( 
.A(n_143),
.B(n_177),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_148),
.C(n_153),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_157),
.B(n_159),
.C(n_402),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_160),
.B(n_162),
.C(n_167),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_169),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_176),
.Y(n_285)
);

INVxp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_179),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_207),
.C(n_210),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_180),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.C(n_194),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2x2_ASAP7_75t_L g270 ( 
.A(n_182),
.B(n_271),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_186),
.B(n_194),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_192),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_187),
.B(n_192),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.C(n_202),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_195),
.A2(n_200),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_200),
.A2(n_257),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_200),
.B(n_344),
.C(n_347),
.Y(n_369)
);

XOR2x1_ASAP7_75t_L g254 ( 
.A(n_202),
.B(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_207),
.B(n_210),
.Y(n_279)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_286),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_280),
.C(n_282),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_272),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_218),
.B(n_272),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_252),
.C(n_270),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_219),
.B(n_389),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_234),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_220),
.B(n_235),
.C(n_248),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_221),
.B(n_378),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_226),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_222),
.B(n_226),
.Y(n_320)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_222),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_222),
.A2(n_337),
.B1(n_338),
.B2(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_229),
.Y(n_247)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_229),
.Y(n_340)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_248),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_250),
.B(n_295),
.C(n_296),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_253),
.B(n_270),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_258),
.C(n_268),
.Y(n_253)
);

XOR2x1_ASAP7_75t_L g383 ( 
.A(n_254),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_259),
.B(n_269),
.Y(n_384)
);

XOR2x1_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_265),
.Y(n_409)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_275),
.C(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_281),
.B(n_283),
.Y(n_392)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND3xp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.C(n_392),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_387),
.B(n_391),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_372),
.B(n_386),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_333),
.B(n_371),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_316),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_292),
.B(n_316),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.C(n_306),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_293),
.B(n_367),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_299),
.B1(n_306),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_305),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_300),
.B(n_305),
.Y(n_348)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

AO22x1_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_310),
.B1(n_314),
.B2(n_315),
.Y(n_306)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_314),
.Y(n_318)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_328),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_317),
.B(n_329),
.C(n_330),
.Y(n_385)
);

XOR2x1_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_320),
.C(n_321),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

AOI21x1_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_365),
.B(n_370),
.Y(n_333)
);

OAI21x1_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_349),
.B(n_364),
.Y(n_334)
);

NOR2x1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_341),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_338),
.Y(n_355)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_342),
.A2(n_343),
.B1(n_347),
.B2(n_348),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI21x1_ASAP7_75t_SL g349 ( 
.A1(n_350),
.A2(n_356),
.B(n_363),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_354),
.Y(n_363)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_369),
.Y(n_365)
);

NOR2x1_ASAP7_75t_SL g370 ( 
.A(n_366),
.B(n_369),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_385),
.Y(n_372)
);

NOR2x1_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_385),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_375),
.B1(n_382),
.B2(n_383),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_380),
.B2(n_381),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_381),
.C(n_382),
.Y(n_390)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_388),
.B(n_390),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_444),
.Y(n_394)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_400),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_397),
.B(n_400),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_435),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_417),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.Y(n_406)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.Y(n_420)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_432),
.Y(n_425)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_443),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_442),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_438),
.A2(n_439),
.B1(n_440),
.B2(n_441),
.Y(n_437)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_438),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_439),
.Y(n_440)
);


endmodule