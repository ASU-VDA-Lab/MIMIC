module real_jpeg_9788_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_70;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_202;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_0),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_1),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_1),
.A2(n_46),
.B1(n_56),
.B2(n_57),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_1),
.A2(n_46),
.B1(n_65),
.B2(n_71),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_22),
.B1(n_26),
.B2(n_46),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_1),
.A2(n_3),
.B(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_1),
.B(n_96),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_1),
.A2(n_6),
.B(n_22),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_51),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g186 ( 
.A1(n_1),
.A2(n_53),
.B(n_57),
.C(n_187),
.Y(n_186)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_3),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_6),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_37),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_6),
.A2(n_22),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_25),
.B1(n_37),
.B2(n_43),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_10),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_10),
.A2(n_44),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_10),
.A2(n_44),
.B1(n_65),
.B2(n_71),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_22),
.B1(n_26),
.B2(n_44),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_120),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_118),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_102),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_15),
.B(n_102),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_84),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_74),
.B2(n_75),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_47),
.B1(n_48),
.B2(n_73),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_34),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_20),
.A2(n_34),
.B1(n_35),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_20),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_26),
.B(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_27),
.B(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_28),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_28),
.A2(n_29),
.B1(n_90),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_29),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_29),
.B(n_46),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_30),
.A2(n_89),
.B(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_34),
.A2(n_35),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_34),
.A2(n_35),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_35),
.B(n_116),
.C(n_177),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_35),
.B(n_194),
.C(n_200),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_36),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_36),
.B(n_40),
.Y(n_130)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_43),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_37),
.A2(n_46),
.B(n_54),
.Y(n_187)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_40),
.B(n_46),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_41),
.A2(n_43),
.B(n_46),
.C(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_42),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_45),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_46),
.A2(n_65),
.B(n_66),
.C(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_49),
.A2(n_50),
.B1(n_128),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_49),
.A2(n_50),
.B1(n_91),
.B2(n_92),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_50),
.B(n_95),
.C(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_50),
.B(n_92),
.C(n_189),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B(n_58),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_51),
.A2(n_55),
.B1(n_101),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_53),
.B(n_57),
.C(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_57),
.Y(n_61)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_59),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_110),
.C(n_112),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_62),
.A2(n_63),
.B1(n_110),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_72),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_72),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_83),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_78),
.B(n_90),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.C(n_98),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_86),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_91),
.A2(n_92),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_92),
.B(n_161),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_105),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.C(n_108),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_106),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_109),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_148),
.C(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_110),
.A2(n_133),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_116),
.B(n_169),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_116),
.A2(n_145),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_152),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_137),
.B(n_151),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_123),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_134),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_134),
.Y(n_151)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.CI(n_131),
.CON(n_124),
.SN(n_124)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_138),
.B(n_139),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_146),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_140),
.B(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_144),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_148),
.A2(n_149),
.B1(n_165),
.B2(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_159),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_208),
.C(n_209),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_202),
.B(n_207),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_191),
.B(n_201),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_180),
.B(n_190),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_172),
.B(n_179),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_163),
.B(n_171),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_168),
.B(n_170),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_173),
.B(n_174),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_182),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_189),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_185),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_193),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);


endmodule