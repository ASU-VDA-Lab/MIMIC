module fake_jpeg_15906_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_57),
.B1(n_20),
.B2(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_53),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_19),
.B1(n_38),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_74),
.B1(n_27),
.B2(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_53),
.Y(n_66)
);

INVxp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_0),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_17),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_40),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_82),
.Y(n_96)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_76),
.B1(n_83),
.B2(n_66),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_86),
.B1(n_58),
.B2(n_17),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_38),
.B1(n_20),
.B2(n_16),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_45),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_78),
.B(n_80),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_39),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_54),
.A2(n_18),
.B1(n_32),
.B2(n_26),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_30),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_30),
.C(n_24),
.Y(n_88)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_41),
.A2(n_34),
.A3(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_26),
.A3(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_34),
.B1(n_56),
.B2(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_91),
.B1(n_94),
.B2(n_98),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_29),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_0),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_71),
.B1(n_67),
.B2(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_99),
.B(n_24),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_53),
.B1(n_31),
.B2(n_23),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_100),
.A2(n_104),
.B1(n_112),
.B2(n_62),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_65),
.B1(n_80),
.B2(n_72),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_63),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_28),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_107),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_28),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_93),
.B1(n_97),
.B2(n_89),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_0),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_68),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_100),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_90),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_128),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_92),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_123),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_1),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_139),
.B(n_2),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_96),
.B(n_64),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_89),
.B1(n_81),
.B2(n_60),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_64),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_130),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_127),
.A2(n_112),
.B1(n_89),
.B2(n_107),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_135),
.C(n_99),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_110),
.B(n_10),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_110),
.B(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_62),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_104),
.B(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_95),
.B(n_63),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_138),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_60),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_114),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_128),
.B1(n_136),
.B2(n_127),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_142),
.A2(n_146),
.B1(n_159),
.B2(n_61),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_144),
.C(n_154),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_97),
.C(n_105),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_113),
.A2(n_87),
.B1(n_108),
.B2(n_94),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_148),
.Y(n_184)
);

NOR2x1_ASAP7_75t_SL g149 ( 
.A(n_120),
.B(n_107),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_151),
.B(n_166),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_157),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_111),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_122),
.A2(n_8),
.B(n_12),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_125),
.B(n_115),
.C(n_132),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_61),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_170),
.B(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_115),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_174),
.B(n_180),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_192),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_138),
.C(n_117),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_178),
.C(n_179),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_117),
.C(n_121),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_121),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_153),
.B(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_118),
.Y(n_185)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_150),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_178),
.C(n_174),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_153),
.B(n_8),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_205),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_206),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_149),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_164),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_207),
.B(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_171),
.A2(n_167),
.B1(n_152),
.B2(n_159),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_208),
.A2(n_181),
.B1(n_189),
.B2(n_187),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_142),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_211),
.C(n_184),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_147),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_177),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_186),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_215),
.C(n_218),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_214),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_181),
.B(n_189),
.Y(n_216)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_169),
.B1(n_184),
.B2(n_164),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_169),
.B1(n_158),
.B2(n_146),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_162),
.B1(n_158),
.B2(n_180),
.Y(n_221)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_190),
.C(n_117),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_226),
.C(n_2),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_212),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_194),
.B1(n_206),
.B2(n_208),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_233),
.B1(n_227),
.B2(n_3),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_214),
.A2(n_197),
.B(n_201),
.C(n_203),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_236),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_211),
.B1(n_200),
.B2(n_209),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_196),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.C(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_2),
.C(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_239),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_221),
.CI(n_217),
.CON(n_240),
.SN(n_240)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_5),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_244),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_218),
.C(n_226),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_229),
.C(n_7),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_246),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_235),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_232),
.A2(n_4),
.B(n_5),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_237),
.C(n_6),
.Y(n_251)
);

OAI221xp5_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_231),
.B1(n_230),
.B2(n_233),
.C(n_238),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_251),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_254),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_244),
.B(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_258),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_253),
.A2(n_240),
.B(n_242),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_255),
.A2(n_252),
.B(n_257),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_255),
.A2(n_250),
.B(n_240),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_9),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_12),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_262),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_260),
.Y(n_267)
);


endmodule