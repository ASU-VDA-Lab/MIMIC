module real_aes_13904_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g111 ( .A1(n_0), .A2(n_48), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g146 ( .A(n_0), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_1), .B(n_140), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_2), .A2(n_23), .B1(n_533), .B2(n_534), .Y(n_532) );
OAI222xp33_ASAP7_75t_SL g578 ( .A1(n_2), .A2(n_42), .B1(n_76), .B2(n_579), .C1(n_583), .C2(n_588), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_3), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_4), .B(n_203), .Y(n_264) );
BUFx3_ASAP7_75t_L g566 ( .A(n_5), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_6), .B(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g485 ( .A(n_7), .Y(n_485) );
INVx2_ASAP7_75t_L g573 ( .A(n_8), .Y(n_573) );
INVx1_ASAP7_75t_L g582 ( .A(n_8), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_9), .B(n_142), .Y(n_218) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_10), .A2(n_45), .B1(n_497), .B2(n_502), .C(n_507), .Y(n_496) );
INVx1_ASAP7_75t_L g606 ( .A(n_10), .Y(n_606) );
INVx1_ASAP7_75t_L g528 ( .A(n_11), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_12), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_13), .B(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_14), .Y(n_244) );
INVx1_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
BUFx3_ASAP7_75t_L g121 ( .A(n_15), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_16), .B(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_17), .Y(n_258) );
BUFx10_ASAP7_75t_L g683 ( .A(n_18), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_19), .A2(n_42), .B1(n_544), .B2(n_547), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g635 ( .A1(n_19), .A2(n_636), .B(n_642), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_20), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g549 ( .A(n_21), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_22), .Y(n_238) );
INVx1_ASAP7_75t_L g630 ( .A(n_23), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_24), .B(n_140), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_25), .B(n_116), .Y(n_126) );
XNOR2xp5_ASAP7_75t_L g473 ( .A(n_26), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g486 ( .A(n_27), .B(n_487), .Y(n_486) );
INVxp33_ASAP7_75t_L g495 ( .A(n_27), .Y(n_495) );
AND2x2_ASAP7_75t_L g520 ( .A(n_27), .B(n_39), .Y(n_520) );
INVx1_ASAP7_75t_L g542 ( .A(n_27), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_28), .B(n_128), .Y(n_159) );
INVx1_ASAP7_75t_L g660 ( .A(n_28), .Y(n_660) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_29), .B(n_120), .Y(n_185) );
INVx1_ASAP7_75t_L g85 ( .A(n_30), .Y(n_85) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_31), .A2(n_162), .B(n_235), .C(n_237), .Y(n_234) );
INVx2_ASAP7_75t_L g482 ( .A(n_32), .Y(n_482) );
INVx1_ASAP7_75t_L g526 ( .A(n_33), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_34), .B(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_35), .B(n_93), .Y(n_217) );
INVx1_ASAP7_75t_L g508 ( .A(n_36), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_37), .B(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_38), .Y(n_513) );
INVx2_ASAP7_75t_L g487 ( .A(n_39), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_39), .B(n_542), .Y(n_541) );
AO221x1_ASAP7_75t_L g133 ( .A1(n_40), .A2(n_64), .B1(n_116), .B2(n_123), .C(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g692 ( .A(n_40), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_41), .B(n_158), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_43), .Y(n_669) );
AND2x4_ASAP7_75t_L g84 ( .A(n_44), .B(n_85), .Y(n_84) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_44), .Y(n_655) );
INVx1_ASAP7_75t_L g622 ( .A(n_45), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g164 ( .A(n_46), .B(n_162), .C(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g571 ( .A(n_47), .Y(n_571) );
INVx1_ASAP7_75t_L g587 ( .A(n_47), .Y(n_587) );
INVx1_ASAP7_75t_L g147 ( .A(n_48), .Y(n_147) );
INVx1_ASAP7_75t_L g112 ( .A(n_49), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g209 ( .A1(n_50), .A2(n_210), .B(n_212), .C(n_214), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_51), .Y(n_242) );
INVx2_ASAP7_75t_L g213 ( .A(n_52), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_53), .B(n_110), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_54), .B(n_197), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_55), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_55), .Y(n_670) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_56), .Y(n_662) );
AND2x2_ASAP7_75t_L g206 ( .A(n_57), .B(n_110), .Y(n_206) );
INVx1_ASAP7_75t_L g150 ( .A(n_58), .Y(n_150) );
INVx1_ASAP7_75t_L g522 ( .A(n_59), .Y(n_522) );
OAI22xp33_ASAP7_75t_L g139 ( .A1(n_60), .A2(n_62), .B1(n_140), .B2(n_142), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_60), .A2(n_474), .B1(n_700), .B2(n_703), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_61), .B(n_162), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_63), .Y(n_666) );
AND2x2_ASAP7_75t_L g220 ( .A(n_65), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g89 ( .A(n_66), .Y(n_89) );
BUFx3_ASAP7_75t_L g124 ( .A(n_66), .Y(n_124) );
INVx1_ASAP7_75t_L g138 ( .A(n_66), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_67), .B(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_68), .B(n_246), .Y(n_245) );
INVx2_ASAP7_75t_L g483 ( .A(n_69), .Y(n_483) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_69), .Y(n_500) );
AND2x2_ASAP7_75t_L g512 ( .A(n_69), .B(n_482), .Y(n_512) );
INVx1_ASAP7_75t_L g488 ( .A(n_70), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_71), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_72), .B(n_110), .Y(n_187) );
OAI21xp5_ASAP7_75t_SL g560 ( .A1(n_73), .A2(n_561), .B(n_577), .Y(n_560) );
INVx2_ASAP7_75t_L g565 ( .A(n_74), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_75), .Y(n_170) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_76), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_96), .B(n_472), .Y(n_77) );
CKINVDCx20_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_86), .Y(n_80) );
BUFx2_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx3_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
INVx2_ASAP7_75t_L g232 ( .A(n_84), .Y(n_232) );
BUFx6f_ASAP7_75t_SL g265 ( .A(n_84), .Y(n_265) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_85), .Y(n_653) );
INVxp67_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AO21x2_ASAP7_75t_L g705 ( .A1(n_87), .A2(n_652), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_90), .Y(n_87) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_88), .A2(n_195), .B(n_196), .Y(n_194) );
BUFx3_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g205 ( .A(n_89), .Y(n_205) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
INVx1_ASAP7_75t_L g211 ( .A(n_94), .Y(n_211) );
INVx2_ASAP7_75t_L g263 ( .A(n_94), .Y(n_263) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g117 ( .A(n_95), .Y(n_117) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
HB1xp67_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NOR2x1_ASAP7_75t_L g98 ( .A(n_99), .B(n_402), .Y(n_98) );
NAND4xp25_ASAP7_75t_L g99 ( .A(n_100), .B(n_309), .C(n_345), .D(n_370), .Y(n_99) );
NOR3xp33_ASAP7_75t_L g100 ( .A(n_101), .B(n_276), .C(n_292), .Y(n_100) );
OAI221xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_188), .B1(n_247), .B2(n_252), .C(n_267), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_152), .Y(n_103) );
INVx2_ASAP7_75t_L g361 ( .A(n_104), .Y(n_361) );
AND2x4_ASAP7_75t_L g393 ( .A(n_104), .B(n_315), .Y(n_393) );
AND2x2_ASAP7_75t_L g471 ( .A(n_104), .B(n_337), .Y(n_471) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_132), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_105), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g335 ( .A(n_105), .Y(n_335) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_106), .B(n_174), .Y(n_269) );
AND2x2_ASAP7_75t_L g295 ( .A(n_106), .B(n_249), .Y(n_295) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_106), .Y(n_313) );
OR2x2_ASAP7_75t_L g317 ( .A(n_106), .B(n_132), .Y(n_317) );
AND2x2_ASAP7_75t_L g330 ( .A(n_106), .B(n_174), .Y(n_330) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_110), .B(n_131), .Y(n_130) );
INVx2_ASAP7_75t_L g168 ( .A(n_110), .Y(n_168) );
INVx1_ASAP7_75t_L g176 ( .A(n_110), .Y(n_176) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g172 ( .A(n_111), .Y(n_172) );
INVx1_ASAP7_75t_L g222 ( .A(n_111), .Y(n_222) );
INVx1_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_125), .B(n_130), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_118), .B(n_122), .Y(n_114) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx3_ASAP7_75t_L g184 ( .A(n_117), .Y(n_184) );
INVx2_ASAP7_75t_L g163 ( .A(n_119), .Y(n_163) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx3_ASAP7_75t_L g128 ( .A(n_120), .Y(n_128) );
INVx3_ASAP7_75t_L g134 ( .A(n_120), .Y(n_134) );
INVx2_ASAP7_75t_L g203 ( .A(n_120), .Y(n_203) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g141 ( .A(n_121), .Y(n_141) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_121), .Y(n_143) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_122), .A2(n_241), .B(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g129 ( .A(n_124), .Y(n_129) );
INVx2_ASAP7_75t_L g162 ( .A(n_124), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B(n_129), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_129), .A2(n_157), .B(n_159), .Y(n_156) );
O2A1O1Ixp5_ASAP7_75t_L g257 ( .A1(n_129), .A2(n_258), .B(n_259), .C(n_260), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g144 ( .A(n_131), .B(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
OR2x2_ASAP7_75t_L g248 ( .A(n_132), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g270 ( .A(n_132), .B(n_251), .Y(n_270) );
BUFx3_ASAP7_75t_L g283 ( .A(n_132), .Y(n_283) );
INVx2_ASAP7_75t_SL g303 ( .A(n_132), .Y(n_303) );
AND2x2_ASAP7_75t_L g344 ( .A(n_132), .B(n_335), .Y(n_344) );
AND2x2_ASAP7_75t_L g367 ( .A(n_132), .B(n_279), .Y(n_367) );
AO31x2_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_135), .A3(n_144), .B(n_149), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_139), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_137), .A2(n_179), .B(n_181), .Y(n_178) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g186 ( .A(n_138), .Y(n_186) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
INVx2_ASAP7_75t_L g201 ( .A(n_141), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_142), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx2_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
AOI21x1_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_148), .Y(n_145) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_146), .A2(n_147), .B(n_148), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_L g312 ( .A(n_152), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_152), .B(n_334), .Y(n_374) );
AND2x2_ASAP7_75t_L g428 ( .A(n_152), .B(n_303), .Y(n_428) );
AND2x2_ASAP7_75t_L g442 ( .A(n_152), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OR2x2_ASAP7_75t_L g408 ( .A(n_153), .B(n_317), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_173), .Y(n_153) );
INVx2_ASAP7_75t_L g251 ( .A(n_154), .Y(n_251) );
BUFx2_ASAP7_75t_SL g291 ( .A(n_154), .Y(n_291) );
AND2x2_ASAP7_75t_L g315 ( .A(n_154), .B(n_174), .Y(n_315) );
INVx1_ASAP7_75t_L g337 ( .A(n_154), .Y(n_337) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_160), .B(n_166), .C(n_169), .Y(n_155) );
INVx2_ASAP7_75t_SL g197 ( .A(n_158), .Y(n_197) );
OAI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_163), .B(n_164), .Y(n_160) );
NAND2x1_ASAP7_75t_L g193 ( .A(n_166), .B(n_194), .Y(n_193) );
AOI21x1_ASAP7_75t_L g198 ( .A1(n_166), .A2(n_199), .B(n_206), .Y(n_198) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_167), .A2(n_178), .B(n_182), .Y(n_177) );
AOI21xp33_ASAP7_75t_L g223 ( .A1(n_167), .A2(n_171), .B(n_220), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVxp67_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx3_ASAP7_75t_L g255 ( .A(n_172), .Y(n_255) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g249 ( .A(n_174), .Y(n_249) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_174), .Y(n_280) );
INVx1_ASAP7_75t_L g302 ( .A(n_174), .Y(n_302) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_177), .B(n_187), .Y(n_174) );
INVx1_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B(n_186), .Y(n_182) );
INVx2_ASAP7_75t_L g236 ( .A(n_184), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_184), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g259 ( .A(n_184), .Y(n_259) );
INVx1_ASAP7_75t_L g214 ( .A(n_186), .Y(n_214) );
OR2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_224), .Y(n_188) );
OR2x2_ASAP7_75t_L g284 ( .A(n_189), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g440 ( .A(n_189), .Y(n_440) );
OR2x2_ASAP7_75t_L g464 ( .A(n_189), .B(n_325), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_207), .Y(n_189) );
AND2x2_ASAP7_75t_L g275 ( .A(n_190), .B(n_208), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_190), .B(n_225), .Y(n_357) );
OR2x2_ASAP7_75t_L g386 ( .A(n_190), .B(n_299), .Y(n_386) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g308 ( .A(n_191), .B(n_208), .Y(n_308) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g253 ( .A(n_192), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g289 ( .A(n_192), .Y(n_289) );
AND2x2_ASAP7_75t_L g369 ( .A(n_192), .B(n_300), .Y(n_369) );
OR2x2_ASAP7_75t_L g422 ( .A(n_192), .B(n_208), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_193), .B(n_198), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_202), .B(n_204), .Y(n_199) );
INVx1_ASAP7_75t_L g219 ( .A(n_204), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_204), .A2(n_262), .B(n_264), .Y(n_261) );
BUFx10_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g298 ( .A(n_207), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g323 ( .A(n_208), .Y(n_323) );
INVx2_ASAP7_75t_L g349 ( .A(n_208), .Y(n_349) );
AND2x2_ASAP7_75t_L g376 ( .A(n_208), .B(n_226), .Y(n_376) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_215), .B(n_223), .Y(n_208) );
NOR2xp67_ASAP7_75t_L g212 ( .A(n_210), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_211), .B(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_219), .B(n_220), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
BUFx2_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g285 ( .A(n_225), .Y(n_285) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g340 ( .A(n_226), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g385 ( .A(n_226), .B(n_349), .Y(n_385) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_227), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g391 ( .A(n_227), .B(n_299), .Y(n_391) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_233), .B(n_239), .Y(n_227) );
AO21x1_ASAP7_75t_SL g274 ( .A1(n_228), .A2(n_233), .B(n_239), .Y(n_274) );
INVxp67_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
OAI21x1_ASAP7_75t_SL g239 ( .A1(n_229), .A2(n_240), .B(n_245), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g246 ( .A(n_230), .Y(n_246) );
INVx2_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
OR2x2_ASAP7_75t_L g290 ( .A(n_248), .B(n_291), .Y(n_290) );
NOR2x1_ASAP7_75t_SL g411 ( .A(n_248), .B(n_291), .Y(n_411) );
INVx2_ASAP7_75t_L g354 ( .A(n_250), .Y(n_354) );
INVx2_ASAP7_75t_L g279 ( .A(n_251), .Y(n_279) );
INVx6_ASAP7_75t_L g328 ( .A(n_252), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_252), .B(n_468), .Y(n_467) );
INVx4_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g375 ( .A(n_253), .B(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_253), .Y(n_444) );
INVx2_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
INVxp33_ASAP7_75t_L g341 ( .A(n_254), .Y(n_341) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_266), .Y(n_254) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_261), .B(n_265), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVxp67_ASAP7_75t_L g387 ( .A(n_269), .Y(n_387) );
AND2x4_ASAP7_75t_L g294 ( .A(n_270), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g332 ( .A(n_271), .Y(n_332) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_272), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g413 ( .A(n_272), .Y(n_413) );
AND2x2_ASAP7_75t_L g420 ( .A(n_272), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g456 ( .A(n_272), .B(n_457), .Y(n_456) );
INVx5_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g347 ( .A(n_273), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g401 ( .A(n_273), .B(n_308), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_273), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g427 ( .A(n_273), .B(n_421), .Y(n_427) );
AND2x4_ASAP7_75t_SL g433 ( .A(n_273), .B(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_273), .B(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVxp67_ASAP7_75t_L g287 ( .A(n_274), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_284), .B1(n_286), .B2(n_290), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_281), .Y(n_277) );
OR2x2_ASAP7_75t_L g395 ( .A(n_278), .B(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g399 ( .A(n_279), .Y(n_399) );
AND2x2_ASAP7_75t_L g462 ( .A(n_279), .B(n_329), .Y(n_462) );
AND2x2_ASAP7_75t_L g380 ( .A(n_280), .B(n_381), .Y(n_380) );
INVxp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g378 ( .A(n_282), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g338 ( .A(n_283), .Y(n_338) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_283), .Y(n_351) );
INVx1_ASAP7_75t_L g396 ( .A(n_283), .Y(n_396) );
AND2x4_ASAP7_75t_L g392 ( .A(n_285), .B(n_308), .Y(n_392) );
OR2x2_ASAP7_75t_L g417 ( .A(n_285), .B(n_368), .Y(n_417) );
OR2x2_ASAP7_75t_L g296 ( .A(n_286), .B(n_297), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x4_ASAP7_75t_L g383 ( .A(n_288), .B(n_298), .Y(n_383) );
INVx1_ASAP7_75t_L g407 ( .A(n_288), .Y(n_407) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g461 ( .A(n_289), .B(n_307), .Y(n_461) );
AND2x2_ASAP7_75t_L g447 ( .A(n_291), .B(n_330), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B1(n_301), .B2(n_304), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_294), .A2(n_433), .B(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g366 ( .A(n_295), .B(n_367), .Y(n_366) );
NAND2x1_ASAP7_75t_L g466 ( .A(n_295), .B(n_399), .Y(n_466) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g348 ( .A(n_299), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g307 ( .A(n_300), .Y(n_307) );
INVx1_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g353 ( .A(n_302), .Y(n_353) );
AOI211x1_ASAP7_75t_L g429 ( .A1(n_302), .A2(n_430), .B(n_435), .C(n_441), .Y(n_429) );
AND2x4_ASAP7_75t_SL g329 ( .A(n_303), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g443 ( .A(n_303), .B(n_335), .Y(n_443) );
INVx2_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AO22x1_ASAP7_75t_L g469 ( .A1(n_305), .A2(n_392), .B1(n_470), .B2(n_471), .Y(n_469) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
OR2x2_ASAP7_75t_L g414 ( .A(n_306), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g432 ( .A(n_306), .Y(n_432) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g436 ( .A(n_307), .B(n_422), .Y(n_436) );
INVx1_ASAP7_75t_L g415 ( .A(n_308), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_318), .B1(n_326), .B2(n_329), .C(n_331), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI221xp5_ASAP7_75t_SL g345 ( .A1(n_312), .A2(n_346), .B1(n_350), .B2(n_355), .C(n_360), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR2x1_ASAP7_75t_L g424 ( .A(n_317), .B(n_337), .Y(n_424) );
INVx2_ASAP7_75t_L g434 ( .A(n_317), .Y(n_434) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_324), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_322), .Y(n_364) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_SL g457 ( .A(n_325), .B(n_451), .Y(n_457) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g418 ( .A(n_329), .Y(n_418) );
AND2x2_ASAP7_75t_L g372 ( .A(n_330), .B(n_337), .Y(n_372) );
OAI22xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B1(n_339), .B2(n_342), .Y(n_331) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g410 ( .A(n_334), .Y(n_410) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g381 ( .A(n_335), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx2_ASAP7_75t_L g343 ( .A(n_337), .Y(n_343) );
AND2x2_ASAP7_75t_L g470 ( .A(n_337), .B(n_434), .Y(n_470) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g446 ( .A(n_340), .B(n_421), .Y(n_446) );
AND2x2_ASAP7_75t_L g359 ( .A(n_341), .B(n_349), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g438 ( .A(n_343), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_343), .B(n_344), .Y(n_455) );
AND2x2_ASAP7_75t_L g398 ( .A(n_344), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_348), .B(n_357), .Y(n_426) );
NAND2xp33_ASAP7_75t_L g449 ( .A(n_348), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
AND2x4_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_356), .B(n_358), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_405), .B(n_408), .C(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B(n_365), .C(n_368), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_377), .C(n_394), .Y(n_370) );
OA21x2_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g465 ( .A(n_372), .Y(n_465) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g445 ( .A(n_376), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B1(n_384), .B2(n_387), .C(n_388), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g468 ( .A(n_385), .Y(n_468) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_392), .B(n_393), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_397), .B(n_400), .Y(n_394) );
INVx1_ASAP7_75t_L g454 ( .A(n_396), .Y(n_454) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
NAND4xp75_ASAP7_75t_L g402 ( .A(n_403), .B(n_429), .C(n_448), .D(n_458), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_412), .B(n_416), .Y(n_403) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g412 ( .A(n_408), .B(n_413), .C(n_414), .Y(n_412) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_409), .A2(n_436), .B1(n_437), .B2(n_439), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_423), .C(n_425), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g451 ( .A(n_422), .Y(n_451) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_424), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_425) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AO32x1_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_444), .A3(n_445), .B1(n_446), .B2(n_447), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_447), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_452), .B1(n_455), .B2(n_456), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI211xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_462), .B(n_463), .C(n_469), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp33_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_465), .B1(n_466), .B2(n_467), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_474), .B1(n_646), .B2(n_656), .C(n_699), .Y(n_472) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_560), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_477), .B(n_521), .C(n_531), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_488), .B1(n_489), .B2(n_496), .C(n_517), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_484), .Y(n_478) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g516 ( .A(n_480), .Y(n_516) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_480), .Y(n_548) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_483), .Y(n_480) );
INVx1_ASAP7_75t_L g501 ( .A(n_481), .Y(n_501) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_481), .Y(n_554) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g505 ( .A(n_482), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_482), .B(n_483), .Y(n_576) );
INVx2_ASAP7_75t_L g506 ( .A(n_483), .Y(n_506) );
AND2x2_ASAP7_75t_L g525 ( .A(n_484), .B(n_504), .Y(n_525) );
AND2x6_ASAP7_75t_L g527 ( .A(n_484), .B(n_499), .Y(n_527) );
AND2x4_ASAP7_75t_L g529 ( .A(n_484), .B(n_530), .Y(n_529) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
AND3x1_ASAP7_75t_L g492 ( .A(n_485), .B(n_493), .C(n_495), .Y(n_492) );
AND2x4_ASAP7_75t_SL g519 ( .A(n_485), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g539 ( .A(n_485), .Y(n_539) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_485), .B(n_520), .Y(n_552) );
OR2x2_ASAP7_75t_L g563 ( .A(n_485), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g494 ( .A(n_487), .Y(n_494) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_488), .A2(n_598), .B1(n_620), .B2(n_622), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx4_ASAP7_75t_L g533 ( .A(n_498), .Y(n_533) );
INVx5_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g558 ( .A(n_500), .Y(n_558) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g518 ( .A(n_504), .B(n_519), .Y(n_518) );
BUFx2_ASAP7_75t_L g534 ( .A(n_504), .Y(n_534) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_513), .B2(n_514), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_508), .A2(n_606), .B1(n_607), .B2(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx4f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_512), .Y(n_530) );
BUFx3_ASAP7_75t_L g546 ( .A(n_512), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_513), .A2(n_522), .B1(n_613), .B2(n_616), .C(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g555 ( .A(n_519), .B(n_556), .Y(n_555) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_526), .B2(n_527), .C1(n_528), .C2(n_529), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_526), .A2(n_528), .B1(n_596), .B2(n_598), .C(n_600), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_535), .A3(n_543), .B1(n_549), .B2(n_550), .C1(n_555), .C2(n_559), .Y(n_531) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g645 ( .A(n_538), .Y(n_645) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_549), .A2(n_624), .B1(n_630), .B2(n_631), .Y(n_623) );
INVx5_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OR2x6_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OR2x2_ASAP7_75t_L g574 ( .A(n_552), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_567), .B(n_574), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g579 ( .A(n_564), .B(n_580), .Y(n_579) );
OR2x6_ASAP7_75t_SL g583 ( .A(n_564), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g590 ( .A(n_564), .Y(n_590) );
OR2x6_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
BUFx2_ASAP7_75t_L g603 ( .A(n_565), .Y(n_603) );
INVx1_ASAP7_75t_L g629 ( .A(n_565), .Y(n_629) );
INVx1_ASAP7_75t_L g604 ( .A(n_566), .Y(n_604) );
AND2x4_ASAP7_75t_L g618 ( .A(n_566), .B(n_603), .Y(n_618) );
AND2x2_ASAP7_75t_L g628 ( .A(n_566), .B(n_629), .Y(n_628) );
OR2x2_ASAP7_75t_L g685 ( .A(n_566), .B(n_629), .Y(n_685) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx12f_ASAP7_75t_L g599 ( .A(n_570), .Y(n_599) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x4_ASAP7_75t_L g581 ( .A(n_571), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g611 ( .A(n_571), .Y(n_611) );
AND2x4_ASAP7_75t_L g585 ( .A(n_572), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g593 ( .A(n_573), .B(n_586), .Y(n_593) );
AND2x2_ASAP7_75t_L g640 ( .A(n_573), .B(n_587), .Y(n_640) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI31xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_594), .A3(n_635), .B(n_645), .Y(n_577) );
BUFx3_ASAP7_75t_L g607 ( .A(n_580), .Y(n_607) );
BUFx3_ASAP7_75t_L g616 ( .A(n_580), .Y(n_616) );
INVx8_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g610 ( .A(n_582), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g625 ( .A(n_582), .Y(n_625) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_585), .Y(n_597) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_585), .Y(n_615) );
INVx1_ASAP7_75t_L g633 ( .A(n_586), .Y(n_633) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx4_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g594 ( .A1(n_595), .A2(n_605), .B1(n_612), .B2(n_619), .C(n_623), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
BUFx3_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g621 ( .A(n_609), .Y(n_621) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_SL g690 ( .A(n_624), .Y(n_690) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g681 ( .A(n_625), .B(n_682), .C(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g634 ( .A(n_627), .Y(n_634) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g641 ( .A(n_628), .Y(n_641) );
AND2x4_ASAP7_75t_L g631 ( .A(n_632), .B(n_634), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx3_ASAP7_75t_L g643 ( .A(n_641), .Y(n_643) );
OR2x6_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
CKINVDCx16_ASAP7_75t_R g646 ( .A(n_647), .Y(n_646) );
CKINVDCx16_ASAP7_75t_R g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_654), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g679 ( .A(n_653), .Y(n_679) );
AND2x2_ASAP7_75t_L g706 ( .A(n_654), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_655), .B(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_673), .B1(n_691), .B2(n_693), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_657), .A2(n_691), .B1(n_701), .B2(n_702), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_664), .B2(n_672), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_660), .Y(n_663) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g672 ( .A(n_664), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g671 ( .A(n_669), .Y(n_671) );
INVx3_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx3_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx5_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g701 ( .A(n_676), .Y(n_701) );
AND2x6_ASAP7_75t_L g676 ( .A(n_677), .B(n_686), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVxp67_ASAP7_75t_L g697 ( .A(n_678), .Y(n_697) );
INVx1_ASAP7_75t_L g707 ( .A(n_679), .Y(n_707) );
INVxp67_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_681), .B(n_690), .Y(n_698) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
CKINVDCx11_ASAP7_75t_R g688 ( .A(n_683), .Y(n_688) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_687), .B(n_689), .Y(n_686) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx3_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx4f_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
BUFx3_ASAP7_75t_L g702 ( .A(n_695), .Y(n_702) );
INVx4_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_704), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_705), .Y(n_704) );
endmodule