module fake_jpeg_27904_n_141 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_141);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_141;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_7),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_69),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_52),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_64),
.Y(n_73)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_50),
.B1(n_53),
.B2(n_46),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_70),
.A2(n_71),
.B1(n_61),
.B2(n_48),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_57),
.B1(n_45),
.B2(n_55),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_44),
.B1(n_60),
.B2(n_48),
.Y(n_74)
);

OR2x4_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_81),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_77),
.Y(n_87)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_43),
.B1(n_51),
.B2(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_60),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_45),
.B1(n_57),
.B2(n_62),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_61),
.B(n_45),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_86),
.B1(n_90),
.B2(n_4),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_0),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_98),
.B(n_3),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_73),
.B(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_97),
.Y(n_102)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_44),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_83),
.C(n_72),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_104),
.B(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_26),
.B1(n_41),
.B2(n_39),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_90),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_106),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_91),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_101),
.C(n_87),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_111),
.B(n_112),
.Y(n_118)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_28),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_27),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_20),
.Y(n_126)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_114),
.Y(n_119)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_96),
.B1(n_100),
.B2(n_103),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_125),
.B1(n_89),
.B2(n_5),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_117),
.B(n_121),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_25),
.B(n_42),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_16),
.B1(n_36),
.B2(n_35),
.C(n_33),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_126),
.B1(n_19),
.B2(n_38),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_100),
.B1(n_89),
.B2(n_24),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_125),
.C(n_117),
.Y(n_133)
);

AO21x1_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_130),
.B(n_118),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_131),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_122),
.C(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_130),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_10),
.C(n_32),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_37),
.C(n_29),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_15),
.Y(n_141)
);


endmodule