module fake_jpeg_20132_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_6),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_58),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_67),
.B1(n_53),
.B2(n_74),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_67),
.B1(n_58),
.B2(n_61),
.Y(n_100)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_75),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_2),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_102),
.B1(n_108),
.B2(n_111),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_77),
.C(n_68),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_109),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_76),
.B1(n_57),
.B2(n_55),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_51),
.B(n_72),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_103),
.A2(n_55),
.B1(n_54),
.B2(n_69),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_73),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_63),
.B1(n_56),
.B2(n_66),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_32),
.B(n_42),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_70),
.B1(n_60),
.B2(n_66),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_122),
.C(n_3),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_110),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_121),
.Y(n_131)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_70),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_65),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_64),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_2),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_65),
.C(n_102),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_129),
.C(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_64),
.C(n_54),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_112),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_23),
.B(n_45),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_28),
.B(n_13),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_18),
.C(n_44),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_9),
.B1(n_14),
.B2(n_15),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_5),
.B(n_7),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_142),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_146),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_148),
.B1(n_146),
.B2(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_150),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_148)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_130),
.C(n_129),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_153),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_166),
.B(n_155),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_159),
.B(n_156),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_162),
.Y(n_169)
);

AOI321xp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_154),
.A3(n_33),
.B1(n_35),
.B2(n_38),
.C(n_29),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_39),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_43),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_49),
.Y(n_173)
);


endmodule