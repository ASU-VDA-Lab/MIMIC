module fake_jpeg_21301_n_98 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_29),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_51),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_45),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_38),
.B1(n_46),
.B2(n_44),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_56),
.A2(n_59),
.B1(n_37),
.B2(n_1),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_38),
.B1(n_43),
.B2(n_39),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_3),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_57),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_70),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_36),
.B1(n_1),
.B2(n_2),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_62),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_72),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_18),
.C(n_32),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_SL g78 ( 
.A(n_71),
.B(n_74),
.C(n_15),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_17),
.C(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_2),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_3),
.B(n_4),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_16),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_19),
.C(n_30),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_80),
.C(n_20),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

XNOR2x1_ASAP7_75t_L g85 ( 
.A(n_83),
.B(n_73),
.Y(n_85)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_4),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_89),
.B1(n_79),
.B2(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_81),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_87),
.B(n_77),
.C(n_82),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_84),
.B1(n_5),
.B2(n_12),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_34),
.C(n_8),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_13),
.B(n_23),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_25),
.B(n_28),
.Y(n_98)
);


endmodule