module fake_jpeg_27161_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_SL g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_21),
.B(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_46),
.A2(n_51),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_50),
.B(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_58),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_56),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_36),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_79),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_44),
.B1(n_60),
.B2(n_52),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_70),
.B1(n_84),
.B2(n_88),
.Y(n_115)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_44),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_40),
.C(n_38),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_23),
.B1(n_37),
.B2(n_18),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_92),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_76),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_18),
.B1(n_25),
.B2(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_65),
.B1(n_68),
.B2(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_32),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_41),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_83),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_41),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_85),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_42),
.B1(n_41),
.B2(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_90),
.Y(n_124)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_30),
.B1(n_29),
.B2(n_16),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_91),
.A2(n_96),
.B1(n_27),
.B2(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_40),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_53),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_19),
.B1(n_24),
.B2(n_33),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_97),
.B1(n_24),
.B2(n_33),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_52),
.A2(n_24),
.B1(n_19),
.B2(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_31),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_62),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_99),
.B(n_101),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_125),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_69),
.A2(n_0),
.B(n_1),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_40),
.C(n_38),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_121),
.C(n_126),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_38),
.A3(n_36),
.B1(n_43),
.B2(n_17),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_70),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_0),
.B(n_1),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_38),
.B(n_36),
.C(n_43),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_122),
.B1(n_85),
.B2(n_86),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_17),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_L g123 ( 
.A(n_64),
.B(n_36),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_123),
.B(n_71),
.Y(n_136)
);

OAI22x1_ASAP7_75t_L g125 ( 
.A1(n_63),
.A2(n_27),
.B1(n_31),
.B2(n_28),
.Y(n_125)
);

OAI22x1_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_80),
.B1(n_66),
.B2(n_83),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_31),
.B(n_12),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_135),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_142),
.Y(n_164)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_136),
.B(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_117),
.B1(n_106),
.B2(n_104),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_96),
.B1(n_93),
.B2(n_77),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_143),
.B1(n_102),
.B2(n_113),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_139),
.A2(n_112),
.B1(n_100),
.B2(n_104),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_88),
.B1(n_81),
.B2(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_152),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_82),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_87),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_148),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_66),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

OA21x2_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_112),
.B(n_106),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_28),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_20),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_72),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_157)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_20),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_124),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_174),
.B(n_181),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_166),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_121),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_183),
.B1(n_184),
.B2(n_175),
.Y(n_210)
);

AOI22x1_ASAP7_75t_SL g170 ( 
.A1(n_151),
.A2(n_125),
.B1(n_109),
.B2(n_114),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_170),
.A2(n_185),
.B1(n_141),
.B2(n_140),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_102),
.B1(n_122),
.B2(n_119),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_171),
.A2(n_186),
.B1(n_187),
.B2(n_10),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_130),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_177),
.B(n_188),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_101),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_140),
.B(n_150),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_2),
.B(n_3),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_10),
.C(n_14),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g192 ( 
.A1(n_170),
.A2(n_157),
.B1(n_143),
.B2(n_133),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_135),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_197),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_196),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_160),
.B(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_157),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_209),
.Y(n_236)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_203),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_142),
.Y(n_204)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_152),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_214),
.B1(n_215),
.B2(n_218),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_220),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_150),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_165),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_169),
.B1(n_180),
.B2(n_171),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_15),
.A3(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_216),
.A2(n_176),
.B(n_185),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_172),
.B(n_15),
.Y(n_217)
);

NOR4xp25_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_11),
.C(n_3),
.D(n_4),
.Y(n_242)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_2),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_219),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_169),
.B(n_11),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_221),
.A2(n_187),
.B1(n_182),
.B2(n_175),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_223),
.A2(n_216),
.B1(n_219),
.B2(n_215),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_228),
.A2(n_231),
.B(n_240),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_190),
.B(n_182),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_229),
.B(n_242),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_191),
.C(n_186),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_178),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_235),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_210),
.C(n_198),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_198),
.C(n_214),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_163),
.B(n_179),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_193),
.B(n_163),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_220),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_179),
.B(n_3),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_200),
.B1(n_4),
.B2(n_5),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_208),
.C(n_205),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_247),
.C(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_206),
.C(n_209),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_192),
.B1(n_211),
.B2(n_204),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_256),
.B1(n_227),
.B2(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_254),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_236),
.B(n_197),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_192),
.B1(n_211),
.B2(n_201),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_255),
.A2(n_257),
.B1(n_223),
.B2(n_232),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_194),
.B1(n_201),
.B2(n_211),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

XOR2x2_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_221),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_234),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_257),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_241),
.C(n_240),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_248),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_247),
.C(n_250),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_230),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_224),
.C(n_225),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_243),
.B(n_232),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_251),
.Y(n_285)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_230),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_268),
.A2(n_252),
.B(n_224),
.Y(n_281)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_249),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_226),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_286),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_276),
.Y(n_296)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_288),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_226),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_271),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_290),
.A2(n_284),
.B1(n_269),
.B2(n_270),
.Y(n_297)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_278),
.A2(n_248),
.B(n_4),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_299),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_272),
.C(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_272),
.C(n_273),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_6),
.C(n_304),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_286),
.A2(n_266),
.B(n_274),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_303),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_265),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_306),
.B(n_311),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_291),
.A3(n_290),
.B1(n_293),
.B2(n_285),
.C1(n_5),
.C2(n_2),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_307),
.A2(n_298),
.B(n_310),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_5),
.B1(n_6),
.B2(n_296),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_6),
.B(n_300),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_312),
.B(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_313),
.Y(n_317)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_298),
.B(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_316),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_315),
.B(n_312),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_317),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_308),
.Y(n_322)
);


endmodule