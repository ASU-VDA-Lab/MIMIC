module fake_jpeg_7871_n_228 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_36),
.Y(n_52)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_14),
.B(n_21),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_34),
.B(n_38),
.C(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_15),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_25),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_29),
.B(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_23),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_27),
.B1(n_23),
.B2(n_18),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_15),
.B1(n_19),
.B2(n_18),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_36),
.B1(n_33),
.B2(n_39),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_63),
.B1(n_67),
.B2(n_55),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_59),
.A2(n_60),
.B1(n_43),
.B2(n_49),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_36),
.B1(n_39),
.B2(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_24),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_74),
.B(n_56),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_30),
.B1(n_23),
.B2(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_71),
.Y(n_87)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_72),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_77),
.B(n_79),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_88),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_31),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_48),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_86),
.B(n_91),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_48),
.B(n_56),
.C(n_51),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_SL g95 ( 
.A(n_85),
.B(n_66),
.C(n_73),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_43),
.B(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_95),
.A2(n_101),
.B1(n_107),
.B2(n_88),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_105),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_38),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_1),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_66),
.B(n_73),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_86),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_1),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_42),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_90),
.C(n_84),
.Y(n_123)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_110),
.A2(n_76),
.B1(n_93),
.B2(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_85),
.B1(n_76),
.B2(n_31),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_78),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_113),
.B(n_115),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_91),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_114),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_124),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_117),
.B(n_120),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_118),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_137)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_101),
.C(n_102),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_126),
.B(n_108),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_128),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_75),
.C(n_68),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_121),
.A2(n_100),
.B(n_99),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_136),
.B(n_137),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_103),
.B1(n_100),
.B2(n_109),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_138),
.A2(n_140),
.B1(n_148),
.B2(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_109),
.B1(n_95),
.B2(n_101),
.Y(n_140)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_147),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_105),
.B1(n_76),
.B2(n_107),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_120),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_153),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_163),
.C(n_165),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_123),
.B1(n_116),
.B2(n_130),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_166),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_161),
.B(n_144),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_125),
.B1(n_75),
.B2(n_64),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_125),
.B1(n_68),
.B2(n_14),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_150),
.C(n_145),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_135),
.C(n_147),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_181),
.C(n_182),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_16),
.B1(n_14),
.B2(n_20),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_159),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_20),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_150),
.C(n_64),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_40),
.C(n_53),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_184),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_173),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_189),
.B1(n_193),
.B2(n_21),
.Y(n_203)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_192),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_179),
.A2(n_151),
.B1(n_53),
.B2(n_40),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_191),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_2),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_12),
.B1(n_13),
.B2(n_20),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_12),
.Y(n_199)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_172),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_181),
.C(n_168),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_187),
.C(n_193),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

OAI321xp33_ASAP7_75t_L g207 ( 
.A1(n_198),
.A2(n_202),
.A3(n_192),
.B1(n_21),
.B2(n_16),
.C(n_38),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_3),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_13),
.B1(n_20),
.B2(n_16),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_203),
.A2(n_195),
.B(n_200),
.C(n_183),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_207),
.Y(n_213)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_4),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_201),
.A2(n_21),
.B1(n_16),
.B2(n_7),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_3),
.C(n_4),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_203),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_3),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_4),
.Y(n_215)
);

AOI31xp67_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_206),
.A3(n_211),
.B(n_201),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_7),
.C(n_8),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_218),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_221),
.B(n_222),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_213),
.C(n_215),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_53),
.C(n_10),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_224),
.B(n_10),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_8),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_11),
.Y(n_228)
);


endmodule