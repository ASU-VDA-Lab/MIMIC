module real_jpeg_30859_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_682, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_682;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_553;
wire n_290;
wire n_121;
wire n_234;
wire n_666;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_634;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_667;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_0),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g368 ( 
.A(n_0),
.Y(n_368)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_0),
.Y(n_639)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_2),
.A2(n_103),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_2),
.A2(n_103),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_2),
.A2(n_103),
.B1(n_370),
.B2(n_374),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_66),
.B1(n_91),
.B2(n_94),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_3),
.A2(n_66),
.B1(n_168),
.B2(n_172),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_3),
.A2(n_66),
.B1(n_309),
.B2(n_314),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_4),
.A2(n_154),
.B1(n_155),
.B2(n_160),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_4),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_4),
.A2(n_154),
.B1(n_249),
.B2(n_252),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_4),
.A2(n_154),
.B1(n_410),
.B2(n_414),
.Y(n_409)
);

AO22x1_ASAP7_75t_L g467 ( 
.A1(n_4),
.A2(n_154),
.B1(n_363),
.B2(n_468),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_5),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_5),
.A2(n_182),
.B1(n_225),
.B2(n_228),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_5),
.A2(n_160),
.B1(n_182),
.B2(n_272),
.Y(n_271)
);

AO22x1_ASAP7_75t_L g360 ( 
.A1(n_5),
.A2(n_182),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_6),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_7),
.A2(n_54),
.B1(n_57),
.B2(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_7),
.A2(n_60),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_7),
.A2(n_60),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_7),
.A2(n_60),
.B1(n_277),
.B2(n_282),
.Y(n_276)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_8),
.Y(n_96)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_8),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_9),
.Y(n_195)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_10),
.A2(n_54),
.B1(n_397),
.B2(n_398),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_10),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_10),
.A2(n_397),
.B1(n_450),
.B2(n_452),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_10),
.A2(n_397),
.B1(n_542),
.B2(n_546),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g631 ( 
.A1(n_10),
.A2(n_397),
.B1(n_632),
.B2(n_634),
.Y(n_631)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_11),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_12),
.A2(n_258),
.B1(n_259),
.B2(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_12),
.A2(n_258),
.B1(n_381),
.B2(n_384),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_12),
.A2(n_134),
.B1(n_258),
.B2(n_500),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_SL g571 ( 
.A1(n_12),
.A2(n_258),
.B1(n_572),
.B2(n_575),
.Y(n_571)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_13),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_14),
.B(n_678),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_14),
.B(n_680),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_15),
.Y(n_106)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_15),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_15),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_16),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_16),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_16),
.A2(n_150),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_16),
.A2(n_150),
.B1(n_432),
.B2(n_433),
.Y(n_431)
);

OAI22x1_ASAP7_75t_L g526 ( 
.A1(n_16),
.A2(n_150),
.B1(n_527),
.B2(n_529),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_17),
.B(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_17),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_17),
.B(n_63),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_SL g550 ( 
.A1(n_17),
.A2(n_446),
.B1(n_551),
.B2(n_553),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_17),
.B(n_216),
.Y(n_569)
);

OAI21xp33_ASAP7_75t_L g645 ( 
.A1(n_17),
.A2(n_237),
.B(n_580),
.Y(n_645)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_18),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_18),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_72),
.B(n_676),
.C(n_679),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_22),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_52),
.B1(n_61),
.B2(n_64),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_23),
.A2(n_61),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_24),
.A2(n_62),
.B(n_65),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_24),
.A2(n_62),
.B1(n_153),
.B2(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_24),
.A2(n_53),
.B1(n_62),
.B2(n_329),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_25),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_25),
.B(n_257),
.Y(n_256)
);

AO22x1_ASAP7_75t_L g421 ( 
.A1(n_25),
.A2(n_63),
.B1(n_257),
.B2(n_396),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_25),
.B(n_442),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_42),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_34),
.B2(n_38),
.Y(n_26)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_27),
.Y(n_398)
);

INVx4_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_29),
.Y(n_151)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_29),
.Y(n_445)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_37),
.Y(n_149)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_37),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_37),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_41),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_41),
.Y(n_358)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_48),
.B2(n_50),
.Y(n_42)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_44),
.Y(n_253)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_45),
.Y(n_392)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_46),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_47),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_47),
.Y(n_281)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_48),
.Y(n_554)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g264 ( 
.A(n_56),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_59),
.Y(n_161)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_63),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_63),
.B(n_146),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_63),
.B(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_71),
.B(n_333),
.Y(n_678)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AO21x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_334),
.B(n_665),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_319),
.C(n_330),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_290),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_266),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_77),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_163),
.C(n_219),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_78),
.B(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_142),
.Y(n_78)
);

OA21x2_ASAP7_75t_SL g289 ( 
.A1(n_79),
.A2(n_144),
.B(n_162),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_97),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_80),
.A2(n_143),
.B1(n_144),
.B2(n_162),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_80),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_80),
.A2(n_97),
.B1(n_162),
.B2(n_480),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B(n_90),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_82),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_84),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_84),
.A2(n_360),
.B1(n_365),
.B2(n_369),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_84),
.A2(n_360),
.B1(n_365),
.B2(n_467),
.Y(n_466)
);

NAND2x1_ASAP7_75t_SL g525 ( 
.A(n_84),
.B(n_526),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_87),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_87),
.Y(n_244)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_87),
.Y(n_373)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_87),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_87),
.Y(n_592)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_89),
.Y(n_649)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_90),
.Y(n_236)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_93),
.Y(n_377)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_93),
.Y(n_633)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_95),
.Y(n_364)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_95),
.Y(n_528)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_96),
.Y(n_609)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_97),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_107),
.B1(n_133),
.B2(n_141),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_98),
.A2(n_107),
.B1(n_141),
.B2(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_106),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_106),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_106),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_106),
.Y(n_614)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_107),
.A2(n_141),
.B1(n_224),
.B2(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_107),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_107),
.A2(n_141),
.B1(n_499),
.B2(n_541),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_107),
.A2(n_541),
.B1(n_566),
.B2(n_567),
.Y(n_565)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_120),
.Y(n_107)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

OAI22x1_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_116),
.B2(n_118),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_115),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_124),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_125),
.Y(n_438)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_132),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_132),
.Y(n_545)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_137),
.Y(n_432)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_140),
.Y(n_515)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_140),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_145),
.B(n_395),
.Y(n_394)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_157),
.Y(n_273)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_163),
.B(n_220),
.Y(n_476)
);

XNOR2x1_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_176),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_164),
.B(n_176),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_164),
.B(n_176),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_167),
.B2(n_175),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_165),
.A2(n_167),
.B(n_175),
.Y(n_284)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_175),
.A2(n_430),
.B1(n_431),
.B2(n_439),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_175),
.B(n_431),
.Y(n_502)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_175),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_188),
.B1(n_209),
.B2(n_216),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_188),
.B1(n_218),
.B2(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_179),
.Y(n_451)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_180),
.Y(n_552)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_181),
.Y(n_346)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_187),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_187),
.Y(n_251)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_187),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_187),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_188),
.A2(n_209),
.B1(n_216),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_188),
.A2(n_216),
.B1(n_276),
.B2(n_308),
.Y(n_307)
);

OA21x2_ASAP7_75t_SL g327 ( 
.A1(n_188),
.A2(n_216),
.B(n_308),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_188),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_188),
.A2(n_216),
.B1(n_449),
.B2(n_454),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g464 ( 
.A(n_188),
.B(n_388),
.Y(n_464)
);

AND2x4_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_202),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_192),
.B1(n_196),
.B2(n_199),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_193),
.Y(n_521)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_198),
.Y(n_203)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_199),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_199),
.Y(n_355)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

INVx5_ASAP7_75t_L g519 ( 
.A(n_200),
.Y(n_519)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_201),
.Y(n_453)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_204),
.Y(n_500)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

OAI22x1_ASAP7_75t_L g418 ( 
.A1(n_217),
.A2(n_386),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_217),
.A2(n_463),
.B(n_464),
.Y(n_462)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_218),
.B(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_245),
.C(n_254),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_222),
.B(n_485),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_223),
.Y(n_401)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_227),
.Y(n_507)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2x2_ASAP7_75t_L g400 ( 
.A(n_232),
.B(n_401),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_237),
.A2(n_238),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_237),
.A2(n_571),
.B(n_580),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_237),
.A2(n_571),
.B1(n_631),
.B2(n_648),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_240),
.Y(n_362)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_247),
.B(n_255),
.Y(n_485)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_248),
.Y(n_420)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_251),
.Y(n_385)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_265),
.B(n_441),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_266),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_289),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_267)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_280),
.Y(n_383)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_284),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_294),
.C(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.C(n_289),
.Y(n_291)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_290),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_291),
.Y(n_672)
);

INVxp33_ASAP7_75t_L g671 ( 
.A(n_292),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_294),
.A2(n_297),
.B1(n_298),
.B2(n_318),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_305),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_299),
.B(n_306),
.C(n_325),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_321),
.C(n_322),
.Y(n_320)
);

OAI321xp33_ASAP7_75t_L g665 ( 
.A1(n_319),
.A2(n_666),
.A3(n_667),
.B1(n_670),
.B2(n_673),
.C(n_682),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_320),
.B(n_323),
.Y(n_674)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_327),
.C(n_328),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND3xp33_ASAP7_75t_L g667 ( 
.A(n_331),
.B(n_668),
.C(n_669),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g670 ( 
.A(n_331),
.B(n_671),
.C(n_672),
.Y(n_670)
);

AOI21xp33_ASAP7_75t_SL g673 ( 
.A1(n_331),
.A2(n_674),
.B(n_675),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_332),
.B(n_333),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_656),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_490),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_473),
.Y(n_336)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_422),
.B(n_455),
.Y(n_337)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_338),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_399),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_339),
.B(n_400),
.C(n_402),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_378),
.C(n_393),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_340),
.B(n_425),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_359),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_341),
.B(n_359),
.Y(n_459)
);

AOI32xp33_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_347),
.A3(n_350),
.B1(n_351),
.B2(n_354),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_346),
.Y(n_389)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_351),
.Y(n_447)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_366),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx8_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_376),
.Y(n_574)
);

INVx4_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_378),
.A2(n_379),
.B1(n_393),
.B2(n_394),
.Y(n_425)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_386),
.B(n_387),
.Y(n_379)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_386),
.A2(n_387),
.B(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_402),
.Y(n_399)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_417),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_403),
.B(n_418),
.C(n_421),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_408),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_406),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_407),
.Y(n_581)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx4_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_416),
.Y(n_622)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_421),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_423),
.B(n_659),
.C(n_660),
.Y(n_658)
);

MAJx2_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_426),
.C(n_427),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_424),
.B(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_426),
.B(n_428),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_440),
.C(n_448),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_429),
.B(n_448),
.Y(n_458)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_431),
.Y(n_566)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_438),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_440),
.B(n_458),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_446),
.B(n_447),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_446),
.B(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_512),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_446),
.B(n_602),
.Y(n_601)
);

OA21x2_ASAP7_75t_R g620 ( 
.A1(n_446),
.A2(n_601),
.B(n_621),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_446),
.B(n_567),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_446),
.B(n_644),
.Y(n_643)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_449),
.Y(n_463)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_471),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_456),
.B(n_471),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.C(n_460),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_457),
.B(n_535),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_459),
.B(n_460),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.C(n_466),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_462),
.B(n_496),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_466),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_467),
.B(n_524),
.Y(n_523)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_468),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_468),
.B(n_643),
.Y(n_642)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_473),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_477),
.B(n_486),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_474),
.B(n_477),
.Y(n_664)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_475),
.B(n_478),
.Y(n_663)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_481),
.C(n_483),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_484),
.Y(n_488)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_488),
.Y(n_487)
);

INVxp33_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_487),
.B(n_489),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_491),
.A2(n_536),
.B(n_654),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_534),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_493),
.B(n_655),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_497),
.C(n_503),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_495),
.B(n_559),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_497),
.A2(n_498),
.B1(n_503),
.B2(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_501),
.B(n_502),
.Y(n_498)
);

OA21x2_ASAP7_75t_SL g619 ( 
.A1(n_501),
.A2(n_502),
.B(n_620),
.Y(n_619)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_503),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_522),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_504),
.B(n_522),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_505),
.A2(n_508),
.B1(n_511),
.B2(n_516),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_520),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

NAND2x1_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_525),
.A2(n_631),
.B(n_635),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g580 ( 
.A(n_526),
.B(n_581),
.Y(n_580)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_533),
.Y(n_579)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_534),
.Y(n_655)
);

AOI21x1_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_586),
.B(n_653),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_561),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_558),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_539),
.B(n_558),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_548),
.C(n_555),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_540),
.B(n_549),
.Y(n_584)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_556),
.A2(n_557),
.B1(n_583),
.B2(n_584),
.Y(n_582)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_585),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_582),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_582),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_568),
.C(n_570),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_565),
.B(n_569),
.Y(n_625)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_581),
.Y(n_644)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_585),
.B(n_652),
.Y(n_651)
);

AO21x1_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_626),
.B(n_651),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_588),
.B(n_623),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_588),
.B(n_623),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_619),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_589),
.B(n_619),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_590),
.A2(n_600),
.B1(n_605),
.B2(n_610),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_591),
.B(n_593),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_615),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_625),
.Y(n_623)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_628),
.B(n_647),
.C(n_650),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_629),
.A2(n_641),
.B(n_646),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_640),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_630),
.B(n_640),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_633),
.Y(n_632)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_638),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_642),
.B(n_645),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_649),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_657),
.A2(n_658),
.B(n_661),
.Y(n_656)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_662),
.A2(n_663),
.B(n_664),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g676 ( 
.A(n_677),
.Y(n_676)
);


endmodule