module fake_jpeg_448_n_686 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_19),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_16),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_8),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_4),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_2),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_60),
.Y(n_213)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_62),
.Y(n_218)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g197 ( 
.A(n_66),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_70),
.B(n_75),
.Y(n_177)
);

BUFx12f_ASAP7_75t_SL g71 ( 
.A(n_23),
.Y(n_71)
);

HAxp5_ASAP7_75t_SL g201 ( 
.A(n_71),
.B(n_52),
.CON(n_201),
.SN(n_201)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_72),
.B(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_10),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_77),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_79),
.B(n_105),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_80),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx5_ASAP7_75t_SL g203 ( 
.A(n_81),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_36),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_84),
.B(n_91),
.Y(n_165)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_23),
.Y(n_85)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_86),
.Y(n_192)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_31),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_107),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_94),
.Y(n_147)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_95),
.Y(n_187)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_97),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_98),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_100),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_10),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_101),
.B(n_29),
.C(n_0),
.Y(n_195)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_102),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx16f_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_42),
.B(n_10),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_31),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_108),
.Y(n_232)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_55),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_111),
.B(n_123),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_38),
.Y(n_112)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_42),
.B(n_12),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_113),
.B(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_53),
.B(n_12),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_41),
.Y(n_119)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_31),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_38),
.Y(n_124)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_125),
.Y(n_196)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_126),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_33),
.Y(n_127)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_129),
.Y(n_221)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_130),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_41),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_132),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_81),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_134),
.B(n_169),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_67),
.A2(n_49),
.B1(n_39),
.B2(n_43),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_138),
.A2(n_160),
.B1(n_217),
.B2(n_230),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_69),
.A2(n_49),
.B1(n_39),
.B2(n_58),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_149),
.A2(n_152),
.B1(n_155),
.B2(n_157),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_76),
.A2(n_43),
.B1(n_35),
.B2(n_39),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_78),
.A2(n_35),
.B1(n_39),
.B2(n_49),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_62),
.A2(n_49),
.B1(n_50),
.B2(n_58),
.Y(n_156)
);

OA22x2_ASAP7_75t_L g291 ( 
.A1(n_156),
.A2(n_161),
.B1(n_173),
.B2(n_202),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_101),
.A2(n_56),
.B1(n_27),
.B2(n_47),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_104),
.A2(n_56),
.B(n_27),
.C(n_47),
.Y(n_159)
);

HAxp5_ASAP7_75t_SL g314 ( 
.A(n_159),
.B(n_201),
.CON(n_314),
.SN(n_314)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_80),
.A2(n_92),
.B1(n_129),
.B2(n_127),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_104),
.A2(n_21),
.B1(n_46),
.B2(n_45),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_60),
.B(n_44),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_82),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_206),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_59),
.A2(n_40),
.B1(n_52),
.B2(n_45),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_90),
.A2(n_40),
.B1(n_21),
.B2(n_46),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_174),
.A2(n_176),
.B1(n_200),
.B2(n_215),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_94),
.A2(n_44),
.B1(n_34),
.B2(n_30),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_99),
.A2(n_34),
.B1(n_30),
.B2(n_29),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_182),
.A2(n_141),
.B1(n_173),
.B2(n_175),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_18),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_0),
.B1(n_1),
.B2(n_52),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_130),
.A2(n_12),
.B1(n_17),
.B2(n_2),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_64),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_68),
.A2(n_9),
.B1(n_17),
.B2(n_2),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_208),
.A2(n_168),
.B1(n_170),
.B2(n_104),
.Y(n_318)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_85),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_83),
.B(n_9),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_220),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_116),
.A2(n_9),
.B1(n_16),
.B2(n_3),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_98),
.B(n_18),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_117),
.A2(n_7),
.B1(n_15),
.B2(n_3),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_97),
.B(n_13),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_112),
.A2(n_124),
.B1(n_102),
.B2(n_100),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_222),
.A2(n_121),
.B1(n_1),
.B2(n_15),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_132),
.B(n_13),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_223),
.B(n_224),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_86),
.B(n_4),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_132),
.Y(n_225)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_98),
.Y(n_228)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_228),
.Y(n_266)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_110),
.Y(n_229)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_110),
.A2(n_4),
.B1(n_7),
.B2(n_14),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_131),
.B(n_4),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_119),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_197),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_233),
.B(n_245),
.Y(n_324)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_235),
.Y(n_320)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_236),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_237),
.B(n_293),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_224),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_238),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_154),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g339 ( 
.A(n_240),
.B(n_265),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_241),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_243),
.Y(n_322)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_184),
.Y(n_244)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_244),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_140),
.Y(n_245)
);

INVx3_ASAP7_75t_SL g246 ( 
.A(n_139),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_246),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_247),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_248),
.B(n_257),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_188),
.B(n_0),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_249),
.B(n_261),
.Y(n_327)
);

AND2x2_ASAP7_75t_SL g250 ( 
.A(n_201),
.B(n_131),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_250),
.Y(n_331)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_142),
.Y(n_252)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

OR2x2_ASAP7_75t_SL g254 ( 
.A(n_189),
.B(n_119),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_254),
.Y(n_349)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_197),
.Y(n_255)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_255),
.Y(n_333)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_136),
.B(n_151),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_179),
.B(n_0),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_197),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_262),
.B(n_264),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_181),
.A2(n_222),
.B(n_156),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_263),
.A2(n_305),
.B(n_309),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_165),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_135),
.B(n_121),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_268),
.A2(n_289),
.B1(n_258),
.B2(n_243),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_269),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_180),
.B(n_1),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_285),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_145),
.Y(n_271)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_271),
.Y(n_350)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_143),
.Y(n_272)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_272),
.Y(n_341)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_163),
.Y(n_274)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

OR2x2_ASAP7_75t_SL g277 ( 
.A(n_177),
.B(n_14),
.Y(n_277)
);

AOI21xp33_ASAP7_75t_L g344 ( 
.A1(n_277),
.A2(n_302),
.B(n_307),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_278),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_137),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_279),
.B(n_284),
.Y(n_353)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_280),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_219),
.Y(n_281)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_281),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_283),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_173),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_191),
.B(n_1),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_198),
.B(n_14),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_286),
.B(n_294),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_138),
.A2(n_15),
.B1(n_152),
.B2(n_155),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_287),
.A2(n_298),
.B1(n_299),
.B2(n_304),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_146),
.B(n_15),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_288),
.B(n_290),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_200),
.A2(n_174),
.B1(n_221),
.B2(n_208),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_203),
.B(n_186),
.Y(n_290)
);

BUFx12f_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_292),
.B(n_296),
.Y(n_363)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_207),
.B(n_187),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_172),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_295),
.Y(n_325)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_150),
.B(n_185),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_306),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_133),
.A2(n_153),
.B1(n_205),
.B2(n_226),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_137),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_300),
.B(n_301),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_190),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_203),
.B(n_227),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_164),
.B(n_161),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_303),
.B(n_170),
.C(n_250),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_214),
.A2(n_167),
.B1(n_166),
.B2(n_158),
.Y(n_304)
);

AO22x1_ASAP7_75t_L g305 ( 
.A1(n_175),
.A2(n_210),
.B1(n_183),
.B2(n_147),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_143),
.B(n_144),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_158),
.A2(n_166),
.B1(n_148),
.B2(n_144),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_147),
.B(n_183),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g365 ( 
.A1(n_308),
.A2(n_309),
.B(n_240),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_148),
.B(n_199),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_202),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_310),
.Y(n_346)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_199),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_311),
.B(n_315),
.Y(n_360)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_190),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_312),
.Y(n_347)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_194),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_313),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_194),
.B(n_162),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_209),
.B(n_168),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_316),
.B(n_317),
.Y(n_376)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_209),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_318),
.A2(n_265),
.B(n_306),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_273),
.A2(n_263),
.B1(n_303),
.B2(n_310),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_321),
.A2(n_343),
.B1(n_362),
.B2(n_259),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_323),
.B(n_305),
.Y(n_386)
);

AND2x2_ASAP7_75t_SL g334 ( 
.A(n_238),
.B(n_240),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g416 ( 
.A(n_334),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_254),
.B(n_250),
.C(n_276),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_355),
.C(n_364),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_260),
.A2(n_258),
.B1(n_289),
.B2(n_261),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_352),
.A2(n_375),
.B1(n_252),
.B2(n_317),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_276),
.B(n_249),
.C(n_253),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_297),
.A2(n_251),
.B1(n_244),
.B2(n_275),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_294),
.B(n_237),
.C(n_238),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_L g401 ( 
.A1(n_365),
.A2(n_379),
.B(n_255),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_268),
.A2(n_315),
.B1(n_316),
.B2(n_253),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_372),
.A2(n_313),
.B1(n_312),
.B2(n_300),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_292),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_291),
.A2(n_285),
.B1(n_314),
.B2(n_286),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_239),
.B(n_270),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_337),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_SL g394 ( 
.A1(n_378),
.A2(n_280),
.B(n_296),
.Y(n_394)
);

A2O1A1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_314),
.A2(n_237),
.B(n_277),
.C(n_291),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_265),
.B(n_234),
.C(n_267),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_281),
.C(n_247),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g381 ( 
.A(n_282),
.B(n_291),
.CI(n_305),
.CON(n_381),
.SN(n_381)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_381),
.B(n_323),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_382),
.A2(n_406),
.B1(n_410),
.B2(n_347),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_374),
.A2(n_291),
.B(n_235),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_384),
.A2(n_330),
.B(n_332),
.Y(n_459)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_336),
.Y(n_385)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_385),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_386),
.B(n_417),
.C(n_419),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_367),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_387),
.B(n_413),
.Y(n_465)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_389),
.B(n_394),
.Y(n_467)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_324),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_392),
.B(n_401),
.Y(n_468)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_393),
.Y(n_448)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_354),
.Y(n_395)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_395),
.Y(n_453)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_376),
.Y(n_396)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_396),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_397),
.B(n_404),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_345),
.B(n_311),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_399),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_241),
.Y(n_399)
);

OA21x2_ASAP7_75t_L g400 ( 
.A1(n_353),
.A2(n_375),
.B(n_379),
.Y(n_400)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_400),
.A2(n_361),
.B(n_332),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_352),
.A2(n_283),
.B1(n_271),
.B2(n_272),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_402),
.A2(n_346),
.B1(n_359),
.B2(n_347),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_349),
.A2(n_278),
.B1(n_246),
.B2(n_269),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_403),
.A2(n_414),
.B(n_423),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_335),
.B(n_348),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_341),
.Y(n_405)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_405),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_372),
.A2(n_256),
.B1(n_293),
.B2(n_274),
.Y(n_406)
);

INVx13_ASAP7_75t_L g407 ( 
.A(n_319),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_407),
.Y(n_439)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_411),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_SL g412 ( 
.A1(n_378),
.A2(n_266),
.B(n_267),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_428),
.B(n_339),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_319),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_327),
.B(n_242),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_421),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g417 ( 
.A(n_355),
.B(n_266),
.C(n_242),
.Y(n_417)
);

OAI21xp33_ASAP7_75t_L g418 ( 
.A1(n_338),
.A2(n_236),
.B(n_292),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_424),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_363),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_327),
.B(n_351),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_341),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_422),
.B(n_426),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_344),
.A2(n_331),
.B(n_371),
.Y(n_423)
);

NOR3xp33_ASAP7_75t_L g424 ( 
.A(n_335),
.B(n_377),
.C(n_358),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_322),
.B(n_320),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g436 ( 
.A(n_425),
.Y(n_436)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_427),
.B(n_429),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_319),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_431),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_351),
.B(n_337),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_440),
.A2(n_443),
.B1(n_446),
.B2(n_382),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_442),
.A2(n_451),
.B(n_456),
.Y(n_509)
);

OAI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_384),
.A2(n_381),
.B1(n_346),
.B2(n_328),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_389),
.A2(n_381),
.B1(n_334),
.B2(n_370),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_380),
.B(n_370),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_452),
.A2(n_471),
.B1(n_402),
.B2(n_390),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_364),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_454),
.B(n_455),
.C(n_462),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_383),
.B(n_334),
.C(n_370),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_400),
.A2(n_325),
.B(n_361),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_467),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_459),
.A2(n_464),
.B(n_429),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_357),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_414),
.A2(n_330),
.B(n_325),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_423),
.A2(n_366),
.B(n_359),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_466),
.A2(n_414),
.B(n_403),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_417),
.B(n_431),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_416),
.C(n_419),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_386),
.A2(n_368),
.B1(n_350),
.B2(n_369),
.Y(n_471)
);

AO22x2_ASAP7_75t_SL g474 ( 
.A1(n_446),
.A2(n_406),
.B1(n_409),
.B2(n_411),
.Y(n_474)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_474),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_449),
.B(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_475),
.Y(n_534)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_477),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_478),
.B(n_493),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_479),
.B(n_488),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_480),
.B(n_481),
.C(n_486),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_416),
.C(n_398),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_460),
.A2(n_408),
.B1(n_399),
.B2(n_415),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_482),
.A2(n_499),
.B1(n_511),
.B2(n_453),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_450),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_483),
.B(n_487),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_484),
.Y(n_527)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_465),
.Y(n_485)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_485),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_397),
.C(n_428),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_445),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_467),
.B(n_387),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_489),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_498),
.B1(n_513),
.B2(n_469),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_437),
.B(n_420),
.C(n_391),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_491),
.B(n_497),
.C(n_481),
.Y(n_540)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_492),
.Y(n_546)
);

A2O1A1Ixp33_ASAP7_75t_L g493 ( 
.A1(n_456),
.A2(n_388),
.B(n_393),
.C(n_395),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_444),
.B(n_385),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_494),
.B(n_506),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_495),
.A2(n_502),
.B(n_458),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_445),
.Y(n_496)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_496),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_437),
.B(n_470),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_444),
.A2(n_413),
.B1(n_422),
.B2(n_405),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_460),
.A2(n_427),
.B1(n_426),
.B2(n_430),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_500),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_451),
.B(n_366),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_462),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_459),
.A2(n_320),
.B(n_326),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_442),
.B(n_333),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_504),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_441),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_441),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_505),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_434),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_439),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_508),
.Y(n_537)
);

NOR2x1_ASAP7_75t_L g508 ( 
.A(n_473),
.B(n_333),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_464),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_434),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_463),
.A2(n_368),
.B1(n_350),
.B2(n_369),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_471),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_512),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_466),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g575 ( 
.A(n_514),
.B(n_551),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_490),
.A2(n_449),
.B1(n_463),
.B2(n_473),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_515),
.A2(n_547),
.B1(n_493),
.B2(n_532),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_435),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_516),
.B(n_518),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_476),
.B(n_433),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_489),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_519),
.B(n_523),
.Y(n_576)
);

AOI22x1_ASAP7_75t_L g520 ( 
.A1(n_488),
.A2(n_467),
.B1(n_440),
.B2(n_469),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_520),
.A2(n_502),
.B1(n_474),
.B2(n_506),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_489),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_524),
.A2(n_530),
.B(n_495),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_525),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_476),
.B(n_435),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_528),
.B(n_529),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_486),
.B(n_433),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_509),
.A2(n_458),
.B(n_468),
.Y(n_530)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_531),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_436),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_533),
.B(n_474),
.Y(n_581)
);

XNOR2x2_ASAP7_75t_SL g538 ( 
.A(n_475),
.B(n_501),
.Y(n_538)
);

AOI21xp33_ASAP7_75t_L g567 ( 
.A1(n_538),
.A2(n_474),
.B(n_494),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_540),
.B(n_485),
.C(n_509),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_488),
.A2(n_452),
.B1(n_453),
.B2(n_438),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_499),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_508),
.Y(n_559)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_550),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_491),
.B(n_448),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_552),
.B(n_581),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_477),
.C(n_482),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_554),
.B(n_555),
.C(n_565),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_484),
.C(n_510),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_541),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_557),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_559),
.B(n_561),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_560),
.A2(n_563),
.B(n_556),
.Y(n_606)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_541),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_563),
.A2(n_573),
.B1(n_580),
.B2(n_582),
.Y(n_600)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_531),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_564),
.B(n_566),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_535),
.B(n_528),
.C(n_516),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_546),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_567),
.B(n_530),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_518),
.B(n_505),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_571),
.C(n_583),
.Y(n_599)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_569),
.A2(n_439),
.B(n_407),
.C(n_373),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_R g571 ( 
.A(n_542),
.B(n_478),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_521),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_572),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_SL g573 ( 
.A1(n_527),
.A2(n_544),
.B1(n_536),
.B2(n_537),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_517),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_574),
.B(n_579),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_533),
.B(n_492),
.C(n_500),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_578),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_551),
.B(n_529),
.C(n_514),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_549),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_515),
.Y(n_580)
);

CKINVDCx14_ASAP7_75t_R g582 ( 
.A(n_526),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_526),
.B(n_438),
.Y(n_583)
);

XNOR2x1_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_555),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_576),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_586),
.B(n_596),
.Y(n_624)
);

FAx1_ASAP7_75t_SL g587 ( 
.A(n_552),
.B(n_538),
.CI(n_534),
.CON(n_587),
.SN(n_587)
);

XOR2x1_ASAP7_75t_L g626 ( 
.A(n_587),
.B(n_597),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_558),
.B(n_527),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_605),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_560),
.A2(n_522),
.B(n_539),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g611 ( 
.A1(n_590),
.A2(n_606),
.B(n_609),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_577),
.B(n_539),
.Y(n_591)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_591),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_553),
.A2(n_532),
.B1(n_543),
.B2(n_534),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_593),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_553),
.A2(n_543),
.B1(n_547),
.B2(n_550),
.Y(n_594)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_594),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_564),
.A2(n_543),
.B1(n_524),
.B2(n_520),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_556),
.A2(n_520),
.B(n_506),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_580),
.A2(n_545),
.B1(n_511),
.B2(n_448),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_598),
.B(n_557),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_562),
.A2(n_545),
.B1(n_447),
.B2(n_461),
.Y(n_603)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_603),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_558),
.B(n_447),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_554),
.B(n_461),
.Y(n_607)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_607),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_565),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_613),
.B(n_615),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_595),
.B(n_570),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_621),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_570),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g618 ( 
.A(n_585),
.B(n_581),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_618),
.B(n_630),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g640 ( 
.A(n_619),
.B(n_584),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_595),
.B(n_579),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_608),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_622),
.B(n_625),
.Y(n_637)
);

CKINVDCx16_ASAP7_75t_R g625 ( 
.A(n_595),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_578),
.C(n_575),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_627),
.B(n_629),
.Y(n_639)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_628),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_601),
.B(n_575),
.C(n_561),
.Y(n_629)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_605),
.B(n_574),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_624),
.A2(n_600),
.B1(n_590),
.B2(n_599),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_633),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_613),
.B(n_588),
.C(n_606),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_612),
.B(n_586),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_634),
.B(n_643),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g658 ( 
.A(n_640),
.B(n_647),
.Y(n_658)
);

OAI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_624),
.A2(n_592),
.B(n_587),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_641),
.A2(n_611),
.B(n_619),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_623),
.B(n_592),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_642),
.B(n_646),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_618),
.B(n_629),
.C(n_615),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g644 ( 
.A1(n_616),
.A2(n_597),
.B1(n_602),
.B2(n_593),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_644),
.B(n_645),
.Y(n_661)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_630),
.B(n_602),
.C(n_594),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_620),
.B(n_608),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g647 ( 
.A(n_610),
.B(n_596),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_617),
.B(n_598),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_648),
.B(n_611),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_649),
.B(n_653),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_633),
.B(n_620),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_650),
.B(n_657),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_SL g655 ( 
.A1(n_638),
.A2(n_626),
.B(n_628),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_655),
.B(n_656),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_639),
.B(n_627),
.C(n_626),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_631),
.B(n_604),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_632),
.A2(n_610),
.B(n_587),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_659),
.B(n_640),
.C(n_643),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_647),
.B(n_604),
.Y(n_660)
);

XNOR2xp5_ASAP7_75t_L g668 ( 
.A(n_660),
.B(n_662),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_645),
.A2(n_566),
.B(n_609),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_SL g663 ( 
.A1(n_651),
.A2(n_637),
.B(n_636),
.Y(n_663)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_663),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_665),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_654),
.B(n_635),
.C(n_636),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_666),
.B(n_667),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g667 ( 
.A(n_652),
.B(n_635),
.C(n_644),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_661),
.B(n_326),
.Y(n_669)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_669),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_660),
.B(n_369),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_SL g678 ( 
.A1(n_672),
.A2(n_658),
.B(n_356),
.C(n_373),
.Y(n_678)
);

A2O1A1O1Ixp25_ASAP7_75t_L g673 ( 
.A1(n_671),
.A2(n_655),
.B(n_658),
.C(n_662),
.D(n_329),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_673),
.B(n_678),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_675),
.Y(n_679)
);

AO21x1_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_664),
.B(n_668),
.Y(n_682)
);

A2O1A1Ixp33_ASAP7_75t_SL g681 ( 
.A1(n_676),
.A2(n_670),
.B(n_677),
.C(n_664),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_681),
.Y(n_683)
);

NOR3xp33_ASAP7_75t_L g684 ( 
.A(n_682),
.B(n_680),
.C(n_674),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_684),
.B(n_683),
.Y(n_685)
);

HAxp5_ASAP7_75t_SL g686 ( 
.A(n_685),
.B(n_329),
.CON(n_686),
.SN(n_686)
);


endmodule