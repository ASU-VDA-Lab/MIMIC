module fake_jpeg_20430_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_69),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_81),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_51),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_58),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_52),
.B1(n_40),
.B2(n_53),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_95),
.B1(n_41),
.B2(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_60),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_90),
.A2(n_92),
.B(n_56),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_46),
.B(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_42),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_96),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_61),
.B1(n_47),
.B2(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_103),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_84),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_1),
.C(n_2),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_105),
.B(n_1),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_45),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_64),
.B1(n_57),
.B2(n_50),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_110),
.B(n_21),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_85),
.A2(n_20),
.B1(n_37),
.B2(n_35),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_16),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_113),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_19),
.C(n_33),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_118),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_117),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_2),
.Y(n_118)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_108),
.B1(n_109),
.B2(n_8),
.Y(n_123)
);

XNOR2x2_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_38),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_23),
.B(n_32),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_125),
.A2(n_111),
.B1(n_124),
.B2(n_122),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_121),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_128),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_126),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_123),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_133),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_115),
.B(n_14),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_11),
.Y(n_137)
);


endmodule