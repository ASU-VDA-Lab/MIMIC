module fake_jpeg_16035_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_240;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_39),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_20),
.Y(n_43)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_44),
.C(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_20),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_31),
.B(n_2),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_25),
.C(n_22),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_17),
.B1(n_18),
.B2(n_26),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_18),
.B1(n_37),
.B2(n_27),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_34),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_62),
.B(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_35),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_18),
.B1(n_17),
.B2(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_64),
.A2(n_85),
.B1(n_52),
.B2(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_70),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_35),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_23),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_24),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

OR2x4_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_30),
.Y(n_79)
);

NOR2xp67_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_30),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_34),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_84),
.Y(n_115)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_87),
.Y(n_110)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

OAI22x1_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_40),
.B1(n_36),
.B2(n_30),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_102),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_47),
.C(n_40),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_97),
.C(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_58),
.A2(n_52),
.B1(n_40),
.B2(n_36),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_105),
.B1(n_82),
.B2(n_57),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_27),
.B1(n_19),
.B2(n_22),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_86),
.A2(n_40),
.B1(n_36),
.B2(n_47),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_86),
.B1(n_74),
.B2(n_68),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_25),
.B1(n_60),
.B2(n_21),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_70),
.B(n_67),
.C(n_75),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_111),
.B1(n_107),
.B2(n_108),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_90),
.Y(n_118)
);

INVxp33_ASAP7_75t_SL g162 ( 
.A(n_118),
.Y(n_162)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_91),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_126),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_108),
.B(n_112),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_132),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_94),
.A2(n_69),
.A3(n_71),
.B1(n_25),
.B2(n_32),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_139),
.C(n_99),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_135),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_83),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_72),
.C(n_56),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_93),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_104),
.B(n_21),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_140),
.A2(n_111),
.B(n_92),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_143),
.A2(n_154),
.B(n_167),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_149),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_4),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_111),
.B(n_101),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_133),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_107),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_158),
.B(n_1),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_111),
.C(n_105),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_147),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_168),
.B1(n_31),
.B2(n_4),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_104),
.B1(n_110),
.B2(n_56),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_120),
.B(n_129),
.C(n_122),
.D(n_131),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_124),
.A3(n_136),
.B1(n_132),
.B2(n_130),
.C1(n_139),
.C2(n_116),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_170),
.B(n_172),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_166),
.B(n_98),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_193),
.C(n_151),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_103),
.B(n_110),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_103),
.B(n_32),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_16),
.B(n_73),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_142),
.B(n_163),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_180),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_88),
.B1(n_16),
.B2(n_90),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_181),
.A2(n_184),
.B1(n_187),
.B2(n_155),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_186),
.Y(n_198)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_153),
.A2(n_31),
.B1(n_14),
.B2(n_3),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_1),
.B(n_2),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_167),
.A2(n_31),
.B(n_3),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_4),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_203),
.C(n_193),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_186),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_177),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_202),
.B(n_204),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_153),
.C(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_210),
.A2(n_176),
.B1(n_188),
.B2(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_185),
.B1(n_179),
.B2(n_187),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_215),
.A2(n_224),
.B1(n_226),
.B2(n_208),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_227),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_209),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_220),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_178),
.C(n_188),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_184),
.C(n_200),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_195),
.A2(n_165),
.B(n_192),
.Y(n_223)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_223),
.A2(n_205),
.B(n_207),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_196),
.A2(n_156),
.B1(n_152),
.B2(n_148),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_198),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_148),
.B1(n_156),
.B2(n_149),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_191),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_199),
.B1(n_207),
.B2(n_197),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_230),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_231),
.B(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_211),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_227),
.B(n_164),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_5),
.C(n_6),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_7),
.Y(n_241)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_226),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_239),
.B1(n_244),
.B2(n_221),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_242),
.A2(n_243),
.B(n_245),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_232),
.A2(n_217),
.B(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_212),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_223),
.B(n_220),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_228),
.B(n_237),
.Y(n_251)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_249),
.A2(n_250),
.B(n_10),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_212),
.B(n_234),
.Y(n_250)
);

AO21x1_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_11),
.B(n_12),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_7),
.C(n_8),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_255),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_256),
.Y(n_258)
);

AOI31xp33_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_10),
.A3(n_11),
.B(n_12),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_248),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_259),
.C(n_258),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_13),
.Y(n_262)
);


endmodule