module real_jpeg_208_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_1),
.A2(n_27),
.B1(n_39),
.B2(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_42),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_38),
.B1(n_57),
.B2(n_59),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_56),
.C(n_57),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_38),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_38),
.B1(n_61),
.B2(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_2),
.B(n_54),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_39),
.C(n_71),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_2),
.B(n_24),
.C(n_46),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_69),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_2),
.B(n_30),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_180),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_4),
.A2(n_39),
.B1(n_42),
.B2(n_62),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_62),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_9),
.A2(n_34),
.B1(n_39),
.B2(n_42),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_34),
.B1(n_61),
.B2(n_63),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_9),
.A2(n_34),
.B1(n_57),
.B2(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_132),
.B1(n_251),
.B2(n_252),
.Y(n_13)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_131),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_106),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_17),
.B(n_106),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.C(n_97),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_18),
.A2(n_19),
.B1(n_97),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_51),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_20),
.B(n_68),
.C(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_35),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_21),
.B(n_35),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_28),
.B(n_31),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_22),
.A2(n_29),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_24),
.B(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_28),
.B(n_33),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_28),
.A2(n_29),
.B(n_105),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_28),
.B(n_105),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_28),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_29),
.B(n_209),
.Y(n_223)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_30),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_31),
.B(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_32),
.B(n_208),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_49),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_36),
.B(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.Y(n_36)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_37),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_37),
.B(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_42),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_39),
.B(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_43),
.B(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_43),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_43),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_48),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_49),
.A2(n_100),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_49),
.B(n_181),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_68),
.B1(n_77),
.B2(n_78),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_53),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_54),
.B(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_56),
.B1(n_61),
.B2(n_63),
.Y(n_66)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_59),
.B1(n_71),
.B2(n_72),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_57),
.B(n_176),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_73),
.B(n_76),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_69),
.B(n_90),
.Y(n_150)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_73),
.B(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_74),
.B(n_121),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_79),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_91),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_96),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_97),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_102),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

AOI21x1_ASAP7_75t_SL g145 ( 
.A1(n_99),
.A2(n_129),
.B(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_99),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_101),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_103),
.B(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_124),
.B2(n_125),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_123),
.B(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_126),
.A2(n_127),
.B1(n_174),
.B2(n_175),
.Y(n_196)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_132),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_242),
.B(n_248),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_166),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_152),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_135),
.B(n_152),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_136),
.B(n_139),
.C(n_151),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_151),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_147),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_159),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_154),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_159),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_165),
.B(n_223),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_186),
.B(n_241),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_183),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_168),
.B(n_183),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.C(n_177),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_170),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_173),
.A2(n_177),
.B1(n_178),
.B2(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_180),
.B(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI21x1_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_197),
.B(n_240),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_192),
.Y(n_240)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_196),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_195),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_235),
.B(n_239),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_217),
.B(n_234),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_210),
.B1(n_211),
.B2(n_216),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_206),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_212),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_224),
.B(n_233),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_221),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_229),
.B(n_232),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_247),
.Y(n_250)
);


endmodule