module real_jpeg_20936_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_215;
wire n_221;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_200;
wire n_48;
wire n_56;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_0),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_0),
.A2(n_28),
.B1(n_49),
.B2(n_50),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_0),
.A2(n_28),
.B1(n_64),
.B2(n_65),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_79),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_1),
.A2(n_64),
.B1(n_65),
.B2(n_79),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_4),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_43),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_5),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_198)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_7),
.B(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_7),
.A2(n_184),
.B(n_208),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_9),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_11),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_11),
.A2(n_49),
.B1(n_50),
.B2(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_12),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_30),
.B(n_33),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_60),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_12),
.B(n_98),
.Y(n_138)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_12),
.A2(n_50),
.B(n_81),
.C(n_151),
.D(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_50),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_12),
.B(n_48),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_67),
.B(n_166),
.Y(n_186)
);

A2O1A1O1Ixp25_ASAP7_75t_L g199 ( 
.A1(n_12),
.A2(n_32),
.B(n_45),
.C(n_53),
.D(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_12),
.B(n_32),
.Y(n_200)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_102),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_21),
.B(n_102),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.C(n_88),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_22),
.B(n_143),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_24),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_25),
.A2(n_29),
.B1(n_38),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_29),
.B(n_31),
.C(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_31),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_27),
.A2(n_31),
.B(n_60),
.C(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_35),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_37),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_40),
.B(n_56),
.C(n_57),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B(n_52),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_42),
.A2(n_44),
.B1(n_55),
.B2(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_45),
.B(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_47),
.Y(n_206)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_82),
.B(n_83),
.C(n_84),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_82),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_49),
.B(n_51),
.Y(n_205)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_50),
.A2(n_200),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_55),
.A2(n_101),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_60),
.B(n_87),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_60),
.B(n_107),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_62),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_63),
.A2(n_67),
.B1(n_107),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_65),
.B1(n_82),
.B2(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_64),
.B(n_82),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_64),
.B(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_65),
.A2(n_83),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_69),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_75),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_67),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_67),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_67),
.B(n_168),
.Y(n_184)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_68),
.A2(n_173),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_71),
.B(n_88),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_77),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_77),
.Y(n_113)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_87),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_80),
.A2(n_86),
.B1(n_87),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_80),
.A2(n_87),
.B1(n_163),
.B2(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_80),
.A2(n_198),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_92),
.Y(n_91)
);

CKINVDCx9p33_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_87),
.B(n_93),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_87),
.A2(n_91),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.C(n_99),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_90),
.B1(n_99),
.B2(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_124),
.B2(n_125),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_112),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_107),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_124),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_144),
.B(n_229),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_129),
.B(n_142),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_130),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_132),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_139),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_136),
.A2(n_137),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_138),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_223),
.B(n_228),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_211),
.B(n_222),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_192),
.B(n_210),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_169),
.B(n_191),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_149),
.B(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_153),
.B1(n_154),
.B2(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_164),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_179),
.B(n_190),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_171),
.B(n_177),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_185),
.B(n_189),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_182),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_194),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_203),
.B2(n_209),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_202),
.C(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_207),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_218),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_219),
.C(n_220),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_215),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_225),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);


endmodule