module real_aes_8954_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_705, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_705;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_691;
wire n_498;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g166 ( .A1(n_0), .A2(n_167), .B(n_168), .C(n_172), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_1), .B(n_161), .Y(n_174) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_3), .B(n_146), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_4), .A2(n_135), .B(n_152), .C(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_5), .A2(n_155), .B(n_479), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_6), .A2(n_155), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_7), .B(n_161), .Y(n_485) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_8), .A2(n_127), .B(n_214), .Y(n_213) );
AND2x6_ASAP7_75t_L g152 ( .A(n_9), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_10), .A2(n_135), .B(n_152), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g450 ( .A(n_11), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_12), .B(n_40), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_12), .B(n_40), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_13), .B(n_171), .Y(n_460) );
INVx1_ASAP7_75t_L g132 ( .A(n_14), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_15), .B(n_146), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_16), .A2(n_147), .B(n_469), .C(n_471), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_17), .B(n_161), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g117 ( .A1(n_18), .A2(n_64), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_18), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_19), .B(n_204), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_20), .A2(n_135), .B(n_198), .C(n_203), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_21), .A2(n_170), .B(n_222), .C(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_22), .B(n_171), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_23), .B(n_171), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_24), .Y(n_488) );
INVx1_ASAP7_75t_L g500 ( .A(n_25), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_26), .A2(n_135), .B(n_203), .C(n_217), .Y(n_216) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_27), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_28), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_29), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g517 ( .A(n_30), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_31), .A2(n_155), .B(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g137 ( .A(n_32), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_33), .A2(n_150), .B(n_182), .C(n_183), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_34), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_35), .A2(n_170), .B(n_482), .C(n_484), .Y(n_481) );
INVxp67_ASAP7_75t_L g518 ( .A(n_36), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_37), .B(n_219), .Y(n_218) );
CKINVDCx14_ASAP7_75t_R g480 ( .A(n_38), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_39), .A2(n_135), .B(n_203), .C(n_499), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_41), .A2(n_172), .B(n_448), .C(n_449), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_42), .B(n_196), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_43), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_44), .B(n_146), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_45), .B(n_155), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_46), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_47), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_48), .A2(n_150), .B(n_182), .C(n_243), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_49), .A2(n_421), .B1(n_690), .B2(n_691), .C1(n_694), .C2(n_697), .Y(n_420) );
INVx1_ASAP7_75t_L g169 ( .A(n_50), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_51), .A2(n_82), .B1(n_692), .B2(n_693), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_51), .Y(n_693) );
INVx1_ASAP7_75t_L g244 ( .A(n_52), .Y(n_244) );
INVx1_ASAP7_75t_L g438 ( .A(n_53), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_54), .B(n_155), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_55), .Y(n_207) );
CKINVDCx14_ASAP7_75t_R g446 ( .A(n_56), .Y(n_446) );
INVx1_ASAP7_75t_L g153 ( .A(n_57), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_58), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_59), .B(n_161), .Y(n_262) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_60), .A2(n_142), .B(n_202), .C(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g131 ( .A(n_61), .Y(n_131) );
INVx1_ASAP7_75t_SL g483 ( .A(n_62), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_63), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_64), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_65), .B(n_146), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_66), .B(n_161), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_67), .B(n_147), .Y(n_233) );
INVx1_ASAP7_75t_L g491 ( .A(n_68), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g164 ( .A(n_69), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_70), .B(n_186), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g134 ( .A1(n_71), .A2(n_135), .B(n_140), .C(n_150), .Y(n_134) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_72), .Y(n_258) );
INVx1_ASAP7_75t_L g109 ( .A(n_73), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_74), .A2(n_102), .B1(n_110), .B2(n_703), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_75), .A2(n_155), .B(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_76), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_77), .A2(n_155), .B(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_78), .A2(n_196), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g467 ( .A(n_79), .Y(n_467) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_80), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_81), .B(n_185), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_82), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_83), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_84), .A2(n_155), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g470 ( .A(n_85), .Y(n_470) );
INVx2_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g459 ( .A(n_87), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_88), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_89), .B(n_171), .Y(n_234) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_90), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g413 ( .A(n_90), .B(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g424 ( .A(n_90), .B(n_415), .Y(n_424) );
INVx2_ASAP7_75t_L g428 ( .A(n_90), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_91), .A2(n_135), .B(n_150), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_92), .B(n_155), .Y(n_180) );
INVx1_ASAP7_75t_L g184 ( .A(n_93), .Y(n_184) );
INVxp67_ASAP7_75t_L g261 ( .A(n_94), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_95), .B(n_127), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_96), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g141 ( .A(n_97), .Y(n_141) );
INVx1_ASAP7_75t_L g229 ( .A(n_98), .Y(n_229) );
INVx2_ASAP7_75t_L g441 ( .A(n_99), .Y(n_441) );
AND2x2_ASAP7_75t_L g246 ( .A(n_100), .B(n_189), .Y(n_246) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g703 ( .A(n_103), .Y(n_703) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g415 ( .A(n_106), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AO21x2_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_419), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g702 ( .A(n_114), .Y(n_702) );
OAI21xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_411), .B(n_417), .Y(n_115) );
XNOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx2_ASAP7_75t_L g425 ( .A(n_120), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_120), .A2(n_423), .B1(n_699), .B2(n_700), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g120 ( .A(n_121), .B(n_354), .Y(n_120) );
AND4x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_294), .C(n_309), .D(n_334), .Y(n_121) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_267), .Y(n_122) );
OAI21xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_175), .B(n_247), .Y(n_123) );
AND2x2_ASAP7_75t_L g297 ( .A(n_124), .B(n_193), .Y(n_297) );
AND2x2_ASAP7_75t_L g310 ( .A(n_124), .B(n_192), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_124), .B(n_176), .Y(n_360) );
INVx1_ASAP7_75t_L g364 ( .A(n_124), .Y(n_364) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
INVx2_ASAP7_75t_L g281 ( .A(n_125), .Y(n_281) );
BUFx2_ASAP7_75t_L g308 ( .A(n_125), .Y(n_308) );
AO21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_133), .B(n_158), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_126), .B(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g161 ( .A(n_126), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_126), .B(n_191), .Y(n_190) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_126), .A2(n_228), .B(n_235), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_126), .B(n_463), .Y(n_462) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_126), .A2(n_487), .B(n_493), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_126), .B(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_127), .A2(n_215), .B(n_216), .Y(n_214) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_127), .Y(n_255) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g237 ( .A(n_128), .Y(n_237) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
AND2x2_ASAP7_75t_SL g189 ( .A(n_129), .B(n_130), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_154), .Y(n_133) );
INVx5_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
AND2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
BUFx3_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
INVx1_ASAP7_75t_L g223 ( .A(n_137), .Y(n_223) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_139), .Y(n_144) );
INVx3_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
AND2x2_ASAP7_75t_L g156 ( .A(n_139), .B(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
INVx1_ASAP7_75t_L g219 ( .A(n_139), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_145), .C(n_148), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_143), .B(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_143), .B(n_470), .Y(n_469) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_143), .A2(n_146), .B1(n_517), .B2(n_518), .Y(n_516) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g186 ( .A(n_144), .Y(n_186) );
INVx2_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_146), .B(n_261), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_146), .A2(n_201), .B(n_500), .C(n_501), .Y(n_499) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_147), .B(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx3_ASAP7_75t_L g484 ( .A(n_149), .Y(n_484) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
O2A1O1Ixp33_ASAP7_75t_SL g163 ( .A1(n_151), .A2(n_164), .B(n_165), .C(n_166), .Y(n_163) );
O2A1O1Ixp33_ASAP7_75t_L g257 ( .A1(n_151), .A2(n_165), .B(n_258), .C(n_259), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_SL g437 ( .A1(n_151), .A2(n_165), .B(n_438), .C(n_439), .Y(n_437) );
O2A1O1Ixp33_ASAP7_75t_SL g445 ( .A1(n_151), .A2(n_165), .B(n_446), .C(n_447), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_SL g466 ( .A1(n_151), .A2(n_165), .B(n_467), .C(n_468), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_151), .A2(n_165), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_151), .A2(n_165), .B(n_514), .C(n_515), .Y(n_513) );
INVx4_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g155 ( .A(n_152), .B(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_152), .B(n_156), .Y(n_230) );
BUFx2_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx1_ASAP7_75t_L g202 ( .A(n_157), .Y(n_202) );
AND2x2_ASAP7_75t_L g248 ( .A(n_160), .B(n_193), .Y(n_248) );
INVx2_ASAP7_75t_L g264 ( .A(n_160), .Y(n_264) );
AND2x2_ASAP7_75t_L g273 ( .A(n_160), .B(n_192), .Y(n_273) );
AND2x2_ASAP7_75t_L g352 ( .A(n_160), .B(n_281), .Y(n_352) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_174), .Y(n_160) );
INVx2_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_170), .B(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g448 ( .A(n_171), .Y(n_448) );
INVx2_ASAP7_75t_L g461 ( .A(n_172), .Y(n_461) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_173), .Y(n_188) );
INVx1_ASAP7_75t_L g471 ( .A(n_173), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_209), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_176), .B(n_279), .Y(n_317) );
INVx1_ASAP7_75t_L g405 ( .A(n_176), .Y(n_405) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_192), .Y(n_176) );
AND2x2_ASAP7_75t_L g263 ( .A(n_177), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g277 ( .A(n_177), .B(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_177), .Y(n_306) );
OR2x2_ASAP7_75t_L g338 ( .A(n_177), .B(n_280), .Y(n_338) );
AND2x2_ASAP7_75t_L g346 ( .A(n_177), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g379 ( .A(n_177), .B(n_348), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_177), .B(n_248), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_177), .B(n_308), .Y(n_404) );
AND2x2_ASAP7_75t_L g410 ( .A(n_177), .B(n_297), .Y(n_410) );
INVx5_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx2_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
AND2x2_ASAP7_75t_L g300 ( .A(n_178), .B(n_280), .Y(n_300) );
AND2x2_ASAP7_75t_L g333 ( .A(n_178), .B(n_293), .Y(n_333) );
AND2x2_ASAP7_75t_L g353 ( .A(n_178), .B(n_193), .Y(n_353) );
AND2x2_ASAP7_75t_L g387 ( .A(n_178), .B(n_253), .Y(n_387) );
OR2x6_ASAP7_75t_L g178 ( .A(n_179), .B(n_190), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_189), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_187), .C(n_188), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_185), .A2(n_188), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_185), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_185), .A2(n_461), .B(n_491), .C(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
INVx1_ASAP7_75t_L g208 ( .A(n_189), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_189), .A2(n_241), .B(n_242), .Y(n_240) );
OA21x2_ASAP7_75t_L g443 ( .A1(n_189), .A2(n_444), .B(n_451), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_189), .A2(n_230), .B(n_497), .C(n_498), .Y(n_496) );
AND2x4_ASAP7_75t_L g293 ( .A(n_192), .B(n_264), .Y(n_293) );
AND2x2_ASAP7_75t_L g304 ( .A(n_192), .B(n_300), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_192), .B(n_280), .Y(n_343) );
INVx2_ASAP7_75t_L g358 ( .A(n_192), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_192), .B(n_292), .Y(n_381) );
AND2x2_ASAP7_75t_L g400 ( .A(n_192), .B(n_352), .Y(n_400) );
INVx5_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_193), .Y(n_299) );
AND2x2_ASAP7_75t_L g307 ( .A(n_193), .B(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g348 ( .A(n_193), .B(n_264), .Y(n_348) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_206), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g194 ( .A1(n_195), .A2(n_197), .B(n_204), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .Y(n_198) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_202), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_205), .B(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_208), .A2(n_455), .B(n_462), .Y(n_454) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_224), .Y(n_210) );
AND2x2_ASAP7_75t_L g271 ( .A(n_211), .B(n_254), .Y(n_271) );
INVx1_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_212), .B(n_227), .Y(n_251) );
OR2x2_ASAP7_75t_L g284 ( .A(n_212), .B(n_254), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_212), .B(n_254), .Y(n_289) );
AND2x2_ASAP7_75t_L g316 ( .A(n_212), .B(n_253), .Y(n_316) );
AND2x2_ASAP7_75t_L g368 ( .A(n_212), .B(n_226), .Y(n_368) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_213), .B(n_238), .Y(n_276) );
AND2x2_ASAP7_75t_L g312 ( .A(n_213), .B(n_227), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_220), .B(n_221), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_221), .A2(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_224), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g302 ( .A(n_225), .B(n_284), .Y(n_302) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_238), .Y(n_225) );
OAI322xp33_ASAP7_75t_L g267 ( .A1(n_226), .A2(n_268), .A3(n_272), .B1(n_274), .B2(n_277), .C1(n_282), .C2(n_290), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_226), .B(n_253), .Y(n_275) );
OR2x2_ASAP7_75t_L g285 ( .A(n_226), .B(n_239), .Y(n_285) );
AND2x2_ASAP7_75t_L g287 ( .A(n_226), .B(n_239), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_226), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_226), .B(n_254), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_226), .B(n_383), .Y(n_382) );
INVx5_ASAP7_75t_SL g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_227), .B(n_271), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_231), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_230), .A2(n_456), .B(n_457), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_230), .A2(n_488), .B(n_489), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g511 ( .A(n_237), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_238), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g265 ( .A(n_238), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_238), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g327 ( .A(n_238), .B(n_254), .Y(n_327) );
AOI211xp5_ASAP7_75t_SL g355 ( .A1(n_238), .A2(n_356), .B(n_359), .C(n_371), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_238), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g393 ( .A(n_238), .B(n_368), .Y(n_393) );
INVx5_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g321 ( .A(n_239), .B(n_254), .Y(n_321) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_239), .Y(n_330) );
AND2x2_ASAP7_75t_L g370 ( .A(n_239), .B(n_368), .Y(n_370) );
AND2x2_ASAP7_75t_SL g401 ( .A(n_239), .B(n_271), .Y(n_401) );
AND2x2_ASAP7_75t_L g408 ( .A(n_239), .B(n_367), .Y(n_408) );
OR2x6_ASAP7_75t_L g239 ( .A(n_240), .B(n_246), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B1(n_263), .B2(n_265), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_248), .B(n_270), .Y(n_318) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g266 ( .A(n_251), .Y(n_266) );
OR2x2_ASAP7_75t_L g326 ( .A(n_251), .B(n_327), .Y(n_326) );
OAI221xp5_ASAP7_75t_SL g374 ( .A1(n_251), .A2(n_375), .B1(n_377), .B2(n_378), .C(n_380), .Y(n_374) );
INVx2_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
AND2x2_ASAP7_75t_L g286 ( .A(n_253), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g376 ( .A(n_253), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_253), .B(n_368), .Y(n_389) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVxp67_ASAP7_75t_L g331 ( .A(n_254), .Y(n_331) );
AND2x2_ASAP7_75t_L g367 ( .A(n_254), .B(n_368), .Y(n_367) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_262), .Y(n_254) );
OA21x2_ASAP7_75t_L g435 ( .A1(n_255), .A2(n_436), .B(n_442), .Y(n_435) );
OA21x2_ASAP7_75t_L g464 ( .A1(n_255), .A2(n_465), .B(n_472), .Y(n_464) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_255), .A2(n_478), .B(n_485), .Y(n_477) );
AND2x2_ASAP7_75t_L g369 ( .A(n_263), .B(n_308), .Y(n_369) );
AND2x2_ASAP7_75t_L g279 ( .A(n_264), .B(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_264), .B(n_337), .Y(n_336) );
NOR2xp33_ASAP7_75t_SL g350 ( .A(n_266), .B(n_313), .Y(n_350) );
INVx1_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g356 ( .A(n_269), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
OR2x2_ASAP7_75t_L g342 ( .A(n_270), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g407 ( .A(n_270), .B(n_352), .Y(n_407) );
INVx2_ASAP7_75t_L g340 ( .A(n_271), .Y(n_340) );
NAND4xp25_ASAP7_75t_SL g403 ( .A(n_272), .B(n_404), .C(n_405), .D(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_273), .B(n_337), .Y(n_372) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_SL g409 ( .A(n_276), .Y(n_409) );
O2A1O1Ixp33_ASAP7_75t_SL g371 ( .A1(n_277), .A2(n_340), .B(n_344), .C(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g366 ( .A(n_279), .B(n_358), .Y(n_366) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_280), .Y(n_292) );
INVx1_ASAP7_75t_L g347 ( .A(n_280), .Y(n_347) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_281), .Y(n_324) );
AOI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B(n_286), .C(n_288), .Y(n_282) );
AND2x2_ASAP7_75t_L g303 ( .A(n_283), .B(n_287), .Y(n_303) );
OAI322xp33_ASAP7_75t_SL g341 ( .A1(n_283), .A2(n_342), .A3(n_344), .B1(n_345), .B2(n_349), .C1(n_350), .C2(n_351), .Y(n_341) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g363 ( .A(n_285), .B(n_289), .Y(n_363) );
INVx1_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
INVx1_ASAP7_75t_SL g362 ( .A(n_289), .Y(n_362) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI222xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_301), .B1(n_303), .B2(n_304), .C1(n_305), .C2(n_705), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_296), .B(n_298), .Y(n_295) );
OAI322xp33_ASAP7_75t_L g384 ( .A1(n_296), .A2(n_358), .A3(n_363), .B1(n_385), .B2(n_386), .C1(n_388), .C2(n_389), .Y(n_384) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_297), .A2(n_311), .B1(n_335), .B2(n_339), .C(n_341), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
OAI222xp33_ASAP7_75t_L g314 ( .A1(n_302), .A2(n_315), .B1(n_317), .B2(n_318), .C1(n_319), .C2(n_322), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_304), .A2(n_311), .B1(n_381), .B2(n_382), .Y(n_380) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
AOI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_314), .C(n_325), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g390 ( .A1(n_311), .A2(n_348), .B(n_391), .C(n_394), .Y(n_390) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x2_ASAP7_75t_L g320 ( .A(n_312), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g383 ( .A(n_316), .Y(n_383) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_323), .B(n_348), .Y(n_377) );
BUFx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B(n_332), .Y(n_325) );
OAI221xp5_ASAP7_75t_SL g394 ( .A1(n_326), .A2(n_395), .B1(n_396), .B2(n_397), .C(n_398), .Y(n_394) );
INVxp33_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_337), .B(n_348), .Y(n_388) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g399 ( .A(n_352), .B(n_358), .Y(n_399) );
AND4x1_ASAP7_75t_L g354 ( .A(n_355), .B(n_373), .C(n_390), .D(n_402), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_361), .B1(n_363), .B2(n_364), .C(n_365), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_369), .B2(n_370), .Y(n_365) );
INVx1_ASAP7_75t_L g395 ( .A(n_366), .Y(n_395) );
INVx1_ASAP7_75t_SL g385 ( .A(n_370), .Y(n_385) );
NOR2xp33_ASAP7_75t_SL g373 ( .A(n_374), .B(n_384), .Y(n_373) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_386), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_393), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g418 ( .A(n_413), .Y(n_418) );
NOR2x2_ASAP7_75t_L g696 ( .A(n_414), .B(n_428), .Y(n_696) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g427 ( .A(n_415), .B(n_428), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_417), .A2(n_420), .B(n_701), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B1(n_426), .B2(n_429), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx6_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g699 ( .A(n_427), .Y(n_699) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g700 ( .A(n_430), .Y(n_700) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_616), .Y(n_430) );
NOR4xp25_ASAP7_75t_L g431 ( .A(n_432), .B(n_558), .C(n_588), .D(n_598), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_473), .B(n_521), .C(n_548), .Y(n_432) );
OAI222xp33_ASAP7_75t_L g643 ( .A1(n_433), .A2(n_563), .B1(n_644), .B2(n_645), .C1(n_646), .C2(n_647), .Y(n_643) );
OR2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_452), .Y(n_433) );
AOI33xp33_ASAP7_75t_L g569 ( .A1(n_434), .A2(n_556), .A3(n_557), .B1(n_570), .B2(n_575), .B3(n_577), .Y(n_569) );
OAI211xp5_ASAP7_75t_SL g626 ( .A1(n_434), .A2(n_627), .B(n_629), .C(n_631), .Y(n_626) );
OR2x2_ASAP7_75t_L g642 ( .A(n_434), .B(n_628), .Y(n_642) );
INVx1_ASAP7_75t_L g675 ( .A(n_434), .Y(n_675) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_443), .Y(n_434) );
INVx2_ASAP7_75t_L g552 ( .A(n_435), .Y(n_552) );
AND2x2_ASAP7_75t_L g568 ( .A(n_435), .B(n_464), .Y(n_568) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_435), .Y(n_603) );
AND2x2_ASAP7_75t_L g632 ( .A(n_435), .B(n_443), .Y(n_632) );
INVx2_ASAP7_75t_L g532 ( .A(n_443), .Y(n_532) );
BUFx3_ASAP7_75t_L g540 ( .A(n_443), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_443), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g551 ( .A(n_443), .B(n_552), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_443), .B(n_453), .Y(n_580) );
AND2x2_ASAP7_75t_L g649 ( .A(n_443), .B(n_583), .Y(n_649) );
INVx2_ASAP7_75t_SL g543 ( .A(n_452), .Y(n_543) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_464), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_453), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g585 ( .A(n_453), .Y(n_585) );
AND2x2_ASAP7_75t_L g596 ( .A(n_453), .B(n_552), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_453), .B(n_581), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_453), .B(n_583), .Y(n_628) );
AND2x2_ASAP7_75t_L g687 ( .A(n_453), .B(n_632), .Y(n_687) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g557 ( .A(n_454), .B(n_464), .Y(n_557) );
AND2x2_ASAP7_75t_L g567 ( .A(n_454), .B(n_568), .Y(n_567) );
BUFx3_ASAP7_75t_L g589 ( .A(n_454), .Y(n_589) );
AND3x2_ASAP7_75t_L g648 ( .A(n_454), .B(n_649), .C(n_650), .Y(n_648) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_464), .Y(n_539) );
INVx1_ASAP7_75t_SL g583 ( .A(n_464), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_464), .B(n_532), .C(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_504), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_474), .A2(n_567), .B(n_619), .C(n_621), .Y(n_618) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_476), .B(n_495), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_476), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_SL g635 ( .A(n_476), .Y(n_635) );
AND2x2_ASAP7_75t_L g656 ( .A(n_476), .B(n_506), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_476), .B(n_565), .Y(n_684) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_486), .Y(n_476) );
AND2x2_ASAP7_75t_L g529 ( .A(n_477), .B(n_520), .Y(n_529) );
INVx2_ASAP7_75t_L g536 ( .A(n_477), .Y(n_536) );
AND2x2_ASAP7_75t_L g556 ( .A(n_477), .B(n_506), .Y(n_556) );
AND2x2_ASAP7_75t_L g606 ( .A(n_477), .B(n_495), .Y(n_606) );
INVx1_ASAP7_75t_L g610 ( .A(n_477), .Y(n_610) );
INVx2_ASAP7_75t_SL g520 ( .A(n_486), .Y(n_520) );
BUFx2_ASAP7_75t_L g546 ( .A(n_486), .Y(n_546) );
AND2x2_ASAP7_75t_L g673 ( .A(n_486), .B(n_495), .Y(n_673) );
INVx3_ASAP7_75t_SL g506 ( .A(n_495), .Y(n_506) );
AND2x2_ASAP7_75t_L g528 ( .A(n_495), .B(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g535 ( .A(n_495), .B(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g565 ( .A(n_495), .B(n_525), .Y(n_565) );
OR2x2_ASAP7_75t_L g574 ( .A(n_495), .B(n_520), .Y(n_574) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_495), .Y(n_592) );
AND2x2_ASAP7_75t_L g597 ( .A(n_495), .B(n_550), .Y(n_597) );
AND2x2_ASAP7_75t_L g625 ( .A(n_495), .B(n_508), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_495), .B(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g663 ( .A(n_495), .B(n_507), .Y(n_663) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AND2x2_ASAP7_75t_L g587 ( .A(n_506), .B(n_536), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_506), .B(n_529), .Y(n_615) );
AND2x2_ASAP7_75t_L g633 ( .A(n_506), .B(n_550), .Y(n_633) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
AND2x2_ASAP7_75t_L g534 ( .A(n_508), .B(n_520), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_508), .B(n_563), .Y(n_562) );
BUFx3_ASAP7_75t_L g572 ( .A(n_508), .Y(n_572) );
OR2x2_ASAP7_75t_L g620 ( .A(n_508), .B(n_540), .Y(n_620) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_512), .B(n_519), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_510), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g526 ( .A(n_512), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_519), .Y(n_527) );
AND2x2_ASAP7_75t_L g555 ( .A(n_520), .B(n_525), .Y(n_555) );
INVx1_ASAP7_75t_L g563 ( .A(n_520), .Y(n_563) );
AND2x2_ASAP7_75t_L g658 ( .A(n_520), .B(n_536), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_530), .B1(n_533), .B2(n_537), .C1(n_541), .C2(n_544), .Y(n_521) );
INVx1_ASAP7_75t_L g653 ( .A(n_522), .Y(n_653) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .Y(n_522) );
AND2x2_ASAP7_75t_L g549 ( .A(n_523), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g560 ( .A(n_523), .B(n_529), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_523), .B(n_551), .Y(n_576) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_523), .A2(n_599), .B1(n_604), .B2(n_605), .C1(n_613), .C2(n_615), .Y(n_598) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g586 ( .A(n_525), .B(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_525), .B(n_606), .Y(n_646) );
AND2x2_ASAP7_75t_L g657 ( .A(n_525), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g665 ( .A(n_528), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_530), .B(n_581), .Y(n_644) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_532), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_532), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
INVx3_ASAP7_75t_L g547 ( .A(n_535), .Y(n_547) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_535), .A2(n_638), .B(n_641), .C(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_535), .B(n_572), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_535), .B(n_555), .Y(n_677) );
AND2x2_ASAP7_75t_L g550 ( .A(n_536), .B(n_546), .Y(n_550) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g577 ( .A(n_539), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_540), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g629 ( .A(n_540), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g668 ( .A(n_540), .B(n_568), .Y(n_668) );
INVx1_ASAP7_75t_L g680 ( .A(n_540), .Y(n_680) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_543), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g661 ( .A(n_546), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_SL g548 ( .A1(n_549), .A2(n_551), .B(n_553), .C(n_557), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_549), .A2(n_579), .B1(n_594), .B2(n_597), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_550), .B(n_564), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_550), .B(n_572), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_551), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g614 ( .A(n_551), .Y(n_614) );
AND2x2_ASAP7_75t_L g621 ( .A(n_551), .B(n_601), .Y(n_621) );
INVx2_ASAP7_75t_L g582 ( .A(n_552), .Y(n_582) );
INVxp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NOR4xp25_ASAP7_75t_L g559 ( .A(n_556), .B(n_560), .C(n_561), .D(n_564), .Y(n_559) );
INVx1_ASAP7_75t_SL g630 ( .A(n_557), .Y(n_630) );
AND2x2_ASAP7_75t_L g674 ( .A(n_557), .B(n_675), .Y(n_674) );
OAI211xp5_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_566), .B(n_569), .C(n_578), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_565), .B(n_635), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_567), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_685) );
INVx1_ASAP7_75t_SL g640 ( .A(n_568), .Y(n_640) );
AND2x2_ASAP7_75t_L g679 ( .A(n_568), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_572), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_576), .B(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_577), .B(n_602), .Y(n_662) );
OAI21xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_584), .B(n_586), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g654 ( .A(n_581), .Y(n_654) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
INVx2_ASAP7_75t_L g682 ( .A(n_582), .Y(n_682) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_583), .Y(n_609) );
OAI21xp33_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_593), .Y(n_588) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_589), .Y(n_601) );
OR2x2_ASAP7_75t_L g639 ( .A(n_589), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI21xp33_ASAP7_75t_SL g634 ( .A1(n_592), .A2(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_596), .A2(n_623), .B1(n_626), .B2(n_633), .C(n_634), .Y(n_622) );
INVx1_ASAP7_75t_SL g666 ( .A(n_597), .Y(n_666) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x2_ASAP7_75t_L g613 ( .A(n_601), .B(n_614), .Y(n_613) );
INVxp67_ASAP7_75t_L g650 ( .A(n_603), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_610), .B2(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g645 ( .A(n_606), .Y(n_645) );
INVxp67_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_609), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR4xp25_ASAP7_75t_L g616 ( .A(n_617), .B(n_651), .C(n_664), .D(n_676), .Y(n_616) );
NAND3xp33_ASAP7_75t_SL g617 ( .A(n_618), .B(n_622), .C(n_637), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_620), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_627), .B(n_632), .Y(n_636) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI221xp5_ASAP7_75t_SL g664 ( .A1(n_639), .A2(n_665), .B1(n_666), .B2(n_667), .C(n_669), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g655 ( .A1(n_641), .A2(n_656), .B(n_657), .C(n_659), .Y(n_655) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_642), .A2(n_660), .B1(n_662), .B2(n_663), .Y(n_659) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B(n_654), .C(n_655), .Y(n_651) );
INVx1_ASAP7_75t_L g670 ( .A(n_663), .Y(n_670) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI21xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_671), .B(n_674), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B1(n_681), .B2(n_683), .C(n_685), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx3_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
endmodule