module real_jpeg_25632_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_1),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_34),
.B1(n_52),
.B2(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_1),
.A2(n_34),
.B1(n_62),
.B2(n_64),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_22),
.B1(n_27),
.B2(n_34),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_2),
.A2(n_22),
.B1(n_27),
.B2(n_61),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_2),
.A2(n_31),
.B1(n_61),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_2),
.A2(n_52),
.B1(n_57),
.B2(n_61),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_7),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_7),
.A2(n_22),
.B1(n_27),
.B2(n_80),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_7),
.A2(n_62),
.B1(n_64),
.B2(n_80),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_52),
.B1(n_57),
.B2(n_80),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_8),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_9),
.A2(n_22),
.B1(n_27),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_9),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_62),
.B1(n_64),
.B2(n_94),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_9),
.A2(n_31),
.B1(n_40),
.B2(n_94),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_52),
.B1(n_57),
.B2(n_94),
.Y(n_196)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_11),
.A2(n_40),
.B1(n_79),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_11),
.A2(n_22),
.B1(n_27),
.B2(n_84),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_11),
.A2(n_62),
.B1(n_64),
.B2(n_84),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_11),
.A2(n_52),
.B1(n_57),
.B2(n_84),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_12),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_12),
.A2(n_39),
.B1(n_62),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_12),
.A2(n_39),
.B1(n_52),
.B2(n_57),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_12),
.A2(n_22),
.B1(n_27),
.B2(n_39),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_30),
.B1(n_78),
.B2(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_22),
.B1(n_27),
.B2(n_167),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_13),
.A2(n_62),
.B1(n_64),
.B2(n_167),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_13),
.A2(n_52),
.B1(n_57),
.B2(n_167),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_14),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_14),
.A2(n_22),
.B1(n_27),
.B2(n_117),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_14),
.A2(n_62),
.B1(n_64),
.B2(n_117),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_14),
.A2(n_52),
.B1(n_57),
.B2(n_117),
.Y(n_278)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_15),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_15),
.B(n_21),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_15),
.B(n_62),
.C(n_90),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_15),
.A2(n_22),
.B1(n_27),
.B2(n_191),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_132),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_15),
.A2(n_62),
.B1(n_64),
.B2(n_191),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_52),
.C(n_67),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_15),
.A2(n_51),
.B(n_279),
.Y(n_309)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_16),
.Y(n_107)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_16),
.Y(n_198)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_16),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_43),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_28),
.B(n_33),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_28),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_21),
.A2(n_28),
.B1(n_116),
.B2(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_21),
.A2(n_28),
.B1(n_38),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_22),
.A2(n_27),
.B1(n_90),
.B2(n_91),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_22),
.A2(n_26),
.B(n_190),
.C(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_22),
.B(n_244),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

NAND3xp33_ASAP7_75t_SL g192 ( 
.A(n_25),
.B(n_27),
.C(n_31),
.Y(n_192)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_28),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_28),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_28),
.A2(n_120),
.B(n_190),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_31),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_32),
.A2(n_76),
.B(n_81),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_32),
.B(n_83),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_32),
.A2(n_76),
.B1(n_118),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_32),
.A2(n_118),
.B1(n_140),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_32),
.A2(n_81),
.B(n_182),
.Y(n_181)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_37),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_37),
.B(n_357),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_356),
.B(n_358),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_344),
.B(n_355),
.Y(n_44)
);

OAI31xp33_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_142),
.A3(n_157),
.B(n_341),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_121),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_47),
.B(n_121),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_85),
.C(n_101),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_48),
.A2(n_85),
.B1(n_86),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_48),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_72),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_49),
.A2(n_50),
.B(n_74),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_58),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_50),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_54),
.B(n_56),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_56),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_51),
.A2(n_54),
.B1(n_106),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_51),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_51),
.A2(n_196),
.B1(n_198),
.B2(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_51),
.B(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_51),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_57),
.B1(n_67),
.B2(n_68),
.Y(n_69)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_57),
.B(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_70),
.B2(n_71),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_60),
.A2(n_65),
.B1(n_71),
.B2(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_62),
.A2(n_64),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_62),
.B(n_288),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_65),
.A2(n_71),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_65),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_65),
.A2(n_71),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_69),
.A2(n_97),
.B1(n_111),
.B2(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_69),
.A2(n_177),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_69),
.A2(n_217),
.B(n_252),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_69),
.B(n_191),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_71),
.B(n_218),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g190 ( 
.A(n_79),
.B(n_191),
.CON(n_190),
.SN(n_190)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_96),
.B(n_100),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_95),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_89),
.B1(n_93),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_88),
.A2(n_89),
.B1(n_134),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_88),
.A2(n_184),
.B(n_186),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_88),
.A2(n_186),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_89),
.A2(n_113),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_89),
.A2(n_170),
.B(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_95),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_97),
.A2(n_266),
.B(n_267),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_97),
.A2(n_267),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_101),
.A2(n_102),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.C(n_114),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_103),
.A2(n_104),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_105),
.Y(n_179)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_107),
.Y(n_294)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_112),
.B(n_114),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B(n_119),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_124),
.C(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_139),
.B2(n_141),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_135),
.B1(n_136),
.B2(n_138),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_136),
.C(n_139),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_131),
.A2(n_132),
.B1(n_185),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_131),
.A2(n_132),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_132),
.B(n_171),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_136),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_136),
.B(n_149),
.C(n_154),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_139),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_141),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_139),
.B(n_145),
.C(n_148),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_143),
.A2(n_342),
.B(n_343),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_156),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_144),
.B(n_156),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_150),
.Y(n_351)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_155),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_334),
.B(n_340),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_206),
.B(n_333),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_199),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_160),
.B(n_199),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_178),
.C(n_180),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_161),
.A2(n_162),
.B1(n_178),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_172),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_168),
.B2(n_169),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_168),
.C(n_172),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_176),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_178),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_180),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_187),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_181),
.B(n_183),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_187),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_193),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_189),
.B1(n_193),
.B2(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_191),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_194),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_198),
.Y(n_247)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_198),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_201),
.B(n_202),
.C(n_205),
.Y(n_339)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_236),
.B(n_327),
.C(n_332),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_230),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_230),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_220),
.C(n_223),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_209),
.A2(n_210),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_219),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_215),
.C(n_219),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.C(n_228),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_231),
.B(n_234),
.C(n_235),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_320),
.B(n_326),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_268),
.B(n_319),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_257),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_257),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.C(n_254),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_242),
.B(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_245),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B(n_248),
.Y(n_245)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_249),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_250),
.A2(n_254),
.B1(n_255),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_250),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_253),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_258),
.B(n_264),
.C(n_265),
.Y(n_325)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_313),
.B(n_318),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_289),
.B(n_312),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_283),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_283),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_277),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_276),
.C(n_277),
.Y(n_317)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_285),
.B1(n_287),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_298),
.B(n_311),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_296),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_296),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_293),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_299),
.A2(n_304),
.B(n_310),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_309),
.Y(n_304)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_317),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_329),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_339),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_339),
.Y(n_340)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_346),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_354),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_348),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_350),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_352),
.C(n_354),
.Y(n_357)
);


endmodule