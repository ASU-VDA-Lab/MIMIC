module fake_jpeg_19622_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_26),
.B(n_19),
.C(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_27),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_23),
.A3(n_14),
.B1(n_19),
.B2(n_26),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_27),
.C(n_18),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_24),
.B1(n_23),
.B2(n_14),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_52),
.B1(n_13),
.B2(n_15),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_28),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_35),
.B1(n_25),
.B2(n_21),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_24),
.B1(n_14),
.B2(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_17),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_44),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_64),
.B1(n_48),
.B2(n_46),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_17),
.B1(n_25),
.B2(n_20),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_20),
.C(n_25),
.Y(n_68)
);

FAx1_ASAP7_75t_SL g79 ( 
.A(n_68),
.B(n_0),
.CI(n_1),
.CON(n_79),
.SN(n_79)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_6),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_73),
.B1(n_77),
.B2(n_84),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_44),
.B1(n_50),
.B2(n_2),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_50),
.B1(n_1),
.B2(n_2),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_68),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_66),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_57),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_76),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_54),
.C(n_56),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.C(n_84),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_53),
.C(n_9),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_80),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_106),
.B(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_70),
.B1(n_78),
.B2(n_71),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_76),
.B1(n_82),
.B2(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_103),
.B(n_94),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_75),
.C(n_79),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_113),
.C(n_98),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_111),
.B(n_112),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_77),
.B1(n_86),
.B2(n_71),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_101),
.C(n_99),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_118),
.Y(n_120)
);

NOR3xp33_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_106),
.C(n_110),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_6),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_116),
.A3(n_97),
.B1(n_99),
.B2(n_79),
.C1(n_96),
.C2(n_72),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_83),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_123),
.A2(n_124),
.B(n_119),
.Y(n_126)
);

OAI31xp33_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_8),
.A3(n_10),
.B(n_11),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_5),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_120),
.C(n_4),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);


endmodule