module fake_jpeg_25603_n_217 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_18),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_34),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_15),
.B1(n_27),
.B2(n_19),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_36),
.B1(n_42),
.B2(n_49),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_77),
.B1(n_18),
.B2(n_37),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_55),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_33),
.B1(n_21),
.B2(n_26),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_25),
.B1(n_23),
.B2(n_16),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_70),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_31),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx6p67_ASAP7_75t_R g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_33),
.B1(n_35),
.B2(n_34),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_75),
.B1(n_63),
.B2(n_68),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_44),
.A2(n_26),
.B1(n_23),
.B2(n_16),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_74),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_40),
.B(n_29),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_29),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_21),
.B1(n_28),
.B2(n_33),
.Y(n_77)
);

AO21x2_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_30),
.B(n_37),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_82),
.A2(n_72),
.B1(n_62),
.B2(n_71),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_13),
.C(n_12),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_10),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_66),
.B1(n_77),
.B2(n_58),
.Y(n_104)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_13),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_86),
.B(n_10),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_30),
.B(n_37),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_72),
.B1(n_55),
.B2(n_30),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_53),
.B(n_18),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_73),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_30),
.C(n_37),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_20),
.C(n_2),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_75),
.B(n_74),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_102),
.A2(n_118),
.B(n_119),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_88),
.B1(n_97),
.B2(n_93),
.Y(n_134)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_108),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_115),
.B1(n_124),
.B2(n_82),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_65),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_107),
.B(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_76),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g118 ( 
.A1(n_82),
.A2(n_80),
.B(n_101),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_20),
.B(n_56),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_120),
.B(n_122),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_67),
.B(n_1),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_121),
.A2(n_0),
.B(n_2),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_125),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_24),
.B1(n_30),
.B2(n_20),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_137),
.B1(n_147),
.B2(n_121),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_133),
.A2(n_135),
.B1(n_140),
.B2(n_125),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_124),
.B1(n_119),
.B2(n_103),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_106),
.A2(n_95),
.B1(n_99),
.B2(n_93),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_99),
.B1(n_78),
.B2(n_4),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_0),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_3),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_105),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_150),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_160),
.B1(n_137),
.B2(n_141),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_155),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_102),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_156),
.B(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_117),
.C(n_118),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_134),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_145),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_135),
.B1(n_133),
.B2(n_146),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_128),
.A2(n_103),
.B(n_116),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

AOI22x1_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_126),
.B1(n_129),
.B2(n_140),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_171),
.B1(n_162),
.B2(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_169),
.B(n_154),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_176),
.Y(n_182)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_145),
.CI(n_127),
.CON(n_175),
.SN(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_175),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_157),
.C(n_160),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_183),
.C(n_185),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_144),
.B(n_177),
.Y(n_192)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_181),
.B(n_186),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_132),
.C(n_156),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_188),
.B(n_172),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_132),
.C(n_163),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_151),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_176),
.C(n_151),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_193),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_175),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_149),
.C(n_166),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_172),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_150),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_197),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_153),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_193),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_141),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_191),
.C(n_189),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_205),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_136),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_207),
.B(n_208),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_185),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g210 ( 
.A(n_206),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_136),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_208),
.C(n_198),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_214),
.A2(n_211),
.B(n_184),
.Y(n_215)
);

OAI321xp33_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_120),
.C(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_7),
.Y(n_217)
);


endmodule