module fake_jpeg_27868_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_7),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_53),
.B1(n_47),
.B2(n_45),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_66),
.B1(n_3),
.B2(n_4),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_69),
.B(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_54),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_57),
.B1(n_49),
.B2(n_61),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_67),
.B1(n_65),
.B2(n_55),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_60),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_89),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_59),
.C(n_47),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_59),
.C(n_62),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_103),
.B1(n_104),
.B2(n_86),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_58),
.C(n_63),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.C(n_100),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_63),
.C(n_64),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx5_ASAP7_75t_SL g99 ( 
.A(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_68),
.C(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_79),
.B(n_22),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_105),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_99),
.B1(n_101),
.B2(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_122),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_20),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_9),
.B1(n_43),
.B2(n_12),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_6),
.Y(n_128)
);

BUFx2_ASAP7_75t_SL g124 ( 
.A(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_130),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_132),
.C(n_134),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_6),
.B(n_7),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_135),
.B1(n_136),
.B2(n_18),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_8),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_11),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_25),
.C(n_31),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_42),
.B1(n_26),
.B2(n_27),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_142),
.C(n_144),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_130),
.B1(n_143),
.B2(n_148),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_139),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_127),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_134),
.B(n_142),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_144),
.C(n_146),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_33),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_37),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_38),
.Y(n_158)
);


endmodule