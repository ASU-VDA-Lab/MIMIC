module fake_jpeg_16648_n_349 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_349);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_51),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_0),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_56),
.Y(n_83)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_27),
.Y(n_77)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_23),
.B(n_0),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_35),
.B1(n_32),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_69),
.B1(n_50),
.B2(n_45),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_21),
.B1(n_30),
.B2(n_36),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_76),
.B1(n_52),
.B2(n_0),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_21),
.B1(n_30),
.B2(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_62),
.A2(n_40),
.B1(n_33),
.B2(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_32),
.B1(n_37),
.B2(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_37),
.B1(n_34),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_71),
.A2(n_79),
.B1(n_49),
.B2(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_41),
.B1(n_38),
.B2(n_34),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_77),
.Y(n_102)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_48),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_53),
.Y(n_94)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_96),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_92),
.B(n_18),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_50),
.B1(n_56),
.B2(n_2),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_106),
.B1(n_0),
.B2(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_58),
.B(n_13),
.Y(n_98)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_113),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_80),
.B(n_42),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_108),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_57),
.B1(n_52),
.B2(n_33),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_64),
.B(n_31),
.Y(n_108)
);

NOR2xp67_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_24),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_79),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_110),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_10),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_10),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_116),
.A2(n_66),
.B1(n_65),
.B2(n_63),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_121),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_132),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_137),
.B1(n_143),
.B2(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_89),
.B(n_78),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_84),
.C(n_67),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_106),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_140),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_75),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_139),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_73),
.B1(n_60),
.B2(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_52),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_111),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_95),
.A2(n_86),
.B1(n_63),
.B2(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_9),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_147),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_108),
.B(n_11),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_152),
.B(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_111),
.B(n_93),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_161),
.B(n_170),
.Y(n_186)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_155),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_108),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_167),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_130),
.A2(n_86),
.B1(n_99),
.B2(n_97),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_131),
.B1(n_147),
.B2(n_136),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_132),
.B(n_117),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_112),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_120),
.B(n_99),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_166),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_163),
.A2(n_143),
.B1(n_137),
.B2(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_121),
.B(n_134),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_179),
.A2(n_189),
.B(n_190),
.C(n_181),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_122),
.B(n_123),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_187),
.B(n_192),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_134),
.B1(n_148),
.B2(n_133),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_188),
.B1(n_190),
.B2(n_193),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_121),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_194),
.B(n_180),
.Y(n_198)
);

XOR2x2_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_142),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_165),
.A2(n_160),
.B1(n_150),
.B2(n_161),
.Y(n_188)
);

AND2x4_ASAP7_75t_SL g189 ( 
.A(n_169),
.B(n_156),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_151),
.B(n_160),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_131),
.B1(n_138),
.B2(n_127),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_146),
.B(n_142),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_200),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_210),
.B(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_172),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_201),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_185),
.A2(n_149),
.B1(n_155),
.B2(n_159),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_206),
.A2(n_209),
.B1(n_216),
.B2(n_203),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_162),
.B1(n_145),
.B2(n_127),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_166),
.B(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_158),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_154),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_168),
.B1(n_131),
.B2(n_145),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_218),
.B1(n_221),
.B2(n_189),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_168),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_216),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_146),
.C(n_139),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_171),
.C(n_144),
.Y(n_238)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_126),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_222),
.B(n_191),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_186),
.B(n_179),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_179),
.B(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_183),
.B1(n_176),
.B2(n_189),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_227),
.A2(n_245),
.B1(n_247),
.B2(n_206),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_174),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_228),
.B(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_231),
.A2(n_234),
.B(n_217),
.Y(n_254)
);

XOR2x2_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_202),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_183),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_237),
.C(n_238),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_179),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_176),
.C(n_171),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_243),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_220),
.B(n_128),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_195),
.A2(n_184),
.B1(n_182),
.B2(n_141),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_198),
.B(n_210),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_246),
.B(n_140),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_141),
.B1(n_118),
.B2(n_85),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_218),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_196),
.B1(n_227),
.B2(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_261),
.B1(n_262),
.B2(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_224),
.A2(n_221),
.B1(n_196),
.B2(n_217),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_252),
.B1(n_256),
.B2(n_260),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_224),
.A2(n_217),
.B1(n_209),
.B2(n_197),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_204),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_246),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_263),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_207),
.B(n_118),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_118),
.B1(n_107),
.B2(n_97),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_231),
.A2(n_107),
.B1(n_115),
.B2(n_90),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_267),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_233),
.B(n_111),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_243),
.Y(n_279)
);

XOR2x1_ASAP7_75t_SL g276 ( 
.A(n_269),
.B(n_241),
.Y(n_276)
);

BUFx12_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_275),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_280),
.B(n_269),
.Y(n_294)
);

INVxp33_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_284),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_285),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_236),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_237),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_240),
.C(n_228),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_238),
.C(n_245),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_288),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_247),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_250),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_90),
.Y(n_288)
);

A2O1A1Ixp33_ASAP7_75t_SL g289 ( 
.A1(n_270),
.A2(n_260),
.B(n_255),
.C(n_254),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_289),
.A2(n_297),
.B1(n_105),
.B2(n_103),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_298),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_251),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_303),
.Y(n_317)
);

XNOR2x1_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_276),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_262),
.Y(n_295)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_273),
.A2(n_266),
.B(n_105),
.C(n_103),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_87),
.Y(n_300)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

BUFx12_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_304),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_271),
.B(n_283),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_282),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_299),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_306),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_292),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_281),
.B1(n_277),
.B2(n_273),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_297),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_314),
.C(n_315),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_110),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_312),
.B(n_110),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_290),
.B1(n_289),
.B2(n_302),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_54),
.C(n_5),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_274),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_266),
.B1(n_4),
.B2(n_5),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_310),
.Y(n_319)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_317),
.B(n_307),
.C(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_322),
.B(n_326),
.C(n_328),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_323),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_324),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_318),
.C(n_308),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_309),
.A2(n_3),
.B(n_4),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_3),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_320),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_333),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_5),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_7),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_332),
.B(n_11),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_321),
.C(n_8),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_337),
.Y(n_345)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_7),
.B(n_8),
.Y(n_338)
);

OAI321xp33_ASAP7_75t_L g344 ( 
.A1(n_338),
.A2(n_339),
.A3(n_341),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_8),
.Y(n_341)
);

A2O1A1O1Ixp25_ASAP7_75t_L g343 ( 
.A1(n_340),
.A2(n_336),
.B(n_12),
.C(n_13),
.D(n_14),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_344),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_346),
.A2(n_345),
.B(n_342),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_16),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_16),
.B1(n_18),
.B2(n_333),
.Y(n_349)
);


endmodule