module fake_netlist_1_5687_n_494 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_494);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_494;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g68 ( .A(n_23), .Y(n_68) );
NOR2xp67_ASAP7_75t_L g69 ( .A(n_7), .B(n_40), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_41), .Y(n_70) );
INVxp33_ASAP7_75t_SL g71 ( .A(n_54), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_12), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_3), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_6), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_16), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_28), .Y(n_76) );
CKINVDCx20_ASAP7_75t_R g77 ( .A(n_64), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_21), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_48), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_15), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_56), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_29), .Y(n_82) );
INVxp67_ASAP7_75t_SL g83 ( .A(n_57), .Y(n_83) );
BUFx3_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_27), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_34), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_26), .Y(n_87) );
INVxp67_ASAP7_75t_L g88 ( .A(n_47), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_51), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_12), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_18), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_65), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_58), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_45), .B(n_61), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_55), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_59), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_46), .Y(n_99) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_76), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_90), .B(n_72), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_76), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_97), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_97), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_97), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_78), .Y(n_107) );
INVx3_ASAP7_75t_L g108 ( .A(n_91), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_97), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_97), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_78), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_73), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_74), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
NOR2x1_ASAP7_75t_L g116 ( .A(n_69), .B(n_0), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_74), .B(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_75), .B(n_1), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_100), .Y(n_121) );
BUFx2_ASAP7_75t_L g122 ( .A(n_86), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_81), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_84), .Y(n_124) );
INVx2_ASAP7_75t_SL g125 ( .A(n_122), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_122), .B(n_75), .Y(n_127) );
OR2x2_ASAP7_75t_L g128 ( .A(n_102), .B(n_80), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_104), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
BUFx3_ASAP7_75t_L g131 ( .A(n_124), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_120), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_112), .B(n_88), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_113), .Y(n_134) );
INVx4_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
INVx2_ASAP7_75t_SL g136 ( .A(n_115), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_110), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g138 ( .A(n_115), .B(n_86), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_117), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_104), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
AND2x6_ASAP7_75t_L g144 ( .A(n_118), .B(n_84), .Y(n_144) );
OAI21xp33_ASAP7_75t_L g145 ( .A1(n_117), .A2(n_80), .B(n_71), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_119), .B(n_92), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_104), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_107), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_107), .Y(n_150) );
XOR2xp5_ASAP7_75t_L g151 ( .A(n_116), .B(n_77), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_111), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_140), .A2(n_118), .B1(n_123), .B2(n_119), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_144), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_134), .B(n_123), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_140), .A2(n_124), .B1(n_111), .B2(n_98), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
INVx1_ASAP7_75t_SL g158 ( .A(n_144), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_137), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_137), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_131), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_136), .B(n_71), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_127), .B(n_116), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_136), .B(n_98), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_125), .B(n_108), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_135), .B(n_96), .Y(n_167) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_144), .A2(n_77), .B1(n_114), .B2(n_108), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_142), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_147), .B(n_108), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_144), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_127), .B(n_108), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_135), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_135), .B(n_114), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_143), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_147), .B(n_114), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_147), .B(n_114), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_125), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_147), .B(n_83), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_144), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_145), .B(n_96), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_130), .B(n_95), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_144), .A2(n_89), .B1(n_68), .B2(n_93), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_146), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
AND3x1_ASAP7_75t_SL g190 ( .A(n_163), .B(n_151), .C(n_70), .Y(n_190) );
BUFx10_ASAP7_75t_L g191 ( .A(n_167), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
OR2x6_ASAP7_75t_L g193 ( .A(n_154), .B(n_130), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_157), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_165), .B(n_132), .C(n_150), .Y(n_195) );
INVx5_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_155), .B(n_128), .Y(n_197) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_171), .B(n_166), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_153), .B(n_128), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_183), .A2(n_132), .B(n_126), .C(n_138), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_168), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_157), .Y(n_204) );
BUFx10_ASAP7_75t_L g205 ( .A(n_167), .Y(n_205) );
INVx2_ASAP7_75t_SL g206 ( .A(n_166), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_171), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_162), .A2(n_126), .B(n_146), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_169), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_166), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_167), .B(n_126), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_166), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_173), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_168), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_160), .Y(n_219) );
INVx1_ASAP7_75t_SL g220 ( .A(n_179), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_177), .B(n_126), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_163), .B(n_144), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_220), .B(n_158), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_193), .Y(n_224) );
INVx1_ASAP7_75t_SL g225 ( .A(n_200), .Y(n_225) );
AOI22xp33_ASAP7_75t_SL g226 ( .A1(n_202), .A2(n_185), .B1(n_163), .B2(n_151), .Y(n_226) );
NOR2xp67_ASAP7_75t_L g227 ( .A(n_217), .B(n_186), .Y(n_227) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_200), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_218), .A2(n_163), .B1(n_185), .B2(n_177), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_194), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_212), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_194), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_203), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_190), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_204), .A2(n_164), .B(n_185), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_212), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_208), .A2(n_186), .B(n_180), .C(n_188), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_204), .Y(n_238) );
OAI222xp33_ASAP7_75t_L g239 ( .A1(n_218), .A2(n_156), .B1(n_181), .B2(n_180), .C1(n_175), .C2(n_188), .Y(n_239) );
AOI221xp5_ASAP7_75t_L g240 ( .A1(n_197), .A2(n_172), .B1(n_133), .B2(n_177), .C(n_176), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_212), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_189), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_191), .Y(n_244) );
OAI222xp33_ASAP7_75t_L g245 ( .A1(n_215), .A2(n_175), .B1(n_158), .B2(n_182), .C1(n_170), .C2(n_177), .Y(n_245) );
CKINVDCx8_ASAP7_75t_R g246 ( .A(n_196), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_199), .B(n_172), .Y(n_247) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_240), .A2(n_239), .B1(n_226), .B2(n_247), .C(n_229), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_234), .A2(n_191), .B1(n_205), .B2(n_215), .Y(n_249) );
OAI221xp5_ASAP7_75t_L g250 ( .A1(n_235), .A2(n_222), .B1(n_201), .B2(n_195), .C(n_214), .Y(n_250) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_225), .A2(n_209), .B1(n_214), .B2(n_193), .Y(n_251) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_237), .A2(n_195), .B(n_221), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_224), .A2(n_205), .B1(n_191), .B2(n_221), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_224), .A2(n_193), .B1(n_205), .B2(n_182), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_246), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_230), .A2(n_221), .B1(n_174), .B2(n_152), .C(n_150), .Y(n_257) );
AOI22xp33_ASAP7_75t_SL g258 ( .A1(n_244), .A2(n_193), .B1(n_196), .B2(n_217), .Y(n_258) );
INVx4_ASAP7_75t_L g259 ( .A(n_231), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_232), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_227), .A2(n_221), .B1(n_193), .B2(n_174), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g263 ( .A1(n_227), .A2(n_174), .B1(n_217), .B2(n_216), .Y(n_263) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_174), .B1(n_149), .B2(n_152), .C(n_139), .Y(n_264) );
AO222x2_ASAP7_75t_L g265 ( .A1(n_238), .A2(n_1), .B1(n_2), .B2(n_3), .C1(n_4), .C2(n_5), .Y(n_265) );
AOI22xp33_ASAP7_75t_SL g266 ( .A1(n_231), .A2(n_196), .B1(n_211), .B2(n_203), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_243), .A2(n_149), .B1(n_216), .B2(n_131), .C(n_213), .Y(n_267) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_243), .A2(n_219), .B1(n_211), .B2(n_196), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_254), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_260), .Y(n_270) );
OR2x2_ASAP7_75t_L g271 ( .A(n_261), .B(n_233), .Y(n_271) );
OAI211xp5_ASAP7_75t_L g272 ( .A1(n_248), .A2(n_246), .B(n_82), .C(n_85), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_259), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_249), .B(n_228), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_259), .B(n_233), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_252), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_256), .Y(n_277) );
NAND4xp25_ASAP7_75t_L g278 ( .A(n_265), .B(n_87), .C(n_94), .D(n_99), .Y(n_278) );
OR2x2_ASAP7_75t_L g279 ( .A(n_251), .B(n_233), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_262), .A2(n_231), .B1(n_236), .B2(n_241), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_250), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_257), .A2(n_231), .B1(n_236), .B2(n_241), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_268), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_268), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_253), .B(n_219), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_255), .A2(n_241), .B1(n_236), .B2(n_223), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_263), .B(n_242), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_255), .A2(n_236), .B1(n_241), .B2(n_216), .Y(n_289) );
AOI211x1_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_245), .B(n_4), .C(n_5), .Y(n_290) );
AND2x4_ASAP7_75t_SL g291 ( .A(n_266), .B(n_242), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_267), .A2(n_210), .B(n_198), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_278), .B(n_2), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_270), .Y(n_294) );
NAND2xp33_ASAP7_75t_SL g295 ( .A(n_273), .B(n_242), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_270), .B(n_6), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_270), .B(n_100), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_269), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_269), .B(n_100), .Y(n_299) );
OA211x2_ASAP7_75t_L g300 ( .A1(n_289), .A2(n_264), .B(n_8), .C(n_9), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_273), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_271), .B(n_7), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_276), .Y(n_303) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_278), .A2(n_100), .B1(n_178), .B2(n_184), .C(n_187), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_275), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_271), .B(n_8), .Y(n_306) );
NAND4xp25_ASAP7_75t_L g307 ( .A(n_290), .B(n_110), .C(n_10), .D(n_11), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_276), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_290), .B(n_9), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_285), .B(n_242), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_288), .B(n_242), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_281), .Y(n_316) );
AOI33xp33_ASAP7_75t_L g317 ( .A1(n_282), .A2(n_110), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_273), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_273), .Y(n_319) );
INVx3_ASAP7_75t_SL g320 ( .A(n_273), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_291), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_282), .B(n_11), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_281), .B(n_242), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_277), .B(n_13), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_291), .Y(n_326) );
AOI21xp33_ASAP7_75t_L g327 ( .A1(n_322), .A2(n_272), .B(n_281), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_314), .B(n_284), .Y(n_328) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_326), .B(n_284), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_298), .Y(n_330) );
INVx4_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_298), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_315), .Y(n_333) );
OAI33xp33_ASAP7_75t_L g334 ( .A1(n_307), .A2(n_274), .A3(n_280), .B1(n_283), .B2(n_286), .B3(n_14), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_293), .B(n_104), .C(n_105), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_317), .B(n_104), .C(n_105), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_294), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_305), .B(n_291), .Y(n_339) );
OR2x6_ASAP7_75t_L g340 ( .A(n_326), .B(n_284), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_284), .B1(n_287), .B2(n_292), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_325), .B(n_105), .C(n_106), .Y(n_342) );
OAI322xp33_ASAP7_75t_L g343 ( .A1(n_302), .A2(n_105), .A3(n_106), .B1(n_109), .B2(n_121), .C1(n_187), .C2(n_184), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_307), .B(n_121), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_315), .B(n_121), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_296), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_306), .A2(n_198), .B1(n_206), .B2(n_213), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_312), .B(n_109), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_306), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_312), .B(n_109), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_309), .B(n_105), .C(n_106), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_313), .B(n_109), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_316), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_310), .B(n_106), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_310), .B(n_106), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_311), .B(n_17), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_299), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g358 ( .A1(n_299), .A2(n_184), .B1(n_178), .B2(n_187), .C(n_206), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_311), .B(n_178), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_311), .B(n_19), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_320), .B(n_303), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_297), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_320), .B(n_161), .Y(n_363) );
OAI21xp33_ASAP7_75t_L g364 ( .A1(n_297), .A2(n_129), .B(n_141), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_303), .B(n_161), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_303), .Y(n_366) );
OAI211xp5_ASAP7_75t_SL g367 ( .A1(n_318), .A2(n_173), .B(n_160), .C(n_210), .Y(n_367) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_321), .B(n_308), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_334), .A2(n_308), .B1(n_324), .B2(n_323), .C(n_319), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_333), .B(n_301), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_333), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_349), .B(n_301), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_330), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_332), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_328), .B(n_324), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_331), .A2(n_300), .B1(n_301), .B2(n_323), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_353), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_328), .B(n_20), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_337), .A2(n_295), .B(n_300), .C(n_210), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_355), .B(n_22), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_346), .B(n_24), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_339), .B(n_25), .Y(n_382) );
NOR2x1_ASAP7_75t_L g383 ( .A(n_331), .B(n_207), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_354), .Y(n_384) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_331), .Y(n_385) );
BUFx2_ASAP7_75t_L g386 ( .A(n_361), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_345), .B(n_30), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_362), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_355), .B(n_31), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_345), .B(n_33), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_362), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_335), .B(n_207), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_363), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_348), .B(n_35), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_348), .B(n_36), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_336), .B(n_37), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_357), .B(n_38), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_364), .B(n_196), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_350), .B(n_42), .Y(n_400) );
AOI211xp5_ASAP7_75t_SL g401 ( .A1(n_343), .A2(n_173), .B(n_44), .C(n_49), .Y(n_401) );
AOI32xp33_ASAP7_75t_L g402 ( .A1(n_344), .A2(n_173), .A3(n_50), .B1(n_52), .B2(n_53), .Y(n_402) );
AND2x4_ASAP7_75t_L g403 ( .A(n_340), .B(n_43), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_338), .B(n_60), .Y(n_404) );
INVxp67_ASAP7_75t_L g405 ( .A(n_350), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_352), .B(n_63), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_327), .B(n_66), .Y(n_407) );
NAND2xp33_ASAP7_75t_L g408 ( .A(n_402), .B(n_347), .Y(n_408) );
AOI32xp33_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_356), .A3(n_360), .B1(n_352), .B2(n_367), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_371), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_373), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_388), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_386), .B(n_340), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_391), .B(n_360), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_377), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_388), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_391), .B(n_384), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_398), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_341), .B1(n_340), .B2(n_342), .Y(n_421) );
OAI211xp5_ASAP7_75t_SL g422 ( .A1(n_379), .A2(n_359), .B(n_358), .C(n_351), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_368), .B(n_370), .Y(n_424) );
INVx1_ASAP7_75t_SL g425 ( .A(n_393), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_369), .B(n_365), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_405), .B(n_329), .Y(n_427) );
AOI222xp33_ASAP7_75t_L g428 ( .A1(n_375), .A2(n_129), .B1(n_141), .B2(n_148), .C1(n_161), .C2(n_196), .Y(n_428) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_403), .B(n_207), .Y(n_429) );
XOR2x2_ASAP7_75t_L g430 ( .A(n_401), .B(n_67), .Y(n_430) );
XOR2xp5_ASAP7_75t_L g431 ( .A(n_376), .B(n_198), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_375), .B(n_129), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_392), .B(n_207), .Y(n_433) );
INVxp67_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_396), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_407), .B(n_141), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_399), .A2(n_189), .B1(n_192), .B2(n_207), .Y(n_438) );
XNOR2x1_ASAP7_75t_L g439 ( .A(n_382), .B(n_189), .Y(n_439) );
NAND2xp33_ASAP7_75t_SL g440 ( .A(n_403), .B(n_189), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_403), .B(n_161), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_394), .B(n_148), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_407), .A2(n_148), .B1(n_189), .B2(n_192), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_SL g445 ( .A1(n_379), .A2(n_148), .B(n_192), .C(n_400), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g446 ( .A1(n_381), .A2(n_148), .B(n_192), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_397), .Y(n_447) );
OA22x2_ASAP7_75t_L g448 ( .A1(n_394), .A2(n_148), .B1(n_192), .B2(n_395), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_380), .B(n_389), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_380), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_389), .B(n_395), .Y(n_451) );
AOI322xp5_ASAP7_75t_L g452 ( .A1(n_387), .A2(n_390), .A3(n_406), .B1(n_293), .B2(n_371), .C1(n_385), .C2(n_349), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_371), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g454 ( .A1(n_376), .A2(n_278), .B(n_293), .C(n_391), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_385), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_385), .A2(n_278), .B1(n_293), .B2(n_334), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_371), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_371), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_455), .B(n_420), .Y(n_459) );
AOI221xp5_ASAP7_75t_L g460 ( .A1(n_454), .A2(n_426), .B1(n_423), .B2(n_456), .C(n_424), .Y(n_460) );
XOR2x2_ASAP7_75t_L g461 ( .A(n_439), .B(n_448), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_420), .B(n_425), .Y(n_464) );
XNOR2x2_ASAP7_75t_L g465 ( .A(n_448), .B(n_429), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_417), .B(n_458), .Y(n_466) );
OAI321xp33_ASAP7_75t_L g467 ( .A1(n_409), .A2(n_427), .A3(n_421), .B1(n_424), .B2(n_434), .C(n_449), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_457), .B(n_410), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_434), .B(n_414), .Y(n_469) );
OAI21xp5_ASAP7_75t_SL g470 ( .A1(n_452), .A2(n_431), .B(n_441), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_408), .A2(n_427), .B1(n_450), .B2(n_435), .Y(n_471) );
XNOR2xp5_ASAP7_75t_L g472 ( .A(n_451), .B(n_430), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_418), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_461), .A2(n_447), .B1(n_451), .B2(n_436), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_459), .A2(n_445), .B(n_440), .Y(n_475) );
OAI21xp33_ASAP7_75t_SL g476 ( .A1(n_471), .A2(n_460), .B(n_473), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_470), .B(n_432), .C(n_437), .Y(n_477) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_469), .B(n_444), .C(n_422), .D(n_428), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_472), .A2(n_453), .B1(n_413), .B2(n_411), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_466), .Y(n_480) );
AO22x2_ASAP7_75t_L g481 ( .A1(n_462), .A2(n_416), .B1(n_419), .B2(n_433), .Y(n_481) );
NOR2xp67_ASAP7_75t_SL g482 ( .A(n_475), .B(n_467), .Y(n_482) );
XNOR2xp5_ASAP7_75t_L g483 ( .A(n_479), .B(n_464), .Y(n_483) );
NOR2x1p5_ASAP7_75t_L g484 ( .A(n_477), .B(n_463), .Y(n_484) );
NOR2xp67_ASAP7_75t_L g485 ( .A(n_476), .B(n_469), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_482), .Y(n_486) );
AOI22xp5_ASAP7_75t_SL g487 ( .A1(n_483), .A2(n_465), .B1(n_480), .B2(n_481), .Y(n_487) );
OAI222xp33_ASAP7_75t_L g488 ( .A1(n_483), .A2(n_474), .B1(n_468), .B2(n_478), .C1(n_415), .C2(n_443), .Y(n_488) );
NOR2xp67_ASAP7_75t_L g489 ( .A(n_486), .B(n_485), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_486), .Y(n_490) );
OR3x1_ASAP7_75t_L g491 ( .A(n_490), .B(n_487), .C(n_488), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_491), .A2(n_489), .B(n_484), .Y(n_492) );
XNOR2xp5_ASAP7_75t_L g493 ( .A(n_492), .B(n_442), .Y(n_493) );
AOI221xp5_ASAP7_75t_L g494 ( .A1(n_493), .A2(n_422), .B1(n_438), .B2(n_446), .C(n_433), .Y(n_494) );
endmodule