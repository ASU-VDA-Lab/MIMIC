module fake_jpeg_4525_n_325 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_8),
.B(n_14),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_49),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_52),
.Y(n_69)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_61),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_57),
.A2(n_64),
.B1(n_79),
.B2(n_37),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_60),
.A2(n_62),
.B1(n_75),
.B2(n_83),
.Y(n_135)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_76),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_25),
.B1(n_33),
.B2(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_24),
.B1(n_17),
.B2(n_18),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_77),
.B1(n_80),
.B2(n_87),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_68),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_99),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_19),
.B1(n_24),
.B2(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_35),
.B1(n_31),
.B2(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_29),
.B1(n_33),
.B2(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_86),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_16),
.B1(n_21),
.B2(n_37),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_47),
.B(n_16),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_84),
.A2(n_104),
.B(n_5),
.C(n_6),
.Y(n_136)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_53),
.A2(n_34),
.B1(n_15),
.B2(n_21),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_92),
.Y(n_121)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_16),
.B1(n_21),
.B2(n_37),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_27),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_103),
.Y(n_123)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_97),
.Y(n_126)
);

BUFx12_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_1),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_27),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_2),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_27),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g104 ( 
.A1(n_48),
.A2(n_37),
.B1(n_27),
.B2(n_4),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_118),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_117),
.Y(n_142)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_120),
.B(n_69),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_57),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_133),
.B1(n_100),
.B2(n_102),
.Y(n_144)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_98),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_2),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_129),
.A2(n_109),
.B(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_72),
.B(n_79),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_74),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_84),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_104),
.A2(n_2),
.B(n_3),
.C(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_136),
.B1(n_129),
.B2(n_115),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_136),
.A2(n_94),
.B(n_58),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_71),
.B1(n_88),
.B2(n_90),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_153),
.B1(n_155),
.B2(n_159),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_147),
.B(n_116),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_143),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_92),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_145),
.B1(n_167),
.B2(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_103),
.B1(n_94),
.B2(n_73),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_156),
.Y(n_179)
);

AND2x4_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_103),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_89),
.C(n_85),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_151),
.C(n_119),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_99),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_82),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_173),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_157),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_113),
.A2(n_101),
.B1(n_82),
.B2(n_70),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_86),
.B1(n_66),
.B2(n_61),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_162),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_97),
.B1(n_56),
.B2(n_95),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_168),
.B1(n_170),
.B2(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

INVx13_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_76),
.Y(n_165)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_166),
.A2(n_126),
.B(n_134),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_129),
.B(n_96),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_120),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_113),
.A2(n_136),
.B1(n_117),
.B2(n_109),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_117),
.A2(n_78),
.B1(n_63),
.B2(n_98),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_134),
.B(n_119),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_108),
.B(n_6),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_128),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_194),
.C(n_201),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_180),
.A2(n_184),
.B(n_185),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_181),
.A2(n_189),
.B1(n_205),
.B2(n_150),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_134),
.B(n_133),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_147),
.A2(n_134),
.B(n_105),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_192),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_168),
.B1(n_155),
.B2(n_137),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_105),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_196),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_139),
.B(n_126),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_143),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_204),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g237 ( 
.A(n_197),
.B(n_141),
.C(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_203),
.Y(n_215)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_106),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_106),
.B1(n_132),
.B2(n_112),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_209),
.B(n_145),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_124),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_195),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_214),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_212),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_178),
.B(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_178),
.B(n_166),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

OAI32xp33_ASAP7_75t_L g222 ( 
.A1(n_209),
.A2(n_167),
.A3(n_150),
.B1(n_142),
.B2(n_138),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_229),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_236),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_160),
.B1(n_179),
.B2(n_162),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_142),
.B(n_141),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_233),
.Y(n_248)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_194),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_148),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_186),
.C(n_175),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_157),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_215),
.B(n_196),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_229),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_201),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_250),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_235),
.A2(n_189),
.B1(n_207),
.B2(n_181),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_246),
.A2(n_253),
.B1(n_226),
.B2(n_232),
.Y(n_267)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_218),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_193),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_252),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_175),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_203),
.B1(n_184),
.B2(n_185),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_254),
.A2(n_219),
.B1(n_236),
.B2(n_225),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_156),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_190),
.C(n_191),
.Y(n_258)
);

OAI321xp33_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_176),
.A3(n_134),
.B1(n_190),
.B2(n_206),
.C(n_200),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_230),
.B(n_215),
.C(n_224),
.D(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_266),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_212),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_267),
.A2(n_269),
.B1(n_270),
.B2(n_276),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_216),
.B1(n_221),
.B2(n_220),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_253),
.A2(n_217),
.B1(n_211),
.B2(n_223),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_260),
.B1(n_248),
.B2(n_240),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_271),
.A2(n_254),
.B1(n_239),
.B2(n_243),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_228),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_176),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_274),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_249),
.B1(n_239),
.B2(n_250),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_233),
.B1(n_222),
.B2(n_228),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_214),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_242),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_272),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_285),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_268),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_171),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_283),
.Y(n_298)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_255),
.C(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_282),
.B(n_267),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_291),
.Y(n_301)
);

AOI321xp33_ASAP7_75t_L g285 ( 
.A1(n_261),
.A2(n_243),
.A3(n_245),
.B1(n_252),
.B2(n_257),
.C(n_258),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_265),
.A2(n_241),
.B1(n_247),
.B2(n_182),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_269),
.B1(n_262),
.B2(n_266),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_124),
.C(n_65),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_182),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_293),
.A2(n_299),
.B(n_302),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_264),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_297),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_268),
.B1(n_264),
.B2(n_202),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_183),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_132),
.B(n_183),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_298),
.C(n_301),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_278),
.B(n_290),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_286),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_287),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_310),
.B(n_300),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_169),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_308),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.C(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_154),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_154),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_316),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_318),
.C(n_312),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_202),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_6),
.C(n_7),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_294),
.C(n_292),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_312),
.A2(n_6),
.B(n_7),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_321),
.C(n_314),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_322),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_319),
.Y(n_325)
);


endmodule