module real_aes_17829_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_1672;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1691;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1647;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1330 ( .A(n_0), .Y(n_1330) );
OAI211xp5_ASAP7_75t_L g455 ( .A1(n_1), .A2(n_446), .B(n_456), .C(n_460), .Y(n_455) );
INVx1_ASAP7_75t_L g506 ( .A(n_1), .Y(n_506) );
INVx1_ASAP7_75t_L g655 ( .A(n_2), .Y(n_655) );
OAI211xp5_ASAP7_75t_L g701 ( .A1(n_2), .A2(n_702), .B(n_704), .C(n_713), .Y(n_701) );
INVx1_ASAP7_75t_L g328 ( .A(n_3), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_3), .B(n_338), .Y(n_354) );
AND2x2_ASAP7_75t_L g538 ( .A(n_3), .B(n_485), .Y(n_538) );
AND2x2_ASAP7_75t_L g605 ( .A(n_3), .B(n_229), .Y(n_605) );
OAI211xp5_ASAP7_75t_SL g1348 ( .A1(n_4), .A2(n_1183), .B(n_1257), .C(n_1349), .Y(n_1348) );
INVx1_ASAP7_75t_L g1359 ( .A(n_4), .Y(n_1359) );
INVx1_ASAP7_75t_L g785 ( .A(n_5), .Y(n_785) );
INVx1_ASAP7_75t_L g958 ( .A(n_6), .Y(n_958) );
INVx1_ASAP7_75t_L g1368 ( .A(n_7), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_8), .A2(n_141), .B1(n_1055), .B2(n_1173), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g1189 ( .A1(n_8), .A2(n_141), .B1(n_880), .B2(n_1190), .Y(n_1189) );
OAI22xp33_ASAP7_75t_L g1177 ( .A1(n_9), .A2(n_248), .B1(n_330), .B2(n_821), .Y(n_1177) );
OAI22xp33_ASAP7_75t_L g1185 ( .A1(n_9), .A2(n_248), .B1(n_1049), .B2(n_1100), .Y(n_1185) );
OAI211xp5_ASAP7_75t_L g783 ( .A1(n_10), .A2(n_414), .B(n_671), .C(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g798 ( .A(n_10), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_11), .A2(n_71), .B1(n_680), .B2(n_681), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g976 ( .A1(n_11), .A2(n_19), .B1(n_977), .B2(n_979), .C(n_980), .Y(n_976) );
INVx1_ASAP7_75t_L g1005 ( .A(n_12), .Y(n_1005) );
INVx1_ASAP7_75t_L g522 ( .A(n_13), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_14), .A2(n_167), .B1(n_690), .B2(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g705 ( .A(n_14), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_15), .A2(n_27), .B1(n_632), .B2(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g939 ( .A(n_15), .Y(n_939) );
INVx1_ASAP7_75t_L g1392 ( .A(n_16), .Y(n_1392) );
OAI211xp5_ASAP7_75t_L g1398 ( .A1(n_16), .A2(n_456), .B(n_1399), .C(n_1400), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1098 ( .A1(n_17), .A2(n_156), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_17), .A2(n_156), .B1(n_330), .B2(n_791), .Y(n_1102) );
INVx1_ASAP7_75t_L g1371 ( .A(n_18), .Y(n_1371) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_19), .A2(n_219), .B1(n_898), .B2(n_968), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g1286 ( .A(n_20), .Y(n_1286) );
INVx2_ASAP7_75t_L g405 ( .A(n_21), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g1429 ( .A1(n_22), .A2(n_24), .B1(n_1413), .B2(n_1420), .Y(n_1429) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_23), .A2(n_311), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g627 ( .A(n_23), .Y(n_627) );
INVx1_ASAP7_75t_L g1146 ( .A(n_25), .Y(n_1146) );
INVx1_ASAP7_75t_L g1333 ( .A(n_26), .Y(n_1333) );
AOI221xp5_ASAP7_75t_L g918 ( .A1(n_27), .A2(n_40), .B1(n_613), .B2(n_919), .C(n_921), .Y(n_918) );
INVx1_ASAP7_75t_L g962 ( .A(n_28), .Y(n_962) );
INVx1_ASAP7_75t_L g1022 ( .A(n_29), .Y(n_1022) );
INVx1_ASAP7_75t_L g1377 ( .A(n_30), .Y(n_1377) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_31), .Y(n_323) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_31), .B(n_321), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_32), .A2(n_189), .B1(n_1413), .B2(n_1469), .Y(n_1482) );
INVx1_ASAP7_75t_L g1254 ( .A(n_33), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_34), .A2(n_194), .B1(n_588), .B2(n_590), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_34), .A2(n_239), .B1(n_643), .B2(n_645), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g899 ( .A1(n_35), .A2(n_202), .B1(n_434), .B2(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g924 ( .A(n_35), .Y(n_924) );
INVx1_ASAP7_75t_L g548 ( .A(n_36), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g1679 ( .A(n_37), .Y(n_1679) );
CKINVDCx5p33_ASAP7_75t_R g1290 ( .A(n_38), .Y(n_1290) );
INVx1_ASAP7_75t_L g828 ( .A(n_39), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_40), .A2(n_288), .B1(n_898), .B2(n_906), .Y(n_905) );
INVxp67_ASAP7_75t_SL g961 ( .A(n_41), .Y(n_961) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_41), .A2(n_166), .B1(n_387), .B2(n_986), .Y(n_985) );
INVx1_ASAP7_75t_L g742 ( .A(n_42), .Y(n_742) );
INVx1_ASAP7_75t_L g1014 ( .A(n_43), .Y(n_1014) );
INVx1_ASAP7_75t_L g838 ( .A(n_44), .Y(n_838) );
INVx1_ASAP7_75t_L g1075 ( .A(n_45), .Y(n_1075) );
INVx1_ASAP7_75t_L g972 ( .A(n_46), .Y(n_972) );
INVx1_ASAP7_75t_L g676 ( .A(n_47), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_47), .A2(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_L g1094 ( .A(n_48), .Y(n_1094) );
AOI22xp5_ASAP7_75t_L g1467 ( .A1(n_49), .A2(n_201), .B1(n_1420), .B2(n_1423), .Y(n_1467) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_50), .A2(n_133), .B1(n_472), .B2(n_788), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_50), .A2(n_133), .B1(n_508), .B2(n_800), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_51), .Y(n_960) );
INVx1_ASAP7_75t_L g996 ( .A(n_52), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g1438 ( .A1(n_52), .A2(n_303), .B1(n_1413), .B2(n_1417), .Y(n_1438) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_53), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_54), .A2(n_69), .B1(n_902), .B2(n_904), .Y(n_901) );
INVx1_ASAP7_75t_L g923 ( .A(n_54), .Y(n_923) );
INVx1_ASAP7_75t_L g1071 ( .A(n_55), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_56), .A2(n_99), .B1(n_616), .B2(n_1124), .Y(n_1123) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_56), .A2(n_212), .B1(n_434), .B2(n_965), .Y(n_1156) );
INVx1_ASAP7_75t_L g667 ( .A(n_57), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_57), .A2(n_280), .B1(n_698), .B2(n_700), .Y(n_697) );
XNOR2xp5_ASAP7_75t_L g1000 ( .A(n_58), .B(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1258 ( .A(n_59), .Y(n_1258) );
INVx1_ASAP7_75t_L g1196 ( .A(n_60), .Y(n_1196) );
AOI21xp33_ASAP7_75t_L g1639 ( .A1(n_61), .A2(n_585), .B(n_1640), .Y(n_1639) );
AOI221xp5_ASAP7_75t_L g1654 ( .A1(n_61), .A2(n_241), .B1(n_900), .B2(n_1655), .C(n_1657), .Y(n_1654) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_62), .Y(n_889) );
XOR2x2_ASAP7_75t_L g1111 ( .A(n_63), .B(n_1112), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1468 ( .A1(n_64), .A2(n_287), .B1(n_1413), .B2(n_1469), .Y(n_1468) );
OAI22xp33_ASAP7_75t_L g1300 ( .A1(n_65), .A2(n_112), .B1(n_330), .B2(n_791), .Y(n_1300) );
OAI22xp33_ASAP7_75t_L g1310 ( .A1(n_65), .A2(n_112), .B1(n_452), .B2(n_1049), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1419 ( .A1(n_66), .A2(n_120), .B1(n_1420), .B2(n_1423), .Y(n_1419) );
OAI222xp33_ASAP7_75t_L g1620 ( .A1(n_67), .A2(n_75), .B1(n_80), .B2(n_524), .C1(n_1621), .C2(n_1622), .Y(n_1620) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_68), .A2(n_609), .B(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_68), .A2(n_194), .B1(n_629), .B2(n_632), .Y(n_628) );
INVx1_ASAP7_75t_L g944 ( .A(n_69), .Y(n_944) );
INVx1_ASAP7_75t_L g1047 ( .A(n_70), .Y(n_1047) );
OAI211xp5_ASAP7_75t_L g1060 ( .A1(n_70), .A2(n_793), .B(n_812), .C(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g995 ( .A(n_71), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g822 ( .A1(n_72), .A2(n_76), .B1(n_823), .B2(n_824), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g878 ( .A1(n_72), .A2(n_76), .B1(n_879), .B2(n_880), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g1627 ( .A(n_73), .Y(n_1627) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_74), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_77), .A2(n_275), .B1(n_362), .B2(n_387), .Y(n_932) );
INVx1_ASAP7_75t_L g946 ( .A(n_77), .Y(n_946) );
INVx1_ASAP7_75t_L g849 ( .A(n_78), .Y(n_849) );
XOR2x2_ASAP7_75t_L g1224 ( .A(n_79), .B(n_1225), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g1646 ( .A1(n_80), .A2(n_309), .B1(n_700), .B2(n_1647), .Y(n_1646) );
INVx1_ASAP7_75t_L g1325 ( .A(n_81), .Y(n_1325) );
INVx1_ASAP7_75t_L g1350 ( .A(n_82), .Y(n_1350) );
AOI22xp5_ASAP7_75t_L g1445 ( .A1(n_83), .A2(n_308), .B1(n_1420), .B2(n_1423), .Y(n_1445) );
AOI22xp33_ASAP7_75t_SL g1665 ( .A1(n_83), .A2(n_1666), .B1(n_1715), .B2(n_1718), .Y(n_1665) );
XNOR2xp5_ASAP7_75t_L g1668 ( .A(n_83), .B(n_1669), .Y(n_1668) );
INVx1_ASAP7_75t_L g1230 ( .A(n_84), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g1641 ( .A1(n_85), .A2(n_153), .B1(n_590), .B2(n_612), .Y(n_1641) );
INVx1_ASAP7_75t_L g1652 ( .A(n_85), .Y(n_1652) );
INVx1_ASAP7_75t_L g1012 ( .A(n_86), .Y(n_1012) );
XNOR2xp5_ASAP7_75t_L g737 ( .A(n_87), .B(n_738), .Y(n_737) );
CKINVDCx5p33_ASAP7_75t_R g971 ( .A(n_88), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_89), .A2(n_290), .B1(n_902), .B2(n_965), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g992 ( .A1(n_89), .A2(n_200), .B1(n_613), .B2(n_711), .C(n_993), .Y(n_992) );
OAI211xp5_ASAP7_75t_L g1178 ( .A1(n_90), .A2(n_1179), .B(n_1180), .C(n_1183), .Y(n_1178) );
INVx1_ASAP7_75t_L g1188 ( .A(n_90), .Y(n_1188) );
INVx1_ASAP7_75t_L g749 ( .A(n_91), .Y(n_749) );
AOI22xp5_ASAP7_75t_SL g1446 ( .A1(n_92), .A2(n_208), .B1(n_1413), .B2(n_1417), .Y(n_1446) );
INVx1_ASAP7_75t_L g1072 ( .A(n_93), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g450 ( .A1(n_94), .A2(n_149), .B1(n_451), .B2(n_452), .Y(n_450) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_94), .A2(n_149), .B1(n_330), .B2(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g948 ( .A(n_95), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g1682 ( .A(n_96), .Y(n_1682) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_97), .A2(n_140), .B1(n_820), .B2(n_821), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_97), .A2(n_140), .B1(n_871), .B2(n_873), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g1387 ( .A1(n_98), .A2(n_105), .B1(n_791), .B2(n_1234), .Y(n_1387) );
OAI22xp33_ASAP7_75t_L g1396 ( .A1(n_98), .A2(n_105), .B1(n_871), .B2(n_1050), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_99), .A2(n_118), .B1(n_744), .B2(n_904), .Y(n_1157) );
INVx1_ASAP7_75t_L g359 ( .A(n_100), .Y(n_359) );
INVx1_ASAP7_75t_L g688 ( .A(n_101), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_101), .A2(n_231), .B1(n_711), .B2(n_712), .Y(n_710) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_102), .Y(n_571) );
INVx1_ASAP7_75t_L g321 ( .A(n_103), .Y(n_321) );
INVx1_ASAP7_75t_L g1011 ( .A(n_104), .Y(n_1011) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_106), .A2(n_164), .B1(n_524), .B2(n_1148), .Y(n_1147) );
OAI211xp5_ASAP7_75t_L g1227 ( .A1(n_107), .A2(n_1183), .B(n_1228), .C(n_1229), .Y(n_1227) );
INVx1_ASAP7_75t_L g1242 ( .A(n_107), .Y(n_1242) );
INVx1_ASAP7_75t_L g1182 ( .A(n_108), .Y(n_1182) );
OAI211xp5_ASAP7_75t_L g1186 ( .A1(n_108), .A2(n_446), .B(n_671), .C(n_1187), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g1137 ( .A(n_109), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1158 ( .A1(n_109), .A2(n_251), .B1(n_680), .B2(n_906), .Y(n_1158) );
AOI22xp5_ASAP7_75t_L g1442 ( .A1(n_110), .A2(n_294), .B1(n_1417), .B2(n_1423), .Y(n_1442) );
INVx1_ASAP7_75t_L g1338 ( .A(n_111), .Y(n_1338) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_113), .Y(n_915) );
INVx1_ASAP7_75t_L g388 ( .A(n_114), .Y(n_388) );
INVx1_ASAP7_75t_L g1335 ( .A(n_115), .Y(n_1335) );
INVx1_ASAP7_75t_L g1337 ( .A(n_116), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_117), .A2(n_128), .B1(n_509), .B2(n_1175), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g1360 ( .A1(n_117), .A2(n_128), .B1(n_1097), .B2(n_1237), .Y(n_1360) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_118), .A2(n_212), .B1(n_715), .B2(n_716), .C(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1263 ( .A(n_119), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_121), .A2(n_269), .B1(n_508), .B2(n_1175), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1397 ( .A1(n_121), .A2(n_269), .B1(n_472), .B2(n_879), .Y(n_1397) );
INVx1_ASAP7_75t_L g1391 ( .A(n_122), .Y(n_1391) );
INVx1_ASAP7_75t_L g1352 ( .A(n_123), .Y(n_1352) );
OAI211xp5_ASAP7_75t_L g1357 ( .A1(n_123), .A2(n_456), .B(n_1239), .C(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1327 ( .A(n_124), .Y(n_1327) );
INVx1_ASAP7_75t_L g1362 ( .A(n_125), .Y(n_1362) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_126), .A2(n_252), .B1(n_679), .B2(n_681), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g707 ( .A1(n_126), .A2(n_610), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g1074 ( .A(n_127), .Y(n_1074) );
OAI211xp5_ASAP7_75t_L g1090 ( .A1(n_129), .A2(n_671), .B(n_1091), .C(n_1093), .Y(n_1090) );
INVx1_ASAP7_75t_L g1106 ( .A(n_129), .Y(n_1106) );
AOI221xp5_ASAP7_75t_L g1118 ( .A1(n_130), .A2(n_251), .B1(n_1119), .B2(n_1120), .C(n_1122), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_130), .A2(n_216), .B1(n_968), .B2(n_1154), .Y(n_1153) );
OAI22xp5_ASAP7_75t_L g1232 ( .A1(n_131), .A2(n_299), .B1(n_508), .B2(n_510), .Y(n_1232) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_131), .A2(n_299), .B1(n_1190), .B2(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1082 ( .A(n_132), .Y(n_1082) );
INVx1_ASAP7_75t_L g366 ( .A(n_134), .Y(n_366) );
INVx1_ASAP7_75t_L g372 ( .A(n_135), .Y(n_372) );
OAI211xp5_ASAP7_75t_L g1301 ( .A1(n_136), .A2(n_1183), .B(n_1302), .C(n_1304), .Y(n_1301) );
INVx1_ASAP7_75t_L g1315 ( .A(n_136), .Y(n_1315) );
OAI22xp33_ASAP7_75t_L g1233 ( .A1(n_137), .A2(n_173), .B1(n_791), .B2(n_1234), .Y(n_1233) );
OAI22xp33_ASAP7_75t_L g1243 ( .A1(n_137), .A2(n_173), .B1(n_451), .B2(n_1050), .Y(n_1243) );
OAI22xp33_ASAP7_75t_L g1354 ( .A1(n_138), .A2(n_223), .B1(n_482), .B2(n_1234), .Y(n_1354) );
OAI22xp33_ASAP7_75t_L g1356 ( .A1(n_138), .A2(n_223), .B1(n_451), .B2(n_873), .Y(n_1356) );
INVx1_ASAP7_75t_L g843 ( .A(n_139), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g1680 ( .A(n_142), .Y(n_1680) );
OAI22xp33_ASAP7_75t_L g1700 ( .A1(n_143), .A2(n_186), .B1(n_791), .B2(n_1701), .Y(n_1700) );
OAI22xp33_ASAP7_75t_L g1713 ( .A1(n_143), .A2(n_175), .B1(n_471), .B2(n_474), .Y(n_1713) );
CKINVDCx5p33_ASAP7_75t_R g1673 ( .A(n_144), .Y(n_1673) );
INVx1_ASAP7_75t_L g764 ( .A(n_145), .Y(n_764) );
INVx1_ASAP7_75t_L g756 ( .A(n_146), .Y(n_756) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_147), .A2(n_232), .B1(n_1049), .B2(n_1050), .Y(n_1048) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_147), .A2(n_232), .B1(n_821), .B2(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1374 ( .A(n_148), .Y(n_1374) );
INVx1_ASAP7_75t_L g1181 ( .A(n_150), .Y(n_1181) );
INVx1_ASAP7_75t_L g1008 ( .A(n_151), .Y(n_1008) );
INVx1_ASAP7_75t_L g1018 ( .A(n_152), .Y(n_1018) );
INVxp67_ASAP7_75t_SL g1658 ( .A(n_153), .Y(n_1658) );
INVx1_ASAP7_75t_L g465 ( .A(n_154), .Y(n_465) );
INVx1_ASAP7_75t_L g1079 ( .A(n_155), .Y(n_1079) );
INVx1_ASAP7_75t_L g758 ( .A(n_157), .Y(n_758) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_158), .A2(n_302), .B1(n_452), .B2(n_781), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g790 ( .A1(n_158), .A2(n_302), .B1(n_330), .B2(n_791), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_159), .A2(n_183), .B1(n_788), .B2(n_880), .Y(n_1041) );
OAI22xp33_ASAP7_75t_L g1054 ( .A1(n_159), .A2(n_183), .B1(n_1055), .B2(n_1057), .Y(n_1054) );
OAI211xp5_ASAP7_75t_L g1388 ( .A1(n_160), .A2(n_863), .B(n_1389), .C(n_1390), .Y(n_1388) );
INVx1_ASAP7_75t_L g1401 ( .A(n_160), .Y(n_1401) );
INVx1_ASAP7_75t_L g1698 ( .A(n_161), .Y(n_1698) );
OAI211xp5_ASAP7_75t_L g1706 ( .A1(n_161), .A2(n_456), .B(n_1707), .C(n_1709), .Y(n_1706) );
INVx1_ASAP7_75t_L g747 ( .A(n_162), .Y(n_747) );
INVx1_ASAP7_75t_L g379 ( .A(n_163), .Y(n_379) );
OAI211xp5_ASAP7_75t_L g1114 ( .A1(n_164), .A2(n_1115), .B(n_1117), .C(n_1125), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g580 ( .A1(n_165), .A2(n_300), .B1(n_581), .B2(n_583), .C(n_585), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_165), .A2(n_311), .B1(n_639), .B2(n_640), .Y(n_638) );
INVxp67_ASAP7_75t_SL g974 ( .A(n_166), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_167), .A2(n_252), .B1(n_711), .B2(n_712), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g1694 ( .A1(n_168), .A2(n_1179), .B(n_1389), .C(n_1695), .Y(n_1694) );
INVx1_ASAP7_75t_L g1712 ( .A(n_168), .Y(n_1712) );
INVx1_ASAP7_75t_L g1479 ( .A(n_169), .Y(n_1479) );
AOI22xp5_ASAP7_75t_SL g1412 ( .A1(n_170), .A2(n_179), .B1(n_1413), .B2(n_1417), .Y(n_1412) );
INVx1_ASAP7_75t_L g1256 ( .A(n_171), .Y(n_1256) );
INVx1_ASAP7_75t_L g1231 ( .A(n_172), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1238 ( .A1(n_172), .A2(n_456), .B(n_1239), .C(n_1241), .Y(n_1238) );
OAI22xp33_ASAP7_75t_L g1699 ( .A1(n_174), .A2(n_175), .B1(n_1059), .B2(n_1234), .Y(n_1699) );
OAI22xp33_ASAP7_75t_L g1703 ( .A1(n_174), .A2(n_186), .B1(n_451), .B2(n_1704), .Y(n_1703) );
OAI22xp33_ASAP7_75t_L g1096 ( .A1(n_176), .A2(n_304), .B1(n_880), .B2(n_1097), .Y(n_1096) );
OAI22xp33_ASAP7_75t_L g1103 ( .A1(n_176), .A2(n_304), .B1(n_1055), .B2(n_1057), .Y(n_1103) );
INVx1_ASAP7_75t_L g1638 ( .A(n_177), .Y(n_1638) );
AOI221x1_ASAP7_75t_SL g1650 ( .A1(n_177), .A2(n_236), .B1(n_744), .B2(n_900), .C(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1367 ( .A(n_178), .Y(n_1367) );
INVx1_ASAP7_75t_L g1126 ( .A(n_180), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g1164 ( .A1(n_180), .A2(n_277), .B1(n_1165), .B2(n_1166), .Y(n_1164) );
AOI21xp33_ASAP7_75t_L g1644 ( .A1(n_181), .A2(n_609), .B(n_610), .Y(n_1644) );
INVx1_ASAP7_75t_L g1659 ( .A(n_181), .Y(n_1659) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_182), .A2(n_234), .B1(n_1130), .B2(n_1133), .C(n_1134), .Y(n_1129) );
INVx1_ASAP7_75t_L g1160 ( .A(n_182), .Y(n_1160) );
INVx2_ASAP7_75t_L g1416 ( .A(n_184), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_184), .B(n_272), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_184), .B(n_1422), .Y(n_1424) );
AOI22xp5_ASAP7_75t_SL g1427 ( .A1(n_185), .A2(n_233), .B1(n_1423), .B2(n_1428), .Y(n_1427) );
CKINVDCx5p33_ASAP7_75t_R g1677 ( .A(n_187), .Y(n_1677) );
INVx1_ASAP7_75t_L g816 ( .A(n_188), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_190), .A2(n_291), .B1(n_1413), .B2(n_1428), .Y(n_1434) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_191), .A2(n_520), .B1(n_648), .B2(n_649), .Y(n_519) );
INVxp67_ASAP7_75t_L g649 ( .A(n_191), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g1437 ( .A1(n_192), .A2(n_235), .B1(n_1420), .B2(n_1423), .Y(n_1437) );
OAI211xp5_ASAP7_75t_L g810 ( .A1(n_193), .A2(n_811), .B(n_812), .C(n_813), .Y(n_810) );
INVx1_ASAP7_75t_L g877 ( .A(n_193), .Y(n_877) );
XOR2x2_ASAP7_75t_L g1168 ( .A(n_195), .B(n_1169), .Y(n_1168) );
INVx1_ASAP7_75t_L g468 ( .A(n_196), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g488 ( .A1(n_196), .A2(n_489), .B(n_491), .C(n_497), .Y(n_488) );
XOR2x2_ASAP7_75t_L g1274 ( .A(n_197), .B(n_1275), .Y(n_1274) );
AOI22xp5_ASAP7_75t_L g1443 ( .A1(n_198), .A2(n_253), .B1(n_1413), .B2(n_1420), .Y(n_1443) );
OAI221xp5_ASAP7_75t_SL g557 ( .A1(n_199), .A2(n_267), .B1(n_558), .B2(n_564), .C(n_570), .Y(n_557) );
INVx1_ASAP7_75t_L g600 ( .A(n_199), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_200), .A2(n_279), .B1(n_744), .B2(n_904), .Y(n_955) );
INVx1_ASAP7_75t_L g942 ( .A(n_202), .Y(n_942) );
INVx2_ASAP7_75t_L g404 ( .A(n_203), .Y(n_404) );
INVx1_ASAP7_75t_L g444 ( .A(n_203), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_203), .B(n_405), .Y(n_547) );
INVx1_ASAP7_75t_L g751 ( .A(n_204), .Y(n_751) );
INVx1_ASAP7_75t_L g1378 ( .A(n_205), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1307 ( .A1(n_206), .A2(n_210), .B1(n_800), .B2(n_1308), .Y(n_1307) );
OAI22xp33_ASAP7_75t_L g1316 ( .A1(n_206), .A2(n_210), .B1(n_1097), .B2(n_1317), .Y(n_1316) );
CKINVDCx5p33_ASAP7_75t_R g1284 ( .A(n_207), .Y(n_1284) );
INVx1_ASAP7_75t_L g1372 ( .A(n_209), .Y(n_1372) );
BUFx3_ASAP7_75t_L g411 ( .A(n_211), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g1685 ( .A(n_213), .Y(n_1685) );
INVx1_ASAP7_75t_L g532 ( .A(n_214), .Y(n_532) );
INVx1_ASAP7_75t_L g1095 ( .A(n_215), .Y(n_1095) );
OAI211xp5_ASAP7_75t_L g1104 ( .A1(n_215), .A2(n_793), .B(n_812), .C(n_1105), .Y(n_1104) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_216), .Y(n_1135) );
AOI22xp5_ASAP7_75t_L g1433 ( .A1(n_217), .A2(n_246), .B1(n_1420), .B2(n_1423), .Y(n_1433) );
OAI22xp5_ASAP7_75t_SL g1629 ( .A1(n_218), .A2(n_254), .B1(n_573), .B2(n_577), .Y(n_1629) );
CKINVDCx5p33_ASAP7_75t_R g1636 ( .A(n_218), .Y(n_1636) );
INVx1_ASAP7_75t_L g994 ( .A(n_219), .Y(n_994) );
INVx1_ASAP7_75t_L g1250 ( .A(n_220), .Y(n_1250) );
CKINVDCx5p33_ASAP7_75t_R g1280 ( .A(n_221), .Y(n_1280) );
CKINVDCx5p33_ASAP7_75t_R g1676 ( .A(n_222), .Y(n_1676) );
INVx1_ASAP7_75t_L g1200 ( .A(n_224), .Y(n_1200) );
INVx1_ASAP7_75t_L g836 ( .A(n_225), .Y(n_836) );
INVx1_ASAP7_75t_L g662 ( .A(n_226), .Y(n_662) );
INVx1_ASAP7_75t_L g1021 ( .A(n_227), .Y(n_1021) );
XNOR2xp5_ASAP7_75t_L g1617 ( .A(n_228), .B(n_1618), .Y(n_1617) );
BUFx3_ASAP7_75t_L g338 ( .A(n_229), .Y(n_338) );
INVx1_ASAP7_75t_L g485 ( .A(n_229), .Y(n_485) );
OAI22xp33_ASAP7_75t_L g469 ( .A1(n_230), .A2(n_276), .B1(n_470), .B2(n_472), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_230), .A2(n_276), .B1(n_508), .B2(n_510), .Y(n_507) );
INVx1_ASAP7_75t_L g677 ( .A(n_231), .Y(n_677) );
XNOR2xp5_ASAP7_75t_L g1320 ( .A(n_233), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1162 ( .A(n_234), .Y(n_1162) );
AOI22xp33_ASAP7_75t_L g1645 ( .A1(n_236), .A2(n_241), .B1(n_590), .B2(n_612), .Y(n_1645) );
INVx1_ASAP7_75t_L g1331 ( .A(n_237), .Y(n_1331) );
INVx1_ASAP7_75t_L g1206 ( .A(n_238), .Y(n_1206) );
INVx1_ASAP7_75t_L g607 ( .A(n_239), .Y(n_607) );
INVx1_ASAP7_75t_L g817 ( .A(n_240), .Y(n_817) );
OAI211xp5_ASAP7_75t_L g874 ( .A1(n_240), .A2(n_671), .B(n_752), .C(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g1252 ( .A(n_242), .Y(n_1252) );
CKINVDCx5p33_ASAP7_75t_R g1287 ( .A(n_243), .Y(n_1287) );
INVx1_ASAP7_75t_L g844 ( .A(n_244), .Y(n_844) );
INVx1_ASAP7_75t_L g1205 ( .A(n_245), .Y(n_1205) );
INVx1_ASAP7_75t_L g383 ( .A(n_247), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_249), .Y(n_916) );
CKINVDCx5p33_ASAP7_75t_R g1674 ( .A(n_250), .Y(n_1674) );
INVx1_ASAP7_75t_L g1633 ( .A(n_254), .Y(n_1633) );
INVx1_ASAP7_75t_L g1202 ( .A(n_255), .Y(n_1202) );
INVx1_ASAP7_75t_L g413 ( .A(n_256), .Y(n_413) );
INVx1_ASAP7_75t_L g419 ( .A(n_256), .Y(n_419) );
INVx1_ASAP7_75t_L g786 ( .A(n_257), .Y(n_786) );
OAI211xp5_ASAP7_75t_L g792 ( .A1(n_257), .A2(n_793), .B(n_795), .C(n_797), .Y(n_792) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_258), .A2(n_651), .B1(n_652), .B2(n_732), .Y(n_650) );
INVxp67_ASAP7_75t_L g732 ( .A(n_258), .Y(n_732) );
INVx1_ASAP7_75t_L g1077 ( .A(n_259), .Y(n_1077) );
INVx1_ASAP7_75t_L g1209 ( .A(n_260), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g1305 ( .A(n_261), .Y(n_1305) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_262), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_262), .A2(n_301), .B1(n_720), .B2(n_721), .C(n_724), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g1282 ( .A(n_263), .Y(n_1282) );
INVx1_ASAP7_75t_L g389 ( .A(n_264), .Y(n_389) );
INVx1_ASAP7_75t_L g1643 ( .A(n_265), .Y(n_1643) );
INVx1_ASAP7_75t_L g1046 ( .A(n_266), .Y(n_1046) );
INVx1_ASAP7_75t_L g618 ( .A(n_267), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g664 ( .A(n_268), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_270), .A2(n_807), .B1(n_808), .B2(n_882), .Y(n_806) );
INVxp67_ASAP7_75t_SL g882 ( .A(n_270), .Y(n_882) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_271), .Y(n_911) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_272), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1422 ( .A(n_272), .Y(n_1422) );
OAI211xp5_ASAP7_75t_SL g1042 ( .A1(n_273), .A2(n_671), .B(n_1043), .C(n_1045), .Y(n_1042) );
INVx1_ASAP7_75t_L g1064 ( .A(n_273), .Y(n_1064) );
CKINVDCx5p33_ASAP7_75t_R g1289 ( .A(n_274), .Y(n_1289) );
INVx1_ASAP7_75t_L g893 ( .A(n_275), .Y(n_893) );
INVx1_ASAP7_75t_L g1127 ( .A(n_277), .Y(n_1127) );
INVx1_ASAP7_75t_L g1248 ( .A(n_278), .Y(n_1248) );
INVx1_ASAP7_75t_L g982 ( .A(n_279), .Y(n_982) );
INVx1_ASAP7_75t_L g669 ( .A(n_280), .Y(n_669) );
INVx1_ASAP7_75t_L g1306 ( .A(n_281), .Y(n_1306) );
OAI211xp5_ASAP7_75t_L g1311 ( .A1(n_281), .A2(n_456), .B(n_1312), .C(n_1314), .Y(n_1311) );
INVx1_ASAP7_75t_L g762 ( .A(n_282), .Y(n_762) );
INVx1_ASAP7_75t_L g1481 ( .A(n_283), .Y(n_1481) );
CKINVDCx5p33_ASAP7_75t_R g1697 ( .A(n_284), .Y(n_1697) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_285), .Y(n_686) );
INVx1_ASAP7_75t_L g1208 ( .A(n_286), .Y(n_1208) );
AOI211xp5_ASAP7_75t_SL g936 ( .A1(n_288), .A2(n_937), .B(n_938), .C(n_941), .Y(n_936) );
INVx1_ASAP7_75t_L g1375 ( .A(n_289), .Y(n_1375) );
INVx1_ASAP7_75t_L g981 ( .A(n_290), .Y(n_981) );
XNOR2xp5_ASAP7_75t_L g1066 ( .A(n_291), .B(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1081 ( .A(n_292), .Y(n_1081) );
INVx1_ASAP7_75t_L g356 ( .A(n_293), .Y(n_356) );
XOR2x2_ASAP7_75t_L g345 ( .A(n_294), .B(n_346), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g1279 ( .A(n_295), .Y(n_1279) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
INVx1_ASAP7_75t_L g831 ( .A(n_297), .Y(n_831) );
INVx1_ASAP7_75t_L g850 ( .A(n_298), .Y(n_850) );
INVx1_ASAP7_75t_L g626 ( .A(n_300), .Y(n_626) );
INVx1_ASAP7_75t_L g659 ( .A(n_301), .Y(n_659) );
INVx1_ASAP7_75t_L g1262 ( .A(n_305), .Y(n_1262) );
INVx1_ASAP7_75t_L g1203 ( .A(n_306), .Y(n_1203) );
INVx2_ASAP7_75t_L g353 ( .A(n_307), .Y(n_353) );
INVx1_ASAP7_75t_L g399 ( .A(n_307), .Y(n_399) );
INVx1_ASAP7_75t_L g443 ( .A(n_307), .Y(n_443) );
INVx1_ASAP7_75t_L g1628 ( .A(n_309), .Y(n_1628) );
CKINVDCx5p33_ASAP7_75t_R g894 ( .A(n_310), .Y(n_894) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_339), .B(n_1405), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx4f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_324), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g1717 ( .A(n_318), .B(n_327), .Y(n_1717) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g1664 ( .A(n_320), .B(n_323), .Y(n_1664) );
INVx1_ASAP7_75t_L g1720 ( .A(n_320), .Y(n_1720) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g1723 ( .A(n_323), .B(n_1720), .Y(n_1723) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g514 ( .A(n_327), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g394 ( .A(n_328), .B(n_338), .Y(n_394) );
AND2x4_ASAP7_75t_L g586 ( .A(n_328), .B(n_337), .Y(n_586) );
INVx1_ASAP7_75t_L g820 ( .A(n_329), .Y(n_820) );
INVxp67_ASAP7_75t_SL g1053 ( .A(n_329), .Y(n_1053) );
AND2x4_ASAP7_75t_SL g1716 ( .A(n_329), .B(n_1717), .Y(n_1716) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x6_ASAP7_75t_L g330 ( .A(n_331), .B(n_336), .Y(n_330) );
INVxp67_ASAP7_75t_L g358 ( .A(n_331), .Y(n_358) );
OR2x6_ASAP7_75t_L g509 ( .A(n_331), .B(n_484), .Y(n_509) );
BUFx4f_ASAP7_75t_L g767 ( .A(n_331), .Y(n_767) );
INVx1_ASAP7_75t_L g1037 ( .A(n_331), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1701 ( .A(n_331), .B(n_484), .Y(n_1701) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx3_ASAP7_75t_L g387 ( .A(n_332), .Y(n_387) );
BUFx4f_ASAP7_75t_L g856 ( .A(n_332), .Y(n_856) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
INVx2_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
INVx2_ASAP7_75t_L g371 ( .A(n_334), .Y(n_371) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_334), .B(n_335), .Y(n_375) );
AND2x2_ASAP7_75t_L g486 ( .A(n_334), .B(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g496 ( .A(n_334), .B(n_335), .Y(n_496) );
INVx1_ASAP7_75t_L g505 ( .A(n_334), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_335), .B(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g370 ( .A(n_335), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g487 ( .A(n_335), .Y(n_487) );
BUFx2_ASAP7_75t_L g500 ( .A(n_335), .Y(n_500) );
INVx1_ASAP7_75t_L g540 ( .A(n_335), .Y(n_540) );
AND2x2_ASAP7_75t_L g591 ( .A(n_335), .B(n_364), .Y(n_591) );
OR2x6_ASAP7_75t_L g1234 ( .A(n_336), .B(n_387), .Y(n_1234) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g493 ( .A(n_337), .Y(n_493) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g499 ( .A(n_338), .Y(n_499) );
AND2x4_ASAP7_75t_L g503 ( .A(n_338), .B(n_504), .Y(n_503) );
XNOR2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_1107), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_801), .B2(n_802), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AO22x2_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_734), .B2(n_735), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AO22x2_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_517), .B1(n_518), .B2(n_733), .Y(n_344) );
INVx1_ASAP7_75t_L g733 ( .A(n_345), .Y(n_733) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_449), .C(n_480), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_400), .Y(n_347) );
OAI33xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_355), .A3(n_365), .B1(n_376), .B2(n_384), .B3(n_392), .Y(n_348) );
OAI33xp33_ASAP7_75t_L g1291 ( .A1(n_349), .A2(n_392), .A3(n_1292), .B1(n_1293), .B2(n_1294), .B3(n_1297), .Y(n_1291) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI33xp33_ASAP7_75t_L g1671 ( .A1(n_350), .A2(n_1259), .A3(n_1672), .B1(n_1675), .B2(n_1678), .B3(n_1681), .Y(n_1671) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g769 ( .A(n_351), .Y(n_769) );
INVx1_ASAP7_75t_L g1024 ( .A(n_351), .Y(n_1024) );
INVx2_ASAP7_75t_L g1194 ( .A(n_351), .Y(n_1194) );
INVx4_ASAP7_75t_L g1342 ( .A(n_351), .Y(n_1342) );
INVx2_ASAP7_75t_L g1382 ( .A(n_351), .Y(n_1382) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
INVx1_ASAP7_75t_L g622 ( .A(n_352), .Y(n_622) );
OR2x6_ASAP7_75t_L g908 ( .A(n_352), .B(n_909), .Y(n_908) );
OR2x2_ASAP7_75t_L g1692 ( .A(n_352), .B(n_909), .Y(n_1692) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g731 ( .A(n_353), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B1(n_359), .B2(n_360), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_356), .A2(n_379), .B1(n_407), .B2(n_414), .Y(n_406) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g445 ( .A1(n_359), .A2(n_383), .B1(n_407), .B2(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g1672 ( .A1(n_360), .A2(n_943), .B1(n_1673), .B2(n_1674), .Y(n_1672) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
INVx1_ASAP7_75t_L g768 ( .A(n_361), .Y(n_768) );
INVx4_ASAP7_75t_L g859 ( .A(n_361), .Y(n_859) );
INVx2_ASAP7_75t_L g986 ( .A(n_361), .Y(n_986) );
INVx1_ASAP7_75t_L g1039 ( .A(n_361), .Y(n_1039) );
INVx2_ASAP7_75t_L g1298 ( .A(n_361), .Y(n_1298) );
INVx2_ASAP7_75t_L g1684 ( .A(n_361), .Y(n_1684) );
INVx8_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g512 ( .A(n_362), .B(n_499), .Y(n_512) );
BUFx2_ASAP7_75t_L g1136 ( .A(n_362), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_372), .B2(n_373), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_366), .A2(n_388), .B1(n_422), .B2(n_428), .Y(n_421) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx4_ASAP7_75t_L g771 ( .A(n_368), .Y(n_771) );
INVx2_ASAP7_75t_L g773 ( .A(n_368), .Y(n_773) );
INVx2_ASAP7_75t_L g1087 ( .A(n_368), .Y(n_1087) );
INVx4_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g378 ( .A(n_370), .Y(n_378) );
INVx2_ASAP7_75t_L g862 ( .A(n_370), .Y(n_862) );
BUFx3_ASAP7_75t_L g940 ( .A(n_370), .Y(n_940) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_370), .Y(n_1253) );
AND2x2_ASAP7_75t_L g539 ( .A(n_371), .B(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_371), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_372), .A2(n_389), .B1(n_433), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g794 ( .A(n_373), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g1381 ( .A1(n_373), .A2(n_1253), .B1(n_1371), .B2(n_1374), .Y(n_1381) );
BUFx4f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx4_ASAP7_75t_L g490 ( .A(n_374), .Y(n_490) );
BUFx4f_ASAP7_75t_L g811 ( .A(n_374), .Y(n_811) );
BUFx4f_ASAP7_75t_L g863 ( .A(n_374), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g993 ( .A1(n_374), .A2(n_394), .B1(n_940), .B2(n_994), .C(n_995), .Y(n_993) );
BUFx6f_ASAP7_75t_L g1228 ( .A(n_374), .Y(n_1228) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx3_ASAP7_75t_L g382 ( .A(n_375), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B1(n_380), .B2(n_383), .Y(n_376) );
OAI22xp5_ASAP7_75t_SL g1293 ( .A1(n_377), .A2(n_1228), .B1(n_1282), .B2(n_1286), .Y(n_1293) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI211xp5_ASAP7_75t_L g606 ( .A1(n_380), .A2(n_607), .B(n_608), .C(n_611), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_380), .A2(n_742), .B1(n_762), .B2(n_771), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_380), .A2(n_1011), .B1(n_1014), .B2(n_1029), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g1031 ( .A1(n_380), .A2(n_1008), .B1(n_1022), .B2(n_1032), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_380), .A2(n_1072), .B1(n_1082), .B2(n_1087), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1204 ( .A1(n_380), .A2(n_861), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
INVx5_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g706 ( .A(n_382), .Y(n_706) );
BUFx2_ASAP7_75t_SL g774 ( .A(n_382), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_382), .B(n_935), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_382), .B(n_989), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g1675 ( .A1(n_382), .A2(n_925), .B1(n_1676), .B2(n_1677), .Y(n_1675) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_389), .B2(n_390), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g1134 ( .A1(n_385), .A2(n_1135), .B1(n_1136), .B2(n_1137), .C(n_1138), .Y(n_1134) );
OAI22xp33_ASAP7_75t_L g1292 ( .A1(n_385), .A2(n_390), .B1(n_1279), .B2(n_1289), .Y(n_1292) );
OAI22xp33_ASAP7_75t_L g1297 ( .A1(n_385), .A2(n_1284), .B1(n_1287), .B2(n_1298), .Y(n_1297) );
OAI22xp33_ASAP7_75t_L g1343 ( .A1(n_385), .A2(n_859), .B1(n_1325), .B2(n_1337), .Y(n_1343) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
BUFx3_ASAP7_75t_L g776 ( .A(n_387), .Y(n_776) );
BUFx3_ASAP7_75t_L g1199 ( .A(n_387), .Y(n_1199) );
BUFx6f_ASAP7_75t_L g1249 ( .A(n_387), .Y(n_1249) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_390), .A2(n_1034), .B1(n_1075), .B2(n_1079), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g1261 ( .A1(n_390), .A2(n_767), .B1(n_1262), .B2(n_1263), .Y(n_1261) );
INVx5_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx6_ASAP7_75t_L g777 ( .A(n_391), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g778 ( .A(n_393), .Y(n_778) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx4_ASAP7_75t_L g610 ( .A(n_394), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_394), .B(n_395), .Y(n_867) );
OAI21xp33_ASAP7_75t_L g938 ( .A1(n_394), .A2(n_939), .B(n_940), .Y(n_938) );
INVx1_ASAP7_75t_SL g1122 ( .A(n_394), .Y(n_1122) );
AND2x2_ASAP7_75t_SL g1260 ( .A(n_394), .B(n_397), .Y(n_1260) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g402 ( .A(n_397), .B(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_397), .Y(n_479) );
OR2x2_ASAP7_75t_L g546 ( .A(n_397), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx2_ASAP7_75t_L g516 ( .A(n_398), .Y(n_516) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI33xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_406), .A3(n_421), .B1(n_432), .B2(n_440), .B3(n_445), .Y(n_400) );
OAI33xp33_ASAP7_75t_L g1277 ( .A1(n_401), .A2(n_759), .A3(n_1278), .B1(n_1281), .B2(n_1285), .B3(n_1288), .Y(n_1277) );
BUFx8_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx4f_ASAP7_75t_L g633 ( .A(n_402), .Y(n_633) );
BUFx4f_ASAP7_75t_L g683 ( .A(n_402), .Y(n_683) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_402), .Y(n_1265) );
NAND2xp33_ASAP7_75t_SL g403 ( .A(n_404), .B(n_405), .Y(n_403) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_404), .Y(n_477) );
INVx1_ASAP7_75t_L g529 ( .A(n_404), .Y(n_529) );
AND3x4_ASAP7_75t_L g896 ( .A(n_404), .B(n_463), .C(n_731), .Y(n_896) );
INVx3_ASAP7_75t_L g441 ( .A(n_405), .Y(n_441) );
BUFx3_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
OAI22xp33_ASAP7_75t_L g1278 ( .A1(n_407), .A2(n_752), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g1007 ( .A(n_409), .Y(n_1007) );
BUFx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OR2x4_ASAP7_75t_L g451 ( .A(n_410), .B(n_441), .Y(n_451) );
OR2x4_ASAP7_75t_L g471 ( .A(n_410), .B(n_454), .Y(n_471) );
INVx2_ASAP7_75t_L g543 ( .A(n_410), .Y(n_543) );
BUFx3_ASAP7_75t_L g757 ( .A(n_410), .Y(n_757) );
BUFx4f_ASAP7_75t_L g1214 ( .A(n_410), .Y(n_1214) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_411), .Y(n_420) );
INVx2_ASAP7_75t_L g427 ( .A(n_411), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_411), .B(n_419), .Y(n_431) );
AND2x4_ASAP7_75t_L g458 ( .A(n_411), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g527 ( .A(n_412), .Y(n_527) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVxp67_ASAP7_75t_L g426 ( .A(n_413), .Y(n_426) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVxp67_ASAP7_75t_SL g1092 ( .A(n_415), .Y(n_1092) );
INVxp67_ASAP7_75t_SL g1379 ( .A(n_415), .Y(n_1379) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g1044 ( .A(n_416), .Y(n_1044) );
INVx1_ASAP7_75t_L g1708 ( .A(n_416), .Y(n_1708) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_417), .Y(n_448) );
BUFx3_ASAP7_75t_L g754 ( .A(n_417), .Y(n_754) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
BUFx2_ASAP7_75t_L g467 ( .A(n_418), .Y(n_467) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
BUFx2_ASAP7_75t_L g464 ( .A(n_420), .Y(n_464) );
INVx2_ASAP7_75t_L g563 ( .A(n_420), .Y(n_563) );
AND2x4_ASAP7_75t_L g641 ( .A(n_420), .B(n_569), .Y(n_641) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g551 ( .A(n_423), .B(n_545), .Y(n_551) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g639 ( .A(n_424), .Y(n_639) );
BUFx2_ASAP7_75t_L g685 ( .A(n_424), .Y(n_685) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_425), .Y(n_435) );
BUFx6f_ASAP7_75t_L g746 ( .A(n_425), .Y(n_746) );
BUFx8_ASAP7_75t_L g842 ( .A(n_425), .Y(n_842) );
AND2x4_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
AND2x4_ASAP7_75t_L g526 ( .A(n_427), .B(n_527), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_428), .A2(n_675), .B1(n_676), .B2(n_677), .C(n_678), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g1285 ( .A1(n_428), .A2(n_761), .B1(n_1286), .B2(n_1287), .Y(n_1285) );
CKINVDCx8_ASAP7_75t_R g428 ( .A(n_429), .Y(n_428) );
INVx3_ASAP7_75t_L g687 ( .A(n_429), .Y(n_687) );
INVx3_ASAP7_75t_L g839 ( .A(n_429), .Y(n_839) );
INVx3_ASAP7_75t_L g1019 ( .A(n_429), .Y(n_1019) );
INVx1_ASAP7_75t_L g1270 ( .A(n_429), .Y(n_1270) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g574 ( .A(n_430), .Y(n_574) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g439 ( .A(n_431), .Y(n_439) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g453 ( .A(n_435), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g625 ( .A(n_435), .Y(n_625) );
INVx1_ASAP7_75t_L g1283 ( .A(n_435), .Y(n_1283) );
INVx2_ASAP7_75t_L g1689 ( .A(n_435), .Y(n_1689) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_435), .B(n_454), .Y(n_1705) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_436), .A2(n_625), .B1(n_626), .B2(n_627), .C(n_628), .Y(n_624) );
OAI22xp33_ASAP7_75t_SL g741 ( .A1(n_436), .A2(n_742), .B1(n_743), .B2(n_747), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g1281 ( .A1(n_436), .A2(n_1282), .B1(n_1283), .B2(n_1284), .Y(n_1281) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x6_ASAP7_75t_L g474 ( .A(n_439), .B(n_441), .Y(n_474) );
BUFx3_ASAP7_75t_L g763 ( .A(n_439), .Y(n_763) );
INVx3_ASAP7_75t_L g647 ( .A(n_440), .Y(n_647) );
INVx3_ASAP7_75t_L g847 ( .A(n_440), .Y(n_847) );
NAND3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .C(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g454 ( .A(n_441), .Y(n_454) );
AND2x4_ASAP7_75t_L g457 ( .A(n_441), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g528 ( .A(n_441), .B(n_529), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g909 ( .A(n_441), .B(n_444), .Y(n_909) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g561 ( .A(n_443), .Y(n_561) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g1240 ( .A(n_447), .Y(n_1240) );
INVx1_ASAP7_75t_L g1313 ( .A(n_447), .Y(n_1313) );
INVx2_ASAP7_75t_L g1653 ( .A(n_447), .Y(n_1653) );
INVx4_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OR2x2_ASAP7_75t_L g577 ( .A(n_448), .B(n_546), .Y(n_577) );
BUFx6f_ASAP7_75t_L g834 ( .A(n_448), .Y(n_834) );
INVx3_ASAP7_75t_L g1268 ( .A(n_448), .Y(n_1268) );
OAI31xp33_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_455), .A3(n_469), .B(n_475), .Y(n_449) );
INVx2_ASAP7_75t_SL g668 ( .A(n_451), .Y(n_668) );
INVx1_ASAP7_75t_L g782 ( .A(n_451), .Y(n_782) );
INVx2_ASAP7_75t_SL g872 ( .A(n_451), .Y(n_872) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_451), .Y(n_1099) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_453), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
INVx2_ASAP7_75t_L g873 ( .A(n_453), .Y(n_873) );
INVx1_ASAP7_75t_L g1050 ( .A(n_453), .Y(n_1050) );
INVx1_ASAP7_75t_L g1100 ( .A(n_453), .Y(n_1100) );
CKINVDCx8_ASAP7_75t_R g456 ( .A(n_457), .Y(n_456) );
CKINVDCx8_ASAP7_75t_R g671 ( .A(n_457), .Y(n_671) );
BUFx2_ASAP7_75t_L g632 ( .A(n_458), .Y(n_632) );
BUFx2_ASAP7_75t_L g636 ( .A(n_458), .Y(n_636) );
INVx2_ASAP7_75t_L g646 ( .A(n_458), .Y(n_646) );
BUFx2_ASAP7_75t_L g665 ( .A(n_458), .Y(n_665) );
BUFx2_ASAP7_75t_L g968 ( .A(n_458), .Y(n_968) );
INVx1_ASAP7_75t_L g569 ( .A(n_459), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_465), .B1(n_466), .B2(n_468), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g1241 ( .A1(n_461), .A2(n_466), .B1(n_1230), .B2(n_1242), .Y(n_1241) );
AOI22xp33_ASAP7_75t_SL g1314 ( .A1(n_461), .A2(n_466), .B1(n_1305), .B2(n_1315), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_461), .A2(n_466), .B1(n_1350), .B2(n_1359), .Y(n_1358) );
AOI22xp33_ASAP7_75t_SL g1400 ( .A1(n_461), .A2(n_466), .B1(n_1391), .B2(n_1401), .Y(n_1400) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
AND2x4_ASAP7_75t_L g466 ( .A(n_462), .B(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g661 ( .A(n_462), .B(n_464), .Y(n_661) );
AND2x4_ASAP7_75t_L g1710 ( .A(n_462), .B(n_464), .Y(n_1710) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_462), .B(n_467), .Y(n_1711) );
INVx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_465), .A2(n_498), .B1(n_501), .B2(n_506), .Y(n_497) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_466), .Y(n_663) );
BUFx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_SL g670 ( .A(n_471), .Y(n_670) );
BUFx2_ASAP7_75t_L g788 ( .A(n_471), .Y(n_788) );
BUFx2_ASAP7_75t_L g1190 ( .A(n_471), .Y(n_1190) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g657 ( .A(n_474), .Y(n_657) );
BUFx3_ASAP7_75t_L g880 ( .A(n_474), .Y(n_880) );
INVx1_ASAP7_75t_L g1318 ( .A(n_474), .Y(n_1318) );
OAI31xp33_ASAP7_75t_L g779 ( .A1(n_475), .A2(n_780), .A3(n_783), .B(n_787), .Y(n_779) );
OAI31xp33_ASAP7_75t_L g1040 ( .A1(n_475), .A2(n_1041), .A3(n_1042), .B(n_1048), .Y(n_1040) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
AND2x4_ASAP7_75t_L g672 ( .A(n_476), .B(n_478), .Y(n_672) );
AND2x2_ASAP7_75t_SL g881 ( .A(n_476), .B(n_478), .Y(n_881) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_476), .B(n_478), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1714 ( .A(n_476), .B(n_478), .Y(n_1714) );
INVx1_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI31xp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_488), .A3(n_507), .B(n_513), .Y(n_480) );
INVx4_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g791 ( .A(n_483), .Y(n_791) );
INVx3_ASAP7_75t_SL g821 ( .A(n_483), .Y(n_821) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_486), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_486), .Y(n_555) );
INVx2_ASAP7_75t_L g709 ( .A(n_486), .Y(n_709) );
BUFx3_ASAP7_75t_L g1640 ( .A(n_486), .Y(n_1640) );
OAI22xp5_ASAP7_75t_SL g1251 ( .A1(n_489), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1251) );
NAND2xp5_ASAP7_75t_SL g1634 ( .A(n_489), .B(n_1635), .Y(n_1634) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g922 ( .A(n_490), .Y(n_922) );
INVx1_ASAP7_75t_L g1179 ( .A(n_490), .Y(n_1179) );
INVx2_ASAP7_75t_L g1257 ( .A(n_490), .Y(n_1257) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g1389 ( .A(n_492), .Y(n_1389) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x2_ASAP7_75t_L g796 ( .A(n_493), .B(n_584), .Y(n_796) );
AND2x2_ASAP7_75t_L g1696 ( .A(n_493), .B(n_500), .Y(n_1696) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g602 ( .A(n_495), .Y(n_602) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_496), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_498), .A2(n_501), .B1(n_785), .B2(n_798), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_498), .A2(n_1062), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_498), .A2(n_1350), .B1(n_1351), .B2(n_1352), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_498), .A2(n_1351), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
AND2x4_ASAP7_75t_L g815 ( .A(n_499), .B(n_500), .Y(n_815) );
INVx1_ASAP7_75t_L g599 ( .A(n_500), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_500), .A2(n_596), .B1(n_889), .B2(n_915), .Y(n_935) );
BUFx2_ASAP7_75t_L g990 ( .A(n_500), .Y(n_990) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g818 ( .A(n_503), .Y(n_818) );
INVx2_ASAP7_75t_L g1063 ( .A(n_503), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_503), .A2(n_815), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_504), .B(n_605), .Y(n_726) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_509), .Y(n_823) );
INVx1_ASAP7_75t_L g1056 ( .A(n_509), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1308 ( .A(n_509), .Y(n_1308) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g800 ( .A(n_511), .Y(n_800) );
INVx1_ASAP7_75t_L g824 ( .A(n_511), .Y(n_824) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_512), .Y(n_1059) );
INVx1_ASAP7_75t_L g1176 ( .A(n_512), .Y(n_1176) );
OAI31xp33_ASAP7_75t_L g789 ( .A1(n_513), .A2(n_790), .A3(n_792), .B(n_799), .Y(n_789) );
OAI31xp33_ASAP7_75t_L g1299 ( .A1(n_513), .A2(n_1300), .A3(n_1301), .B(n_1307), .Y(n_1299) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI31xp33_ASAP7_75t_L g809 ( .A1(n_514), .A2(n_810), .A3(n_819), .B(n_822), .Y(n_809) );
BUFx2_ASAP7_75t_SL g1065 ( .A(n_514), .Y(n_1065) );
INVx1_ASAP7_75t_L g1170 ( .A(n_514), .Y(n_1170) );
OAI31xp33_ASAP7_75t_L g1347 ( .A1(n_514), .A2(n_1348), .A3(n_1353), .B(n_1354), .Y(n_1347) );
BUFx2_ASAP7_75t_L g1394 ( .A(n_514), .Y(n_1394) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVxp67_ASAP7_75t_L g530 ( .A(n_516), .Y(n_530) );
INVx1_ASAP7_75t_L g536 ( .A(n_516), .Y(n_536) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_516), .B(n_726), .Y(n_1149) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
XOR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_650), .Y(n_518) );
INVx1_ASAP7_75t_L g648 ( .A(n_520), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .C(n_556), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_523), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_522), .A2(n_615), .B1(n_618), .B2(n_619), .Y(n_614) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx5_ASAP7_75t_L g947 ( .A(n_524), .Y(n_947) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
BUFx3_ASAP7_75t_L g631 ( .A(n_526), .Y(n_631) );
INVx8_ASAP7_75t_L g644 ( .A(n_526), .Y(n_644) );
BUFx3_ASAP7_75t_L g680 ( .A(n_526), .Y(n_680) );
AND2x4_ASAP7_75t_L g560 ( .A(n_528), .B(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B1(n_548), .B2(n_549), .Y(n_531) );
INVxp67_ASAP7_75t_L g1621 ( .A(n_533), .Y(n_1621) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_541), .Y(n_533) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND2x4_ASAP7_75t_L g553 ( .A(n_536), .B(n_554), .Y(n_553) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_537), .Y(n_699) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_L g554 ( .A(n_538), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g615 ( .A(n_538), .B(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_SL g620 ( .A(n_538), .B(n_584), .Y(n_620) );
AND2x4_ASAP7_75t_L g703 ( .A(n_538), .B(n_555), .Y(n_703) );
BUFx2_ASAP7_75t_L g928 ( .A(n_538), .Y(n_928) );
AND2x4_ASAP7_75t_L g1116 ( .A(n_538), .B(n_712), .Y(n_1116) );
INVx3_ASAP7_75t_L g589 ( .A(n_539), .Y(n_589) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_539), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_539), .B(n_605), .Y(n_720) );
OR2x6_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
INVx2_ASAP7_75t_SL g830 ( .A(n_542), .Y(n_830) );
OR2x2_ASAP7_75t_L g1165 ( .A(n_542), .B(n_544), .Y(n_1165) );
OAI22xp33_ASAP7_75t_L g1687 ( .A1(n_542), .A2(n_834), .B1(n_1673), .B2(n_1679), .Y(n_1687) );
OAI22xp33_ASAP7_75t_L g1691 ( .A1(n_542), .A2(n_754), .B1(n_1674), .B2(n_1680), .Y(n_1691) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
INVx3_ASAP7_75t_L g750 ( .A(n_543), .Y(n_750) );
INVxp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g573 ( .A(n_546), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g892 ( .A(n_546), .Y(n_892) );
INVx1_ASAP7_75t_L g1622 ( .A(n_549), .Y(n_1622) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g582 ( .A(n_555), .Y(n_582) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_555), .Y(n_609) );
INVx2_ASAP7_75t_L g931 ( .A(n_555), .Y(n_931) );
NOR3xp33_ASAP7_75t_SL g556 ( .A(n_557), .B(n_578), .C(n_623), .Y(n_556) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_559), .A2(n_565), .B1(n_635), .B2(n_915), .C(n_916), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_559), .A2(n_565), .B1(n_635), .B2(n_971), .C(n_972), .Y(n_970) );
AND2x4_ASAP7_75t_SL g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x4_ASAP7_75t_SL g565 ( .A(n_560), .B(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g635 ( .A(n_560), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_560), .B(n_562), .Y(n_1161) );
AND2x4_ASAP7_75t_L g1163 ( .A(n_560), .B(n_566), .Y(n_1163) );
NAND2x1_ASAP7_75t_L g1626 ( .A(n_560), .B(n_562), .Y(n_1626) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_561), .B(n_720), .Y(n_1145) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_575), .B2(n_576), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_571), .B(n_594), .Y(n_593) );
AOI222xp33_ASAP7_75t_L g888 ( .A1(n_572), .A2(n_576), .B1(n_889), .B2(n_890), .C1(n_893), .C2(n_894), .Y(n_888) );
AOI222xp33_ASAP7_75t_L g959 ( .A1(n_572), .A2(n_576), .B1(n_890), .B2(n_960), .C1(n_961), .C2(n_962), .Y(n_959) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_573), .B(n_1145), .Y(n_1144) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_574), .Y(n_1334) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_575), .A2(n_596), .B1(n_598), .B2(n_600), .C(n_601), .Y(n_595) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_577), .B(n_1149), .Y(n_1148) );
AOI31xp33_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_606), .A3(n_614), .B(n_621), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_587), .B(n_592), .Y(n_579) );
INVx2_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g929 ( .A1(n_583), .A2(n_911), .B1(n_916), .B2(n_930), .C(n_932), .Y(n_929) );
AOI221xp5_ASAP7_75t_L g984 ( .A1(n_583), .A2(n_930), .B1(n_958), .B2(n_972), .C(n_985), .Y(n_984) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x6_ASAP7_75t_L g727 ( .A(n_584), .B(n_605), .Y(n_727) );
BUFx3_ASAP7_75t_L g937 ( .A(n_584), .Y(n_937) );
BUFx3_ASAP7_75t_L g1119 ( .A(n_584), .Y(n_1119) );
INVx1_ASAP7_75t_L g1140 ( .A(n_584), .Y(n_1140) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx3_ASAP7_75t_L g716 ( .A(n_586), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_586), .A2(n_922), .B1(n_923), .B2(n_924), .C(n_925), .Y(n_921) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_586), .A2(n_861), .B1(n_922), .B2(n_981), .C(n_982), .Y(n_980) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx2_ASAP7_75t_SL g594 ( .A(n_589), .Y(n_594) );
INVx1_ASAP7_75t_L g612 ( .A(n_589), .Y(n_612) );
INVx2_ASAP7_75t_L g1124 ( .A(n_589), .Y(n_1124) );
BUFx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx3_ASAP7_75t_L g613 ( .A(n_591), .Y(n_613) );
INVx2_ASAP7_75t_L g617 ( .A(n_591), .Y(n_617) );
BUFx6f_ASAP7_75t_L g712 ( .A(n_591), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B(n_603), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g989 ( .A1(n_596), .A2(n_960), .B1(n_971), .B2(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1635 ( .A1(n_596), .A2(n_990), .B1(n_1627), .B2(n_1636), .Y(n_1635) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NOR2x1_ASAP7_75t_L g722 ( .A(n_599), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g933 ( .A1(n_604), .A2(n_711), .B(n_894), .C(n_934), .Y(n_933) );
A2O1A1Ixp33_ASAP7_75t_L g1632 ( .A1(n_604), .A2(n_979), .B(n_1633), .C(n_1634), .Y(n_1632) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g723 ( .A(n_605), .Y(n_723) );
INVx2_ASAP7_75t_L g700 ( .A(n_615), .Y(n_700) );
INVx3_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI211xp5_ASAP7_75t_SL g718 ( .A1(n_619), .A2(n_662), .B(n_719), .C(n_727), .Y(n_718) );
BUFx3_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g1132 ( .A(n_620), .Y(n_1132) );
BUFx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI211xp5_ASAP7_75t_SL g623 ( .A1(n_624), .A2(n_633), .B(n_634), .C(n_637), .Y(n_623) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI33xp33_ASAP7_75t_L g1003 ( .A1(n_633), .A2(n_694), .A3(n_1004), .B1(n_1010), .B2(n_1013), .B3(n_1020), .Y(n_1003) );
OAI33xp33_ASAP7_75t_L g1069 ( .A1(n_633), .A2(n_694), .A3(n_1070), .B1(n_1073), .B2(n_1076), .B3(n_1080), .Y(n_1069) );
OAI33xp33_ASAP7_75t_L g1210 ( .A1(n_633), .A2(n_694), .A3(n_1211), .B1(n_1215), .B2(n_1216), .B3(n_1219), .Y(n_1210) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_634), .Y(n_1167) );
INVx3_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g1649 ( .A1(n_635), .A2(n_647), .B1(n_1650), .B2(n_1654), .C(n_1660), .Y(n_1649) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .C(n_647), .Y(n_637) );
INVx1_ASAP7_75t_L g675 ( .A(n_639), .Y(n_675) );
BUFx12f_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx3_ASAP7_75t_L g900 ( .A(n_641), .Y(n_900) );
BUFx3_ASAP7_75t_L g904 ( .A(n_641), .Y(n_904) );
INVx5_ASAP7_75t_L g966 ( .A(n_641), .Y(n_966) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g891 ( .A(n_644), .Y(n_891) );
INVx8_ASAP7_75t_L g898 ( .A(n_644), .Y(n_898) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g681 ( .A(n_646), .Y(n_681) );
INVx1_ASAP7_75t_L g906 ( .A(n_646), .Y(n_906) );
INVx2_ASAP7_75t_L g694 ( .A(n_647), .Y(n_694) );
CKINVDCx5p33_ASAP7_75t_R g759 ( .A(n_647), .Y(n_759) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_672), .B(n_673), .C(n_695), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_654), .B(n_658), .C(n_666), .D(n_671), .Y(n_653) );
INVx2_ASAP7_75t_L g1237 ( .A(n_657), .Y(n_1237) );
AOI222xp33_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_662), .B2(n_663), .C1(n_664), .C2(n_665), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_660), .A2(n_663), .B1(n_785), .B2(n_786), .Y(n_784) );
BUFx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx3_ASAP7_75t_L g876 ( .A(n_661), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_663), .A2(n_816), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_663), .A2(n_876), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_663), .A2(n_876), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_663), .A2(n_876), .B1(n_1181), .B2(n_1188), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_664), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g693 ( .A(n_665), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_666) );
INVx2_ASAP7_75t_L g1049 ( .A(n_668), .Y(n_1049) );
INVx1_ASAP7_75t_L g879 ( .A(n_670), .Y(n_879) );
INVx2_ASAP7_75t_L g1097 ( .A(n_670), .Y(n_1097) );
OAI31xp33_ASAP7_75t_L g1089 ( .A1(n_672), .A2(n_1090), .A3(n_1096), .B(n_1098), .Y(n_1089) );
CKINVDCx14_ASAP7_75t_R g1191 ( .A(n_672), .Y(n_1191) );
OAI31xp33_ASAP7_75t_L g1309 ( .A1(n_672), .A2(n_1310), .A3(n_1311), .B(n_1316), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_682), .B1(n_684), .B2(n_694), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g1215 ( .A1(n_675), .A2(n_839), .B1(n_1202), .B2(n_1208), .Y(n_1215) );
BUFx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g691 ( .A(n_680), .Y(n_691) );
INVx2_ASAP7_75t_SL g1155 ( .A(n_680), .Y(n_1155) );
OAI33xp33_ASAP7_75t_L g740 ( .A1(n_682), .A2(n_741), .A3(n_748), .B1(n_755), .B2(n_759), .B3(n_760), .Y(n_740) );
OAI33xp33_ASAP7_75t_L g826 ( .A1(n_682), .A2(n_827), .A3(n_835), .B1(n_840), .B2(n_845), .B3(n_848), .Y(n_826) );
BUFx3_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI33xp33_ASAP7_75t_L g1686 ( .A1(n_683), .A2(n_1687), .A3(n_1688), .B1(n_1690), .B2(n_1691), .B3(n_1692), .Y(n_1686) );
OAI221xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_687), .B2(n_688), .C(n_689), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_685), .A2(n_1252), .B1(n_1262), .B2(n_1270), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_685), .A2(n_687), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
OAI22xp5_ASAP7_75t_L g1332 ( .A1(n_685), .A2(n_1333), .B1(n_1334), .B2(n_1335), .Y(n_1332) );
OAI22xp5_ASAP7_75t_L g1370 ( .A1(n_685), .A2(n_1270), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
OAI211xp5_ASAP7_75t_SL g713 ( .A1(n_686), .A2(n_706), .B(n_714), .C(n_717), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_687), .A2(n_1203), .B1(n_1209), .B2(n_1217), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g1271 ( .A1(n_687), .A2(n_1254), .B1(n_1263), .B2(n_1272), .Y(n_1271) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_687), .A2(n_1272), .B1(n_1374), .B2(n_1375), .Y(n_1373) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_718), .B(n_728), .Y(n_695) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1125 ( .A1(n_699), .A2(n_1126), .B1(n_1127), .B2(n_1128), .Y(n_1125) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_703), .Y(n_1128) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B(n_707), .C(n_710), .Y(n_704) );
INVx1_ASAP7_75t_L g1303 ( .A(n_706), .Y(n_1303) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_706), .A2(n_1253), .B1(n_1330), .B2(n_1333), .Y(n_1344) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_706), .A2(n_1253), .B1(n_1327), .B2(n_1338), .Y(n_1345) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g715 ( .A(n_709), .Y(n_715) );
INVx3_ASAP7_75t_L g920 ( .A(n_711), .Y(n_920) );
BUFx6f_ASAP7_75t_L g979 ( .A(n_711), .Y(n_979) );
A2O1A1Ixp33_ASAP7_75t_L g987 ( .A1(n_711), .A2(n_962), .B(n_988), .C(n_991), .Y(n_987) );
INVx1_ASAP7_75t_L g978 ( .A(n_712), .Y(n_978) );
INVx2_ASAP7_75t_L g1121 ( .A(n_715), .Y(n_1121) );
BUFx2_ASAP7_75t_L g1133 ( .A(n_721), .Y(n_1133) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g991 ( .A(n_723), .Y(n_991) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AOI21xp5_ASAP7_75t_SL g1117 ( .A1(n_727), .A2(n_1118), .B(n_1123), .Y(n_1117) );
INVx1_ASAP7_75t_L g1141 ( .A(n_728), .Y(n_1141) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
HB1xp67_ASAP7_75t_L g1648 ( .A(n_729), .Y(n_1648) );
BUFx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI31xp33_ASAP7_75t_L g917 ( .A1(n_730), .A2(n_918), .A3(n_926), .B(n_936), .Y(n_917) );
OAI31xp33_ASAP7_75t_L g975 ( .A1(n_730), .A2(n_976), .A3(n_983), .B(n_992), .Y(n_975) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND3xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_779), .C(n_789), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_765), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_L g837 ( .A(n_744), .Y(n_837) );
INVx8_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
BUFx3_ASAP7_75t_L g761 ( .A(n_745), .Y(n_761) );
INVx5_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g903 ( .A(n_746), .Y(n_903) );
INVx3_ASAP7_75t_L g1017 ( .A(n_746), .Y(n_1017) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_746), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_747), .A2(n_764), .B1(n_776), .B2(n_777), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_748) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_749), .A2(n_756), .B1(n_767), .B2(n_768), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g1266 ( .A1(n_750), .A2(n_1248), .B1(n_1256), .B2(n_1267), .Y(n_1266) );
OAI22xp33_ASAP7_75t_L g1273 ( .A1(n_750), .A2(n_754), .B1(n_1250), .B2(n_1258), .Y(n_1273) );
BUFx4f_ASAP7_75t_SL g1326 ( .A(n_750), .Y(n_1326) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_750), .A2(n_834), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_751), .A2(n_758), .B1(n_773), .B2(n_774), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g755 ( .A1(n_752), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_752), .A2(n_829), .B1(n_849), .B2(n_850), .Y(n_848) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_752), .A2(n_1006), .B1(n_1081), .B2(n_1082), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g1211 ( .A1(n_752), .A2(n_1196), .B1(n_1205), .B2(n_1212), .Y(n_1211) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g1399 ( .A(n_753), .Y(n_1399) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
BUFx6f_ASAP7_75t_L g1009 ( .A(n_754), .Y(n_1009) );
OAI22xp33_ASAP7_75t_L g1376 ( .A1(n_757), .A2(n_1377), .B1(n_1378), .B2(n_1379), .Y(n_1376) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_763), .A2(n_837), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_763), .A2(n_837), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
OAI33xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_769), .A3(n_770), .B1(n_772), .B2(n_775), .B3(n_778), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_767), .A2(n_1136), .B1(n_1331), .B2(n_1335), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g1384 ( .A1(n_767), .A2(n_1136), .B1(n_1372), .B2(n_1375), .Y(n_1384) );
OAI33xp33_ASAP7_75t_L g851 ( .A1(n_769), .A2(n_852), .A3(n_860), .B1(n_864), .B2(n_865), .B3(n_868), .Y(n_851) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_771), .A2(n_1256), .B1(n_1257), .B2(n_1258), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1385 ( .A1(n_771), .A2(n_1257), .B1(n_1368), .B2(n_1378), .Y(n_1385) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_777), .A2(n_1005), .B1(n_1021), .B2(n_1026), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_777), .A2(n_1026), .B1(n_1071), .B2(n_1081), .Y(n_1084) );
OAI33xp33_ASAP7_75t_L g1023 ( .A1(n_778), .A2(n_1024), .A3(n_1025), .B1(n_1028), .B2(n_1031), .B3(n_1033), .Y(n_1023) );
OAI33xp33_ASAP7_75t_L g1083 ( .A1(n_778), .A2(n_1024), .A3(n_1084), .B1(n_1085), .B2(n_1086), .B3(n_1088), .Y(n_1083) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g812 ( .A(n_796), .Y(n_812) );
INVx3_ASAP7_75t_L g1183 ( .A(n_796), .Y(n_1183) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
XNOR2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_998), .Y(n_802) );
XNOR2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_883), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_825), .C(n_869), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g1085 ( .A1(n_811), .A2(n_940), .B1(n_1074), .B2(n_1077), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_814), .A2(n_1046), .B1(n_1062), .B2(n_1064), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_814), .A2(n_1062), .B1(n_1094), .B2(n_1106), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_814), .A2(n_818), .B1(n_1181), .B2(n_1182), .Y(n_1180) );
BUFx3_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_818), .A2(n_1696), .B1(n_1697), .B2(n_1698), .Y(n_1695) );
NOR2xp33_ASAP7_75t_SL g825 ( .A(n_826), .B(n_851), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_829), .B1(n_831), .B2(n_832), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_828), .A2(n_849), .B1(n_853), .B2(n_857), .Y(n_852) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g1220 ( .A(n_830), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_831), .A2(n_850), .B1(n_861), .B2(n_863), .Y(n_864) );
INVx2_ASAP7_75t_SL g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B1(n_838), .B2(n_839), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_836), .A2(n_843), .B1(n_861), .B2(n_863), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_838), .A2(n_844), .B1(n_853), .B2(n_857), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_839), .A2(n_841), .B1(n_843), .B2(n_844), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g1690 ( .A1(n_839), .A2(n_903), .B1(n_1677), .B2(n_1685), .Y(n_1690) );
INVx3_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
AND2x4_ASAP7_75t_L g912 ( .A(n_842), .B(n_892), .Y(n_912) );
INVx3_ASAP7_75t_L g1078 ( .A(n_842), .Y(n_1078) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_842), .Y(n_1272) );
INVx2_ASAP7_75t_SL g1656 ( .A(n_842), .Y(n_1656) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_SL g854 ( .A(n_855), .Y(n_854) );
INVx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx4_ASAP7_75t_L g943 ( .A(n_856), .Y(n_943) );
BUFx6f_ASAP7_75t_L g1027 ( .A(n_856), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_857), .A2(n_1196), .B1(n_1197), .B2(n_1200), .Y(n_1195) );
OAI22xp5_ASAP7_75t_L g1207 ( .A1(n_857), .A2(n_1197), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_859), .A2(n_942), .B1(n_943), .B2(n_944), .Y(n_941) );
OAI22xp33_ASAP7_75t_L g1247 ( .A1(n_859), .A2(n_1248), .B1(n_1249), .B2(n_1250), .Y(n_1247) );
OAI22xp33_ASAP7_75t_L g1383 ( .A1(n_859), .A2(n_1249), .B1(n_1367), .B2(n_1377), .Y(n_1383) );
INVx1_ASAP7_75t_L g1030 ( .A(n_861), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1201 ( .A1(n_861), .A2(n_863), .B1(n_1202), .B2(n_1203), .Y(n_1201) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
INVx2_ASAP7_75t_L g925 ( .A(n_862), .Y(n_925) );
BUFx2_ASAP7_75t_L g1296 ( .A(n_862), .Y(n_1296) );
OAI33xp33_ASAP7_75t_L g1193 ( .A1(n_865), .A2(n_1194), .A3(n_1195), .B1(n_1201), .B2(n_1204), .B3(n_1207), .Y(n_1193) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OAI31xp33_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_874), .A3(n_878), .B(n_881), .Y(n_869) );
INVx2_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_949), .B1(n_950), .B2(n_997), .Y(n_883) );
INVx1_ASAP7_75t_L g997 ( .A(n_884), .Y(n_997) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
XNOR2x1_ASAP7_75t_L g885 ( .A(n_886), .B(n_948), .Y(n_885) );
OR2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_913), .Y(n_886) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_895), .C(n_910), .Y(n_887) );
AND2x4_ASAP7_75t_L g890 ( .A(n_891), .B(n_892), .Y(n_890) );
AOI33xp33_ASAP7_75t_L g895 ( .A1(n_896), .A2(n_897), .A3(n_899), .B1(n_901), .B2(n_905), .B3(n_907), .Y(n_895) );
NAND3xp33_ASAP7_75t_L g954 ( .A(n_896), .B(n_955), .C(n_956), .Y(n_954) );
AOI33xp33_ASAP7_75t_L g1152 ( .A1(n_896), .A2(n_907), .A3(n_1153), .B1(n_1156), .B2(n_1157), .B3(n_1158), .Y(n_1152) );
BUFx3_ASAP7_75t_L g1660 ( .A(n_896), .Y(n_1660) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
NAND3xp33_ASAP7_75t_L g963 ( .A(n_907), .B(n_964), .C(n_967), .Y(n_963) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI33xp33_ASAP7_75t_L g1264 ( .A1(n_908), .A2(n_1265), .A3(n_1266), .B1(n_1269), .B2(n_1271), .B3(n_1273), .Y(n_1264) );
OAI33xp33_ASAP7_75t_L g1323 ( .A1(n_908), .A2(n_1265), .A3(n_1324), .B1(n_1329), .B2(n_1332), .B3(n_1336), .Y(n_1323) );
OAI33xp33_ASAP7_75t_L g1365 ( .A1(n_908), .A2(n_1265), .A3(n_1366), .B1(n_1370), .B2(n_1373), .B3(n_1376), .Y(n_1365) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_912), .B(n_958), .Y(n_957) );
INVx2_ASAP7_75t_L g1166 ( .A(n_912), .Y(n_1166) );
NAND3xp33_ASAP7_75t_SL g913 ( .A(n_914), .B(n_917), .C(n_945), .Y(n_913) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_922), .A2(n_1280), .B1(n_1290), .B2(n_1295), .Y(n_1294) );
OAI211xp5_ASAP7_75t_L g1642 ( .A1(n_922), .A2(n_1643), .B(n_1644), .C(n_1645), .Y(n_1642) );
OAI22xp5_ASAP7_75t_L g1678 ( .A1(n_925), .A2(n_1228), .B1(n_1679), .B2(n_1680), .Y(n_1678) );
OAI21xp33_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_929), .B(n_933), .Y(n_926) );
OAI21xp5_ASAP7_75t_SL g983 ( .A1(n_927), .A2(n_984), .B(n_987), .Y(n_983) );
INVxp67_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
HB1xp67_ASAP7_75t_L g1032 ( .A(n_940), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g1681 ( .A1(n_943), .A2(n_1682), .B1(n_1683), .B2(n_1685), .Y(n_1681) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_946), .B(n_947), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_947), .B(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
XNOR2x1_ASAP7_75t_L g951 ( .A(n_952), .B(n_996), .Y(n_951) );
OR2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_969), .Y(n_952) );
NAND4xp25_ASAP7_75t_SL g953 ( .A(n_954), .B(n_957), .C(n_959), .D(n_963), .Y(n_953) );
INVx2_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
NAND3xp33_ASAP7_75t_SL g969 ( .A(n_970), .B(n_973), .C(n_975), .Y(n_969) );
INVx1_ASAP7_75t_L g977 ( .A(n_978), .Y(n_977) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
XOR2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1066), .Y(n_999) );
AND3x1_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1040), .C(n_1051), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1023), .Y(n_1002) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1006), .B1(n_1008), .B2(n_1009), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1020 ( .A1(n_1006), .A2(n_1009), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
OAI22xp33_ASAP7_75t_L g1070 ( .A1(n_1006), .A2(n_1009), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
OAI22xp33_ASAP7_75t_L g1288 ( .A1(n_1006), .A2(n_1092), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OAI22xp33_ASAP7_75t_L g1219 ( .A1(n_1009), .A2(n_1200), .B1(n_1206), .B2(n_1220), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1033 ( .A1(n_1012), .A2(n_1018), .B1(n_1034), .B2(n_1038), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1018), .B2(n_1019), .Y(n_1013) );
INVx2_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx2_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_1019), .A2(n_1077), .B1(n_1078), .B2(n_1079), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1688 ( .A1(n_1019), .A2(n_1676), .B1(n_1682), .B2(n_1689), .Y(n_1688) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVxp67_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1044), .Y(n_1328) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1044), .Y(n_1369) );
OAI31xp33_ASAP7_75t_SL g1051 ( .A1(n_1052), .A2(n_1054), .A3(n_1060), .B(n_1065), .Y(n_1051) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_1059), .Y(n_1058) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1063), .Y(n_1351) );
OAI31xp33_ASAP7_75t_L g1101 ( .A1(n_1065), .A2(n_1102), .A3(n_1103), .B(n_1104), .Y(n_1101) );
OAI31xp33_ASAP7_75t_L g1226 ( .A1(n_1065), .A2(n_1227), .A3(n_1232), .B(n_1233), .Y(n_1226) );
AND3x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1089), .C(n_1101), .Y(n_1067) );
NOR2xp33_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1083), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
OA22x2_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1221), .B1(n_1222), .B2(n_1404), .Y(n_1107) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1108), .Y(n_1404) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_1110), .Y(n_1109) );
XNOR2xp5_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1168), .Y(n_1110) );
NAND3xp33_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1142), .C(n_1150), .Y(n_1112) );
OAI21xp33_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1129), .B(n_1141), .Y(n_1113) );
INVx2_ASAP7_75t_SL g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1131), .Y(n_1647) );
INVx4_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AOI21xp33_ASAP7_75t_SL g1142 ( .A1(n_1143), .A2(n_1146), .B(n_1147), .Y(n_1142) );
INVx8_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
NOR3xp33_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1164), .C(n_1167), .Y(n_1150) );
NAND2xp5_ASAP7_75t_SL g1151 ( .A(n_1152), .B(n_1159), .Y(n_1151) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1160), .A2(n_1161), .B1(n_1162), .B2(n_1163), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1624 ( .A1(n_1163), .A2(n_1625), .B1(n_1627), .B2(n_1628), .C(n_1629), .Y(n_1624) );
OAI221xp5_ASAP7_75t_L g1169 ( .A1(n_1170), .A2(n_1171), .B1(n_1184), .B2(n_1191), .C(n_1192), .Y(n_1169) );
NOR3xp33_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1177), .C(n_1178), .Y(n_1171) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
OAI211xp5_ASAP7_75t_L g1637 ( .A1(n_1179), .A2(n_1638), .B(n_1639), .C(n_1641), .Y(n_1637) );
NOR3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .C(n_1189), .Y(n_1184) );
NOR2xp33_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1210), .Y(n_1192) );
OAI33xp33_ASAP7_75t_L g1246 ( .A1(n_1194), .A2(n_1247), .A3(n_1251), .B1(n_1255), .B2(n_1259), .B3(n_1261), .Y(n_1246) );
INVx2_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
OAI22xp5_ASAP7_75t_L g1657 ( .A1(n_1214), .A2(n_1267), .B1(n_1658), .B2(n_1659), .Y(n_1657) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
AOI22xp5_ASAP7_75t_L g1222 ( .A1(n_1223), .A2(n_1319), .B1(n_1402), .B2(n_1403), .Y(n_1222) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1223), .Y(n_1402) );
XNOR2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1274), .Y(n_1223) );
NAND3xp33_ASAP7_75t_L g1225 ( .A(n_1226), .B(n_1235), .C(n_1245), .Y(n_1225) );
OAI31xp33_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1238), .A3(n_1243), .B(n_1244), .Y(n_1235) );
HB1xp67_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
OAI31xp33_ASAP7_75t_L g1355 ( .A1(n_1244), .A2(n_1356), .A3(n_1357), .B(n_1360), .Y(n_1355) );
OAI31xp33_ASAP7_75t_SL g1395 ( .A1(n_1244), .A2(n_1396), .A3(n_1397), .B(n_1398), .Y(n_1395) );
NOR2xp33_ASAP7_75t_SL g1245 ( .A(n_1246), .B(n_1264), .Y(n_1245) );
OAI33xp33_ASAP7_75t_L g1339 ( .A1(n_1259), .A2(n_1340), .A3(n_1343), .B1(n_1344), .B2(n_1345), .B3(n_1346), .Y(n_1339) );
OAI33xp33_ASAP7_75t_L g1380 ( .A1(n_1259), .A2(n_1381), .A3(n_1382), .B1(n_1383), .B2(n_1384), .B3(n_1385), .Y(n_1380) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
NAND3xp33_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1299), .C(n_1309), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1291), .Y(n_1276) );
INVx4_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1403 ( .A(n_1319), .Y(n_1403) );
XOR2xp5_ASAP7_75t_L g1319 ( .A(n_1320), .B(n_1361), .Y(n_1319) );
NAND3xp33_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1347), .C(n_1355), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1339), .Y(n_1322) );
OAI22xp33_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1326), .B1(n_1327), .B2(n_1328), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1366 ( .A1(n_1326), .A2(n_1367), .B1(n_1368), .B2(n_1369), .Y(n_1366) );
OAI22xp5_ASAP7_75t_L g1651 ( .A1(n_1326), .A2(n_1643), .B1(n_1652), .B2(n_1653), .Y(n_1651) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx2_ASAP7_75t_SL g1341 ( .A(n_1342), .Y(n_1341) );
XNOR2xp5_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1363), .Y(n_1361) );
AND3x1_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1386), .C(n_1395), .Y(n_1363) );
NOR2xp33_ASAP7_75t_SL g1364 ( .A(n_1365), .B(n_1380), .Y(n_1364) );
OAI31xp33_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1388), .A3(n_1393), .B(n_1394), .Y(n_1386) );
OAI31xp33_ASAP7_75t_L g1693 ( .A1(n_1394), .A2(n_1694), .A3(n_1699), .B(n_1700), .Y(n_1693) );
OAI221xp5_ASAP7_75t_SL g1405 ( .A1(n_1406), .A2(n_1616), .B1(n_1617), .B2(n_1661), .C(n_1665), .Y(n_1405) );
AND5x1_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1572), .C(n_1589), .D(n_1598), .E(n_1609), .Y(n_1406) );
OAI33xp33_ASAP7_75t_L g1407 ( .A1(n_1408), .A2(n_1500), .A3(n_1517), .B1(n_1526), .B2(n_1553), .B3(n_1567), .Y(n_1407) );
OAI211xp5_ASAP7_75t_SL g1408 ( .A1(n_1409), .A2(n_1430), .B(n_1447), .C(n_1490), .Y(n_1408) );
CKINVDCx5p33_ASAP7_75t_R g1507 ( .A(n_1409), .Y(n_1507) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1425), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_1410), .A2(n_1457), .B1(n_1460), .B2(n_1463), .Y(n_1456) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1410), .B(n_1464), .Y(n_1463) );
OR2x2_ASAP7_75t_L g1499 ( .A(n_1410), .B(n_1426), .Y(n_1499) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1410), .Y(n_1510) );
INVx2_ASAP7_75t_L g1528 ( .A(n_1410), .Y(n_1528) );
OR2x2_ASAP7_75t_L g1542 ( .A(n_1410), .B(n_1466), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1410), .B(n_1465), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1597 ( .A(n_1410), .B(n_1466), .Y(n_1597) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
OR2x2_ASAP7_75t_L g1449 ( .A(n_1411), .B(n_1425), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_1412), .B(n_1419), .Y(n_1411) );
AND2x6_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1415), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1414), .B(n_1418), .Y(n_1417) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_1414), .B(n_1421), .Y(n_1420) );
AND2x6_ASAP7_75t_L g1423 ( .A(n_1414), .B(n_1424), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1414), .B(n_1418), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1414), .B(n_1418), .Y(n_1469) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1414), .B(n_1421), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1416), .B(n_1422), .Y(n_1421) );
HB1xp67_ASAP7_75t_L g1721 ( .A(n_1421), .Y(n_1721) );
INVx2_ASAP7_75t_L g1480 ( .A(n_1423), .Y(n_1480) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1425), .Y(n_1471) );
NOR2xp33_ASAP7_75t_L g1585 ( .A(n_1425), .B(n_1512), .Y(n_1585) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1464 ( .A(n_1426), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1429), .Y(n_1426) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1431), .B(n_1435), .Y(n_1430) );
NOR2xp33_ASAP7_75t_L g1457 ( .A(n_1431), .B(n_1458), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1431), .B(n_1493), .Y(n_1492) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1431), .B(n_1507), .Y(n_1525) );
CKINVDCx5p33_ASAP7_75t_R g1552 ( .A(n_1431), .Y(n_1552) );
AND2x2_ASAP7_75t_L g1559 ( .A(n_1431), .B(n_1461), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1568 ( .A(n_1431), .B(n_1474), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1431), .B(n_1471), .Y(n_1601) );
INVx4_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
O2A1O1Ixp33_ASAP7_75t_L g1483 ( .A1(n_1432), .A2(n_1484), .B(n_1486), .C(n_1489), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1432), .B(n_1488), .Y(n_1487) );
INVx4_ASAP7_75t_L g1503 ( .A(n_1432), .Y(n_1503) );
NOR2xp33_ASAP7_75t_L g1505 ( .A(n_1432), .B(n_1506), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1509 ( .A(n_1432), .B(n_1453), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1511 ( .A(n_1432), .B(n_1501), .Y(n_1511) );
NAND2xp5_ASAP7_75t_SL g1516 ( .A(n_1432), .B(n_1453), .Y(n_1516) );
NOR2xp33_ASAP7_75t_L g1523 ( .A(n_1432), .B(n_1454), .Y(n_1523) );
NOR3xp33_ASAP7_75t_L g1545 ( .A(n_1432), .B(n_1542), .C(n_1546), .Y(n_1545) );
AND2x2_ASAP7_75t_L g1596 ( .A(n_1432), .B(n_1495), .Y(n_1596) );
AND2x4_ASAP7_75t_SL g1432 ( .A(n_1433), .B(n_1434), .Y(n_1432) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1435), .B(n_1534), .Y(n_1571) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1439), .Y(n_1435) );
OR2x2_ASAP7_75t_L g1494 ( .A(n_1436), .B(n_1441), .Y(n_1494) );
OR2x2_ASAP7_75t_L g1539 ( .A(n_1436), .B(n_1540), .Y(n_1539) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1436), .B(n_1488), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1613 ( .A(n_1436), .B(n_1523), .Y(n_1613) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1438), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1437), .B(n_1438), .Y(n_1453) );
OR2x2_ASAP7_75t_L g1563 ( .A(n_1439), .B(n_1452), .Y(n_1563) );
NAND2xp5_ASAP7_75t_L g1610 ( .A(n_1439), .B(n_1611), .Y(n_1610) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1444), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1441), .B(n_1444), .Y(n_1454) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1441), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1474 ( .A(n_1441), .B(n_1444), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1441), .B(n_1462), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1441), .B(n_1453), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1443), .Y(n_1441) );
INVx2_ASAP7_75t_L g1462 ( .A(n_1444), .Y(n_1462) );
NAND2x1p5_ASAP7_75t_L g1444 ( .A(n_1445), .B(n_1446), .Y(n_1444) );
AOI211xp5_ASAP7_75t_L g1447 ( .A1(n_1448), .A2(n_1450), .B(n_1455), .C(n_1483), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1551 ( .A(n_1448), .B(n_1552), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g1448 ( .A(n_1449), .Y(n_1448) );
OR2x2_ASAP7_75t_L g1615 ( .A(n_1449), .B(n_1465), .Y(n_1615) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
NOR2xp33_ASAP7_75t_L g1543 ( .A(n_1451), .B(n_1497), .Y(n_1543) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1452), .B(n_1454), .Y(n_1451) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_1452), .B(n_1462), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1452), .B(n_1488), .Y(n_1495) );
AND2x2_ASAP7_75t_L g1549 ( .A(n_1452), .B(n_1514), .Y(n_1549) );
A2O1A1Ixp33_ASAP7_75t_L g1609 ( .A1(n_1452), .A2(n_1610), .B(n_1612), .C(n_1614), .Y(n_1609) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1458 ( .A(n_1453), .B(n_1459), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1453), .B(n_1474), .Y(n_1473) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1453), .B(n_1459), .Y(n_1485) );
OR2x2_ASAP7_75t_L g1506 ( .A(n_1453), .B(n_1462), .Y(n_1506) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1453), .B(n_1462), .Y(n_1582) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1454), .Y(n_1514) );
OR2x2_ASAP7_75t_L g1575 ( .A(n_1454), .B(n_1509), .Y(n_1575) );
OAI221xp5_ASAP7_75t_SL g1455 ( .A1(n_1456), .A2(n_1465), .B1(n_1470), .B2(n_1472), .C(n_1475), .Y(n_1455) );
HB1xp67_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1463), .Y(n_1556) );
OR2x2_ASAP7_75t_L g1489 ( .A(n_1464), .B(n_1465), .Y(n_1489) );
INVx2_ASAP7_75t_L g1501 ( .A(n_1464), .Y(n_1501) );
OAI221xp5_ASAP7_75t_L g1517 ( .A1(n_1464), .A2(n_1510), .B1(n_1518), .B2(n_1522), .C(n_1524), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1533 ( .A(n_1464), .B(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1464), .B(n_1503), .Y(n_1561) );
A2O1A1Ixp33_ASAP7_75t_L g1589 ( .A1(n_1464), .A2(n_1590), .B(n_1596), .C(n_1597), .Y(n_1589) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_1465), .B(n_1471), .Y(n_1470) );
A2O1A1Ixp33_ASAP7_75t_L g1504 ( .A1(n_1465), .A2(n_1505), .B(n_1507), .C(n_1508), .Y(n_1504) );
CKINVDCx14_ASAP7_75t_R g1566 ( .A(n_1465), .Y(n_1566) );
INVx3_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1466), .Y(n_1498) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_1466), .A2(n_1501), .B1(n_1573), .B2(n_1576), .C(n_1583), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1578 ( .A(n_1466), .B(n_1510), .Y(n_1578) );
OAI21xp33_ASAP7_75t_L g1583 ( .A1(n_1466), .A2(n_1584), .B(n_1586), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1468), .Y(n_1466) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1471), .Y(n_1520) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1473), .Y(n_1472) );
NAND2x1_ASAP7_75t_L g1502 ( .A(n_1473), .B(n_1503), .Y(n_1502) );
OAI21xp33_ASAP7_75t_L g1586 ( .A1(n_1473), .A2(n_1587), .B(n_1588), .Y(n_1586) );
OAI321xp33_ASAP7_75t_L g1508 ( .A1(n_1474), .A2(n_1484), .A3(n_1509), .B1(n_1510), .B2(n_1511), .C(n_1512), .Y(n_1508) );
INVx1_ASAP7_75t_L g1540 ( .A(n_1474), .Y(n_1540) );
OAI21xp5_ASAP7_75t_L g1548 ( .A1(n_1474), .A2(n_1549), .B(n_1550), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1474), .B(n_1515), .Y(n_1580) );
AOI211xp5_ASAP7_75t_L g1557 ( .A1(n_1475), .A2(n_1558), .B(n_1559), .C(n_1560), .Y(n_1557) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1476), .B(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1477), .Y(n_1476) );
OAI221xp5_ASAP7_75t_L g1477 ( .A1(n_1478), .A2(n_1479), .B1(n_1480), .B2(n_1481), .C(n_1482), .Y(n_1477) );
BUFx2_ASAP7_75t_L g1616 ( .A(n_1478), .Y(n_1616) );
NAND2xp5_ASAP7_75t_SL g1538 ( .A(n_1484), .B(n_1539), .Y(n_1538) );
O2A1O1Ixp33_ASAP7_75t_L g1553 ( .A1(n_1484), .A2(n_1554), .B(n_1557), .C(n_1564), .Y(n_1553) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1524 ( .A(n_1485), .B(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1488), .Y(n_1611) );
OAI322xp33_ASAP7_75t_L g1567 ( .A1(n_1489), .A2(n_1494), .A3(n_1498), .B1(n_1507), .B2(n_1568), .C1(n_1569), .C2(n_1570), .Y(n_1567) );
OAI21xp33_ASAP7_75t_L g1490 ( .A1(n_1491), .A2(n_1495), .B(n_1496), .Y(n_1490) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
INVxp67_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1521 ( .A(n_1494), .B(n_1503), .Y(n_1521) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_1495), .B(n_1507), .Y(n_1536) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1495), .Y(n_1606) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1498), .B(n_1499), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1600 ( .A(n_1498), .B(n_1601), .Y(n_1600) );
OAI21xp33_ASAP7_75t_L g1500 ( .A1(n_1501), .A2(n_1502), .B(n_1504), .Y(n_1500) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1501), .B(n_1542), .Y(n_1569) );
CKINVDCx5p33_ASAP7_75t_R g1534 ( .A(n_1503), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1608 ( .A(n_1507), .B(n_1552), .Y(n_1608) );
NOR2xp33_ASAP7_75t_L g1529 ( .A(n_1510), .B(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1558 ( .A(n_1510), .Y(n_1558) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
AOI211xp5_ASAP7_75t_L g1527 ( .A1(n_1513), .A2(n_1528), .B(n_1529), .C(n_1535), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g1605 ( .A(n_1513), .B(n_1520), .Y(n_1605) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1515), .Y(n_1513) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVxp67_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1519 ( .A(n_1520), .B(n_1521), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1520), .B(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
O2A1O1Ixp33_ASAP7_75t_L g1598 ( .A1(n_1525), .A2(n_1599), .B(n_1602), .C(n_1604), .Y(n_1598) );
NAND4xp25_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1537), .C(n_1544), .D(n_1548), .Y(n_1526) );
INVxp33_ASAP7_75t_L g1587 ( .A(n_1530), .Y(n_1587) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1533), .Y(n_1530) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1532), .Y(n_1531) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1532), .B(n_1552), .Y(n_1593) );
AOI31xp33_ASAP7_75t_L g1537 ( .A1(n_1534), .A2(n_1538), .A3(n_1541), .B(n_1543), .Y(n_1537) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_1534), .B(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
CKINVDCx14_ASAP7_75t_R g1541 ( .A(n_1542), .Y(n_1541) );
OAI22xp5_ASAP7_75t_L g1576 ( .A1(n_1542), .A2(n_1577), .B1(n_1579), .B2(n_1581), .Y(n_1576) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1546), .B(n_1595), .Y(n_1603) );
INVx1_ASAP7_75t_L g1546 ( .A(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1549), .Y(n_1595) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVxp67_ASAP7_75t_SL g1554 ( .A(n_1555), .Y(n_1554) );
OAI22xp5_ASAP7_75t_L g1604 ( .A1(n_1558), .A2(n_1605), .B1(n_1606), .B2(n_1607), .Y(n_1604) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1559), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1562), .Y(n_1560) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
CKINVDCx14_ASAP7_75t_R g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1584 ( .A(n_1585), .Y(n_1584) );
NAND2xp5_ASAP7_75t_L g1590 ( .A(n_1591), .B(n_1595), .Y(n_1590) );
INVxp67_ASAP7_75t_SL g1591 ( .A(n_1592), .Y(n_1591) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1593), .B(n_1594), .Y(n_1592) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVxp67_ASAP7_75t_L g1602 ( .A(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
HB1xp67_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
NOR2x1_ASAP7_75t_L g1619 ( .A(n_1620), .B(n_1623), .Y(n_1619) );
NAND3xp33_ASAP7_75t_SL g1623 ( .A(n_1624), .B(n_1630), .C(n_1649), .Y(n_1623) );
INVx2_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
OAI21xp5_ASAP7_75t_L g1630 ( .A1(n_1631), .A2(n_1646), .B(n_1648), .Y(n_1630) );
NAND3xp33_ASAP7_75t_L g1631 ( .A(n_1632), .B(n_1637), .C(n_1642), .Y(n_1631) );
INVx1_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
CKINVDCx5p33_ASAP7_75t_R g1661 ( .A(n_1662), .Y(n_1661) );
BUFx2_ASAP7_75t_SL g1662 ( .A(n_1663), .Y(n_1662) );
BUFx3_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVxp67_ASAP7_75t_SL g1666 ( .A(n_1667), .Y(n_1666) );
HB1xp67_ASAP7_75t_SL g1667 ( .A(n_1668), .Y(n_1667) );
AND3x1_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1693), .C(n_1702), .Y(n_1669) );
NOR2xp33_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1686), .Y(n_1670) );
BUFx6f_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
AOI22xp33_ASAP7_75t_SL g1709 ( .A1(n_1697), .A2(n_1710), .B1(n_1711), .B2(n_1712), .Y(n_1709) );
OAI31xp33_ASAP7_75t_SL g1702 ( .A1(n_1703), .A2(n_1706), .A3(n_1713), .B(n_1714), .Y(n_1702) );
INVx2_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
BUFx4f_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
HB1xp67_ASAP7_75t_L g1718 ( .A(n_1719), .Y(n_1718) );
OAI21xp5_ASAP7_75t_L g1719 ( .A1(n_1720), .A2(n_1721), .B(n_1722), .Y(n_1719) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
endmodule