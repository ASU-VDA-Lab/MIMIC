module fake_jpeg_4228_n_264 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_82;
wire n_258;
wire n_96;

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_2),
.B(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_42),
.B(n_48),
.Y(n_96)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_23),
.B(n_29),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_53),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_47),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_28),
.B(n_0),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_1),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_74),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_37),
.B1(n_20),
.B2(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_75),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_37),
.B1(n_25),
.B2(n_36),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_31),
.B1(n_36),
.B2(n_23),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_34),
.B1(n_33),
.B2(n_35),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_77),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_90),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_61),
.A2(n_34),
.B1(n_35),
.B2(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_100),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_42),
.A2(n_38),
.B1(n_35),
.B2(n_30),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_21),
.B1(n_30),
.B2(n_3),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_15),
.B1(n_11),
.B2(n_12),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_97),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_103),
.Y(n_133)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_118),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_47),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_45),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_113),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

NAND3xp33_ASAP7_75t_SL g116 ( 
.A(n_65),
.B(n_49),
.C(n_48),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_98),
.B(n_4),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_5),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_68),
.B(n_45),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_124),
.B(n_129),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_73),
.A2(n_45),
.B(n_39),
.C(n_10),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_125),
.A2(n_129),
.B(n_130),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_14),
.C(n_15),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_130),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_5),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_8),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_100),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_62),
.B1(n_64),
.B2(n_72),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_145),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_102),
.B(n_114),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_76),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_158),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_111),
.A2(n_84),
.B1(n_95),
.B2(n_82),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_69),
.B1(n_86),
.B2(n_89),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_143),
.A2(n_144),
.B1(n_151),
.B2(n_155),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_122),
.A2(n_82),
.B1(n_84),
.B2(n_64),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_109),
.B(n_63),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_147),
.Y(n_167)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_104),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_80),
.B(n_81),
.C(n_87),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_106),
.A2(n_80),
.B1(n_97),
.B2(n_92),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_154),
.A2(n_140),
.B1(n_158),
.B2(n_160),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_10),
.B1(n_11),
.B2(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_157),
.B(n_134),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_125),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_128),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_103),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_124),
.C(n_127),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_176),
.C(n_170),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_163),
.B(n_179),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_145),
.B1(n_159),
.B2(n_171),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_147),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_114),
.B1(n_107),
.B2(n_120),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_134),
.B(n_156),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_180),
.B(n_170),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_135),
.A2(n_107),
.B1(n_128),
.B2(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g180 ( 
.A1(n_151),
.A2(n_144),
.B(n_141),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_183),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_167),
.B(n_135),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_187),
.B(n_191),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_190),
.B(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_197),
.C(n_162),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_182),
.B(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_194),
.B(n_196),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_205),
.Y(n_207)
);

OAI211xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_174),
.B(n_186),
.C(n_184),
.Y(n_198)
);

NOR3xp33_ASAP7_75t_L g221 ( 
.A(n_198),
.B(n_166),
.C(n_169),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_167),
.B(n_181),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_188),
.B(n_202),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_166),
.Y(n_205)
);

XOR2x2_ASAP7_75t_SL g206 ( 
.A(n_163),
.B(n_180),
.Y(n_206)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_206),
.A2(n_177),
.B(n_175),
.C(n_178),
.D(n_185),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_203),
.B1(n_171),
.B2(n_205),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_212),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_213),
.C(n_214),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_192),
.B(n_168),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_165),
.C(n_172),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_215),
.Y(n_232)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_180),
.Y(n_216)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_216),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_202),
.B(n_199),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_221),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_200),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_197),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_229),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_211),
.C(n_213),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_189),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_241),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g239 ( 
.A(n_228),
.Y(n_239)
);

BUFx24_ASAP7_75t_SL g243 ( 
.A(n_239),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_206),
.C(n_212),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_203),
.B1(n_220),
.B2(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_232),
.Y(n_247)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_244),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_248),
.B(n_249),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_223),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_225),
.B1(n_201),
.B2(n_224),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_253),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_209),
.A3(n_225),
.B1(n_207),
.B2(n_241),
.C1(n_226),
.C2(n_227),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_235),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_210),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_222),
.B(n_217),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_255),
.A2(n_256),
.B(n_258),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_229),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_251),
.B(n_201),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_190),
.B1(n_195),
.B2(n_243),
.Y(n_262)
);

OA21x2_ASAP7_75t_SL g263 ( 
.A1(n_262),
.A2(n_173),
.B(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_173),
.Y(n_264)
);


endmodule