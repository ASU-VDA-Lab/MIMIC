module fake_jpeg_1542_n_79 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_1),
.B(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_35),
.Y(n_39)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_3),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_51),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_28),
.B1(n_26),
.B2(n_33),
.Y(n_48)
);

NAND2x1_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_33),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_43),
.B1(n_28),
.B2(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_1),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_SL g54 ( 
.A(n_49),
.B(n_39),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_54),
.A2(n_5),
.B(n_6),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_4),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_47),
.B1(n_6),
.B2(n_7),
.Y(n_62)
);

AND2x4_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_68),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_56),
.B1(n_54),
.B2(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_64),
.B1(n_63),
.B2(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_71),
.C(n_65),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_74),
.A2(n_66),
.B(n_70),
.C(n_12),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_18),
.A3(n_9),
.B1(n_13),
.B2(n_14),
.C1(n_17),
.C2(n_23),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_19),
.C(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_22),
.B1(n_8),
.B2(n_70),
.Y(n_79)
);


endmodule