module fake_aes_125_n_8 (n_3, n_1, n_2, n_0, n_8);
input n_3;
input n_1;
input n_2;
input n_0;
output n_8;
wire n_6;
wire n_4;
wire n_5;
wire n_7;
NAND2xp5_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_3), .B(n_1), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_4), .B(n_0), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
OAI21x1_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_5), .B(n_2), .Y(n_8) );
endmodule