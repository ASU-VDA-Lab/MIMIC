module real_jpeg_26865_n_16 (n_333, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_333;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_0),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_0),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_0),
.A2(n_35),
.B1(n_63),
.B2(n_66),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_31),
.B1(n_33),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_1),
.A2(n_51),
.B1(n_63),
.B2(n_66),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_124)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_2),
.Y(n_107)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_3),
.A2(n_54),
.B1(n_63),
.B2(n_66),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_54),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_5),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_37),
.B1(n_63),
.B2(n_66),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_8),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_149),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_149),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_8),
.A2(n_63),
.B1(n_66),
.B2(n_149),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_9),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_9),
.A2(n_31),
.B1(n_33),
.B2(n_122),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_122),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_9),
.A2(n_63),
.B1(n_66),
.B2(n_122),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_183),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_183),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_10),
.A2(n_63),
.B1(n_66),
.B2(n_183),
.Y(n_268)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_12),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_12),
.B(n_30),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_33),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_12),
.A2(n_33),
.B(n_220),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_181),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_12),
.A2(n_60),
.B(n_63),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_12),
.B(n_89),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_12),
.A2(n_128),
.B1(n_129),
.B2(n_268),
.Y(n_270)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_15),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_75),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_319),
.Y(n_323)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_70),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_23),
.A2(n_121),
.B(n_123),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_23),
.A2(n_38),
.B1(n_121),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_23),
.A2(n_38),
.B1(n_148),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_24),
.A2(n_86),
.B(n_124),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_24),
.A2(n_30),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_25),
.B(n_33),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g180 ( 
.A(n_27),
.B(n_181),
.CON(n_180),
.SN(n_180)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_29),
.A2(n_31),
.B1(n_180),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_30),
.B(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_31),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_56)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_31),
.A2(n_47),
.A3(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_218)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_34),
.A2(n_38),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_57),
.B2(n_69),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_57),
.C(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_52),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_43),
.A2(n_77),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_44),
.A2(n_55),
.B1(n_79),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_44),
.A2(n_55),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_44),
.A2(n_55),
.B1(n_177),
.B2(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_44),
.A2(n_55),
.B1(n_205),
.B2(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_45),
.Y(n_219)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_45),
.B(n_48),
.Y(n_221)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_48),
.A2(n_61),
.B(n_181),
.C(n_247),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_52),
.A2(n_89),
.B(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_57),
.A2(n_69),
.B1(n_76),
.B2(n_317),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_67),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_58),
.A2(n_62),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_114),
.B(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_58),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_58),
.A2(n_67),
.B(n_132),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_58),
.A2(n_62),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_58),
.A2(n_155),
.B(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_58),
.A2(n_62),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_58),
.A2(n_62),
.B1(n_227),
.B2(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_113),
.B(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_62),
.B(n_181),
.Y(n_266)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_66),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_68),
.B(n_134),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.C(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_71),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_71),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_75),
.B(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_76),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_77),
.A2(n_80),
.B(n_90),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_312),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_333),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_166),
.B(n_311),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_150),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_99),
.B(n_150),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_125),
.C(n_136),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_100),
.A2(n_101),
.B1(n_125),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_115),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_117),
.C(n_119),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_103),
.B(n_112),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_110),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_104),
.A2(n_196),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_105),
.A2(n_111),
.B(n_141),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_105),
.A2(n_106),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_111),
.Y(n_110)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_106),
.Y(n_209)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_107),
.A2(n_128),
.B1(n_139),
.B2(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_129),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_110),
.A2(n_128),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_125),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_135),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_127),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_131),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_127),
.A2(n_160),
.B(n_163),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B(n_130),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_128),
.A2(n_209),
.B1(n_260),
.B2(n_268),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_129),
.B(n_181),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_131),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_133),
.B(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_136),
.B(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.C(n_146),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_137),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_142),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_145),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_164),
.B2(n_165),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_159),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_153),
.B(n_159),
.C(n_165),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B(n_158),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_158),
.B(n_314),
.C(n_320),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_158),
.A2(n_314),
.B1(n_315),
.B2(n_329),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_158),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_164),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_305),
.B(n_310),
.Y(n_166)
);

O2A1O1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_210),
.B(n_291),
.C(n_304),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_197),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_169),
.B(n_197),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_171),
.B(n_172),
.C(n_184),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_179),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_186),
.B(n_190),
.C(n_192),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_198),
.A2(n_199),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_203),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.C(n_208),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_208),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_290),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_283),
.B(n_289),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_238),
.B(n_282),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_229),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_214),
.B(n_229),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.C(n_225),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_215),
.A2(n_216),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_236),
.C(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_276),
.B(n_281),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_256),
.B(n_275),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_241),
.B(n_248),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_264),
.B(n_274),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_258),
.B(n_262),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_269),
.B(n_273),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_267),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_302),
.B2(n_303),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_299),
.C(n_303),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_302),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_313),
.B(n_322),
.Y(n_331)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_316),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_321),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);


endmodule