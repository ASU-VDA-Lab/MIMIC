module fake_ibex_772_n_4818 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_957, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_974, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_922, n_438, n_851, n_689, n_960, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_935, n_869, n_925, n_718, n_801, n_918, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_919, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4818);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_957;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_974;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_922;
input n_438;
input n_851;
input n_689;
input n_960;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4818;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_4557;
wire n_3150;
wire n_992;
wire n_4773;
wire n_4798;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4449;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_4688;
wire n_1110;
wire n_3610;
wire n_2607;
wire n_1382;
wire n_4615;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_4630;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_4632;
wire n_1080;
wire n_2290;
wire n_4607;
wire n_3750;
wire n_3838;
wire n_4514;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_4749;
wire n_1883;
wire n_1125;
wire n_4805;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_4550;
wire n_4668;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_2392;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_4731;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_4343;
wire n_4353;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4648;
wire n_3569;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4421;
wire n_4179;
wire n_4601;
wire n_3340;
wire n_4142;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_4785;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_1782;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_4585;
wire n_3168;
wire n_2396;
wire n_3904;
wire n_3135;
wire n_3440;
wire n_4378;
wire n_4169;
wire n_3729;
wire n_3175;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_4477;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_4654;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_4765;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_4418;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4708;
wire n_4592;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_4431;
wire n_1327;
wire n_2644;
wire n_4771;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_4652;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_4673;
wire n_3315;
wire n_3537;
wire n_4470;
wire n_4690;
wire n_1668;
wire n_3982;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_4781;
wire n_3724;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_4423;
wire n_4584;
wire n_1766;
wire n_3566;
wire n_3184;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_4578;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_3395;
wire n_3839;
wire n_4403;
wire n_1654;
wire n_3242;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_4526;
wire n_4808;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_4746;
wire n_1680;
wire n_2918;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_4304;
wire n_3976;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_4160;
wire n_4382;
wire n_3939;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_4450;
wire n_3969;
wire n_4467;
wire n_1081;
wire n_4437;
wire n_4801;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4491;
wire n_4672;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_4569;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_4723;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_4510;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_4312;
wire n_3699;
wire n_4567;
wire n_4556;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_4214;
wire n_1313;
wire n_3973;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_4430;
wire n_2260;
wire n_3977;
wire n_4724;
wire n_3722;
wire n_3125;
wire n_4769;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_4721;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_4806;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_4650;
wire n_1645;
wire n_3186;
wire n_4433;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_4428;
wire n_4784;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_4766;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_4563;
wire n_3809;
wire n_979;
wire n_4503;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4517;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3221;
wire n_3210;
wire n_3667;
wire n_1672;
wire n_4511;
wire n_1007;
wire n_2253;
wire n_4479;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_4182;
wire n_3858;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_4600;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_4422;
wire n_1219;
wire n_4513;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_4786;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_4735;
wire n_2189;
wire n_3548;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_4667;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_4610;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_4774;
wire n_1388;
wire n_2859;
wire n_4711;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_4799;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_4481;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_4809;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_4671;
wire n_1326;
wire n_4444;
wire n_1350;
wire n_4499;
wire n_3627;
wire n_2957;
wire n_4676;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_3777;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_4595;
wire n_2541;
wire n_4598;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_4553;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_4533;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_4174;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4455;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_4804;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4518;
wire n_4732;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_4480;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_4548;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_4535;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_4252;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4505;
wire n_3909;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_4577;
wire n_2292;
wire n_3573;
wire n_4604;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2444;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_4398;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_4522;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_4692;
wire n_4713;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_4476;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2646;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3963;
wire n_3800;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_4710;
wire n_1407;
wire n_3282;
wire n_4435;
wire n_4680;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_4649;
wire n_4755;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_4757;
wire n_1058;
wire n_4803;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_4693;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_1543;
wire n_4653;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_4568;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4573;
wire n_4549;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_4767;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_4623;
wire n_1041;
wire n_4700;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4523;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_4582;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_4489;
wire n_2236;
wire n_3455;
wire n_4758;
wire n_3957;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_4712;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_4419;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_1987;
wire n_4571;
wire n_1106;
wire n_1312;
wire n_4655;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_4725;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_4570;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_4494;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4681;
wire n_4122;
wire n_4542;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_4572;
wire n_1181;
wire n_3263;
wire n_4374;
wire n_4501;
wire n_1985;
wire n_1140;
wire n_4375;
wire n_3815;
wire n_4205;
wire n_1772;
wire n_4740;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_4768;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_1109;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_4813;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4469;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_4558;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_4460;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4504;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_4527;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_4608;
wire n_4485;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_1877;
wire n_4537;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_4793;
wire n_2468;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_4646;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_4462;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_4540;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_4490;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_2935;
wire n_3503;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1566;
wire n_1464;
wire n_4362;
wire n_3568;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_4626;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_4414;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_4706;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_4747;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_4791;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_4525;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_4443;
wire n_1682;
wire n_4151;
wire n_4625;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_4554;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_4424;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_4674;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4679;
wire n_4596;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4456;
wire n_4587;
wire n_4315;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_3578;
wire n_4734;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_4492;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_4500;
wire n_4559;
wire n_3797;
wire n_998;
wire n_1115;
wire n_1729;
wire n_1395;
wire n_2551;
wire n_4641;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4660;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_4664;
wire n_3829;
wire n_4579;
wire n_1864;
wire n_4624;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_4753;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4321;
wire n_4051;
wire n_4709;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_4552;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1599;
wire n_1400;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4640;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_4779;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4561;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_4642;
wire n_4764;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_4683;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_2185;
wire n_4141;
wire n_4614;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_4800;
wire n_2460;
wire n_2170;
wire n_4694;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_3383;
wire n_2884;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_3659;
wire n_3254;
wire n_4496;
wire n_4717;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4566;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_4719;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_4647;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4636;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4256;
wire n_1683;
wire n_1185;
wire n_4176;
wire n_3575;
wire n_4454;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_4278;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_4609;
wire n_1514;
wire n_2728;
wire n_3772;
wire n_4685;
wire n_2948;
wire n_4458;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_3657;
wire n_4716;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_4276;
wire n_4612;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_4185;
wire n_2422;
wire n_3902;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_4815;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_4441;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_2997;
wire n_3314;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_4704;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_4775;
wire n_4536;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_4633;
wire n_1950;
wire n_4497;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_4593;
wire n_3632;
wire n_3914;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_4512;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_4483;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4488;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4183;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_4814;
wire n_1694;
wire n_1458;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_4621;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3609;
wire n_3269;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4123;
wire n_3154;
wire n_4000;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_4619;
wire n_4645;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_4007;
wire n_3960;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_4707;
wire n_1754;
wire n_4286;
wire n_4429;
wire n_3048;
wire n_3686;
wire n_1991;
wire n_1177;
wire n_1025;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_4695;
wire n_982;
wire n_4438;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_4802;
wire n_3912;
wire n_3778;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_4816;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_4638;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_4498;
wire n_3265;
wire n_2240;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_4750;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2555;
wire n_2639;
wire n_2330;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_4745;
wire n_3057;
wire n_2143;
wire n_4319;
wire n_2410;
wire n_4057;
wire n_3760;
wire n_4637;
wire n_1396;
wire n_4792;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_4373;
wire n_2351;
wire n_2437;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_4543;
wire n_4466;
wire n_2688;
wire n_2881;
wire n_4643;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_4603;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4212;
wire n_4022;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_3162;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_4436;
wire n_4599;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_4697;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_4538;
wire n_3096;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_4783;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_4730;
wire n_1238;
wire n_1415;
wire n_4616;
wire n_3959;
wire n_3743;
wire n_4760;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_4763;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_4434;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_4720;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_4586;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_4583;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_4622;
wire n_3273;
wire n_4367;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_4715;
wire n_1630;
wire n_3408;
wire n_4475;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_4588;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_4698;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_4741;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_4440;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3604;
wire n_1838;
wire n_3540;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_4739;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_4529;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2576;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4162;
wire n_4111;
wire n_4408;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_4575;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_4759;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_4620;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_4666;
wire n_4770;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_4439;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_4722;
wire n_1530;
wire n_4200;
wire n_3215;
wire n_3413;
wire n_4580;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_4565;
wire n_1088;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_4663;
wire n_2471;
wire n_4581;
wire n_1288;
wire n_4058;
wire n_4487;
wire n_4618;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4519;
wire n_4148;
wire n_1622;
wire n_2757;
wire n_4611;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_4541;
wire n_4515;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_4530;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_4463;
wire n_4591;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_4670;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_4265;
wire n_3062;
wire n_4524;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4628;
wire n_4017;
wire n_1547;
wire n_1542;
wire n_1586;
wire n_1362;
wire n_3497;
wire n_4696;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_3368;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_4597;
wire n_4778;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_4789;
wire n_1951;
wire n_1330;
wire n_4574;
wire n_4659;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_4748;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_2593;
wire n_3899;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_4729;
wire n_1798;
wire n_4555;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_4761;
wire n_3549;
wire n_4751;
wire n_4562;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3972;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_4453;
wire n_1098;
wire n_4474;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_3173;
wire n_2872;
wire n_3102;
wire n_2790;
wire n_4281;
wire n_4345;
wire n_4478;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_4473;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_4464;
wire n_3761;
wire n_2526;
wire n_4794;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_4675;
wire n_3083;
wire n_2083;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_4605;
wire n_4737;
wire n_3844;
wire n_2207;
wire n_4210;
wire n_4752;
wire n_4049;
wire n_2044;
wire n_4546;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1572;
wire n_1635;
wire n_4810;
wire n_3149;
wire n_2827;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_4432;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1912;
wire n_1297;
wire n_1369;
wire n_3143;
wire n_1734;
wire n_3655;
wire n_3543;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4461;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_3042;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_4516;
wire n_2913;
wire n_2491;
wire n_4686;
wire n_1529;
wire n_1824;
wire n_1381;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_4682;
wire n_4528;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_4502;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_4705;
wire n_4811;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_4471;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_4733;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_4547;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_4684;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_4807;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_4482;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_4493;
wire n_4797;
wire n_4738;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_980;
wire n_1193;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_1074;
wire n_3557;
wire n_3380;
wire n_3207;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_1180;
wire n_1462;
wire n_4657;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4718;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1904;
wire n_1262;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_4634;
wire n_4644;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_1022;
wire n_4412;
wire n_4796;
wire n_1760;
wire n_4560;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3737;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_4472;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_4639;
wire n_3636;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_4787;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_4635;
wire n_4521;
wire n_1230;
wire n_4459;
wire n_1516;
wire n_1027;
wire n_4551;
wire n_3893;
wire n_4484;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_2148;
wire n_2104;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_4354;
wire n_4448;
wire n_3938;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_4532;
wire n_4727;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_4701;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4627;
wire n_4743;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_4726;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_2802;
wire n_3052;
wire n_3189;
wire n_4544;
wire n_4728;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_2961;
wire n_4589;
wire n_1915;
wire n_2836;
wire n_3924;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_4631;
wire n_3283;
wire n_4468;
wire n_1736;
wire n_4617;
wire n_4442;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_4689;
wire n_4772;
wire n_3613;
wire n_1383;
wire n_990;
wire n_4108;
wire n_1968;
wire n_3675;
wire n_2057;
wire n_4594;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_4613;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_4629;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_4539;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_4776;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_4702;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_4486;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_4506;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_1551;
wire n_4153;
wire n_3793;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_4817;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_4780;
wire n_4327;
wire n_2656;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_4465;
wire n_1355;
wire n_3691;
wire n_4452;
wire n_2544;
wire n_3193;
wire n_4534;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_4590;
wire n_2915;
wire n_1579;
wire n_4446;
wire n_1280;
wire n_4602;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_4576;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_4606;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_4782;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_4777;
wire n_3851;
wire n_4508;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_3654;
wire n_4425;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_4703;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_4691;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_4662;
wire n_2658;

INVx2_ASAP7_75t_L g979 ( 
.A(n_647),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_173),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_451),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_44),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_946),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_842),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_899),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_829),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_937),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_582),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_635),
.Y(n_989)
);

BUFx10_ASAP7_75t_L g990 ( 
.A(n_417),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_953),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_921),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_855),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_929),
.Y(n_994)
);

CKINVDCx16_ASAP7_75t_R g995 ( 
.A(n_365),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_420),
.Y(n_996)
);

CKINVDCx16_ASAP7_75t_R g997 ( 
.A(n_744),
.Y(n_997)
);

BUFx8_ASAP7_75t_SL g998 ( 
.A(n_935),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_905),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_430),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_917),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_915),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_948),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_756),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_529),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_901),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_484),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_967),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_745),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_641),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_909),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_569),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_274),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_427),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_549),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_87),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_908),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_665),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_614),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_569),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_881),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_424),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_155),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_954),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_930),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_692),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_974),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_907),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_303),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_311),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_678),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_545),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_225),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_894),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_87),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_210),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_888),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_438),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_707),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_904),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_936),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_653),
.Y(n_1042)
);

BUFx2_ASAP7_75t_SL g1043 ( 
.A(n_961),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_110),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_455),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_115),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_912),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_386),
.Y(n_1048)
);

INVxp67_ASAP7_75t_SL g1049 ( 
.A(n_253),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_234),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_669),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_66),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_42),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_487),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_298),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_609),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_966),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_259),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_658),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_24),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_641),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_147),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_971),
.Y(n_1063)
);

CKINVDCx20_ASAP7_75t_R g1064 ( 
.A(n_926),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_252),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_244),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_113),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_574),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_827),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_958),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_923),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_104),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_308),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_909),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_101),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_115),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_395),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_753),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_922),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_890),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_889),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_718),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_39),
.Y(n_1083)
);

BUFx10_ASAP7_75t_L g1084 ( 
.A(n_128),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_327),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_745),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

CKINVDCx16_ASAP7_75t_R g1088 ( 
.A(n_949),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_769),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_397),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_306),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_854),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_373),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_740),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_264),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_465),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_211),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_760),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_15),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_352),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_528),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_550),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_314),
.Y(n_1103)
);

BUFx3_ASAP7_75t_L g1104 ( 
.A(n_957),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_758),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_903),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_660),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_263),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_754),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_689),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_696),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_314),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_65),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_593),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_167),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_408),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_330),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_259),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_919),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_902),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_810),
.Y(n_1121)
);

CKINVDCx20_ASAP7_75t_R g1122 ( 
.A(n_939),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_446),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_90),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_658),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_249),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_180),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_249),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_14),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_900),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_215),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_548),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_303),
.Y(n_1133)
);

BUFx5_ASAP7_75t_L g1134 ( 
.A(n_934),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_5),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_435),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_206),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_598),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_571),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_898),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_254),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_298),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_248),
.Y(n_1143)
);

BUFx10_ASAP7_75t_L g1144 ( 
.A(n_121),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_504),
.Y(n_1145)
);

BUFx10_ASAP7_75t_L g1146 ( 
.A(n_584),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_316),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_707),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_716),
.Y(n_1149)
);

INVx1_ASAP7_75t_SL g1150 ( 
.A(n_358),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_244),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_405),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_300),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_856),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_844),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_940),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_461),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_812),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_364),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_227),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_176),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_174),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_731),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_97),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_814),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_623),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_674),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_366),
.Y(n_1168)
);

CKINVDCx14_ASAP7_75t_R g1169 ( 
.A(n_796),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_575),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_416),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_2),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_437),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_95),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_898),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_267),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_911),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_920),
.Y(n_1178)
);

BUFx5_ASAP7_75t_L g1179 ( 
.A(n_145),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_610),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_557),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_945),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_509),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_901),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_321),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_36),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_410),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_747),
.Y(n_1188)
);

CKINVDCx20_ASAP7_75t_R g1189 ( 
.A(n_394),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_513),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_574),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_634),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_268),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_197),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_561),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_968),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_771),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_777),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_67),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_524),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_842),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_740),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_71),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_623),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_752),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_665),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_941),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_897),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_944),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_428),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_689),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_20),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_804),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_807),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_343),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_925),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_249),
.Y(n_1217)
);

CKINVDCx16_ASAP7_75t_R g1218 ( 
.A(n_950),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_750),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_833),
.Y(n_1220)
);

BUFx10_ASAP7_75t_L g1221 ( 
.A(n_262),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_650),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_88),
.Y(n_1223)
);

BUFx10_ASAP7_75t_L g1224 ( 
.A(n_418),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_24),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_451),
.Y(n_1226)
);

INVx1_ASAP7_75t_SL g1227 ( 
.A(n_235),
.Y(n_1227)
);

BUFx3_ASAP7_75t_L g1228 ( 
.A(n_918),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_896),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_21),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_966),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_925),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_895),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_797),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_963),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_192),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_533),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_591),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_816),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_412),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_761),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_140),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_109),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_605),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_773),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_943),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_118),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_525),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_483),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_58),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_916),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_392),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_688),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_682),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_759),
.Y(n_1255)
);

BUFx10_ASAP7_75t_L g1256 ( 
.A(n_710),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_886),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_381),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_698),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_247),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_517),
.Y(n_1261)
);

INVx1_ASAP7_75t_SL g1262 ( 
.A(n_932),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_572),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_112),
.Y(n_1264)
);

BUFx2_ASAP7_75t_SL g1265 ( 
.A(n_724),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_573),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_219),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_394),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_725),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_917),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_528),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_345),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_779),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_737),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_820),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_157),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_52),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_526),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_30),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_924),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_187),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_406),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_799),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_906),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_713),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_135),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_294),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_748),
.Y(n_1288)
);

CKINVDCx20_ASAP7_75t_R g1289 ( 
.A(n_967),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_813),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_929),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_113),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_423),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_613),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_489),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_756),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_877),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_956),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_819),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_94),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_410),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_970),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_928),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_108),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_956),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_111),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_108),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_87),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_521),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_213),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_947),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_843),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_124),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_960),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_915),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_181),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_965),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_910),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_301),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_231),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_307),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_426),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_178),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_34),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_148),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_797),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_655),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_165),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_782),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_188),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_920),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_409),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_46),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_404),
.Y(n_1334)
);

BUFx2_ASAP7_75t_L g1335 ( 
.A(n_914),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_682),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_964),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_219),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_633),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_155),
.Y(n_1340)
);

CKINVDCx16_ASAP7_75t_R g1341 ( 
.A(n_536),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_7),
.Y(n_1342)
);

CKINVDCx20_ASAP7_75t_R g1343 ( 
.A(n_31),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_865),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_51),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_959),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_811),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_972),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_285),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_146),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_412),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_601),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_647),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_244),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_141),
.Y(n_1355)
);

BUFx2_ASAP7_75t_L g1356 ( 
.A(n_119),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_199),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_666),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_318),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_594),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_325),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_972),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_942),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_951),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_364),
.Y(n_1365)
);

BUFx10_ASAP7_75t_L g1366 ( 
.A(n_266),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_34),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_864),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_962),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_701),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_60),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_147),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_263),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_892),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_480),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_110),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_741),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_685),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_156),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_342),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_390),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_695),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_179),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_434),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_253),
.Y(n_1385)
);

BUFx5_ASAP7_75t_L g1386 ( 
.A(n_459),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_323),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_644),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_664),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_523),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_653),
.Y(n_1391)
);

BUFx6f_ASAP7_75t_L g1392 ( 
.A(n_965),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_166),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_453),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_973),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_97),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_130),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_779),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_188),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_695),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_509),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_220),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_281),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_397),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_465),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_969),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_892),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_713),
.Y(n_1408)
);

INVxp33_ASAP7_75t_R g1409 ( 
.A(n_574),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_607),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_750),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_938),
.Y(n_1412)
);

CKINVDCx14_ASAP7_75t_R g1413 ( 
.A(n_183),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_192),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_140),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_927),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_836),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_130),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_48),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_177),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_177),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_787),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_162),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_751),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_518),
.Y(n_1425)
);

INVx1_ASAP7_75t_SL g1426 ( 
.A(n_690),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_198),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_636),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_921),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_969),
.Y(n_1430)
);

BUFx8_ASAP7_75t_SL g1431 ( 
.A(n_354),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_749),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_135),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_931),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_761),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_415),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_163),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_501),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_819),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_891),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_893),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_280),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_705),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_448),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_454),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_931),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_232),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_913),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_343),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_539),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_807),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_456),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_608),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_492),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_43),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_467),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_610),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_133),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_734),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_809),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_335),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_908),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_342),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_214),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_526),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_513),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_537),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_314),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_156),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_7),
.Y(n_1470)
);

CKINVDCx16_ASAP7_75t_R g1471 ( 
.A(n_542),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_515),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_294),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_107),
.Y(n_1474)
);

INVx1_ASAP7_75t_SL g1475 ( 
.A(n_381),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_674),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_747),
.Y(n_1477)
);

CKINVDCx14_ASAP7_75t_R g1478 ( 
.A(n_652),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_306),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_207),
.Y(n_1480)
);

BUFx5_ASAP7_75t_L g1481 ( 
.A(n_155),
.Y(n_1481)
);

BUFx2_ASAP7_75t_SL g1482 ( 
.A(n_952),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_18),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_757),
.Y(n_1484)
);

BUFx5_ASAP7_75t_L g1485 ( 
.A(n_496),
.Y(n_1485)
);

CKINVDCx16_ASAP7_75t_R g1486 ( 
.A(n_357),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_310),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_237),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_955),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_995),
.B(n_0),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1413),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1413),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1478),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1010),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1048),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1023),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1051),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1431),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1026),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1083),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1014),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1014),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1335),
.B(n_0),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1328),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1380),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1022),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1455),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1133),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_1169),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1039),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1110),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1324),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1133),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1169),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_998),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1160),
.Y(n_1516)
);

BUFx2_ASAP7_75t_SL g1517 ( 
.A(n_990),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1356),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1048),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1341),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1379),
.Y(n_1521)
);

INVxp67_ASAP7_75t_SL g1522 ( 
.A(n_1136),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1471),
.Y(n_1523)
);

INVxp33_ASAP7_75t_SL g1524 ( 
.A(n_1487),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1486),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_980),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_988),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_989),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_981),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_982),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_996),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1019),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1000),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_1135),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1135),
.Y(n_1535)
);

CKINVDCx5p33_ASAP7_75t_R g1536 ( 
.A(n_1005),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1136),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1030),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1134),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1031),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1189),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1033),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1042),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1044),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1050),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1007),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1104),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1189),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1058),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1075),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1076),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1191),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1191),
.Y(n_1553)
);

CKINVDCx14_ASAP7_75t_R g1554 ( 
.A(n_990),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1097),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1266),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1100),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1108),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1114),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1012),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1117),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1213),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1013),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1016),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1118),
.Y(n_1565)
);

CKINVDCx20_ASAP7_75t_R g1566 ( 
.A(n_1276),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1134),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1018),
.Y(n_1568)
);

INVxp67_ASAP7_75t_SL g1569 ( 
.A(n_1170),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1123),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_L g1571 ( 
.A(n_1311),
.B(n_1182),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1029),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1134),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_1276),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1364),
.B(n_2),
.Y(n_1575)
);

INVxp33_ASAP7_75t_SL g1576 ( 
.A(n_1032),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1336),
.Y(n_1577)
);

CKINVDCx5p33_ASAP7_75t_R g1578 ( 
.A(n_1035),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1125),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1036),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1170),
.Y(n_1581)
);

BUFx2_ASAP7_75t_L g1582 ( 
.A(n_1263),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1038),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1126),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1336),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1129),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1134),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_997),
.B(n_1),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1132),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_1045),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1138),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1263),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1046),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1147),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_1052),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1157),
.Y(n_1596)
);

CKINVDCx20_ASAP7_75t_R g1597 ( 
.A(n_1343),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1466),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1547),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1581),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1582),
.Y(n_1601)
);

NOR2xp67_ASAP7_75t_L g1602 ( 
.A(n_1499),
.B(n_1225),
.Y(n_1602)
);

BUFx2_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

AND2x6_ASAP7_75t_L g1604 ( 
.A(n_1510),
.B(n_1466),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1537),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1506),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1537),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1576),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1498),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1539),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1054),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1512),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1567),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1526),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1491),
.B(n_1492),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1527),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1592),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_1528),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1533),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1494),
.Y(n_1621)
);

CKINVDCx20_ASAP7_75t_R g1622 ( 
.A(n_1501),
.Y(n_1622)
);

CKINVDCx20_ASAP7_75t_R g1623 ( 
.A(n_1502),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1508),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1587),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1496),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1536),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1495),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1055),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_1546),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1511),
.Y(n_1631)
);

CKINVDCx16_ASAP7_75t_R g1632 ( 
.A(n_1517),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1560),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1497),
.Y(n_1634)
);

BUFx6f_ASAP7_75t_L g1635 ( 
.A(n_1495),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1563),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1522),
.Y(n_1637)
);

CKINVDCx16_ASAP7_75t_R g1638 ( 
.A(n_1513),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1529),
.A2(n_1020),
.B(n_979),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1564),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1569),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1500),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1568),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1495),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1524),
.B(n_1056),
.Y(n_1645)
);

CKINVDCx20_ASAP7_75t_R g1646 ( 
.A(n_1534),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1535),
.Y(n_1647)
);

INVx6_ASAP7_75t_L g1648 ( 
.A(n_1575),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1504),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1505),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1572),
.Y(n_1651)
);

AND2x2_ASAP7_75t_SL g1652 ( 
.A(n_1562),
.B(n_1088),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1507),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1530),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_R g1655 ( 
.A(n_1515),
.B(n_1218),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1531),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1532),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1538),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1540),
.Y(n_1659)
);

CKINVDCx20_ASAP7_75t_R g1660 ( 
.A(n_1541),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1519),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1519),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1519),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1578),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1580),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1542),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1543),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1544),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1545),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1583),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1590),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1593),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1549),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1516),
.B(n_1207),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1550),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1595),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1551),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1520),
.Y(n_1678)
);

NOR2xp67_ASAP7_75t_L g1679 ( 
.A(n_1518),
.B(n_1162),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1523),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1525),
.Y(n_1681)
);

BUFx6f_ASAP7_75t_L g1682 ( 
.A(n_1519),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1555),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1557),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1558),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1548),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1552),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1521),
.B(n_990),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_1553),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1556),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1559),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1561),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1571),
.B(n_1207),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1565),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1570),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1509),
.B(n_1059),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1566),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1579),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1584),
.A2(n_1020),
.B(n_979),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1574),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1586),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1589),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1490),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_SL g1704 ( 
.A(n_1493),
.B(n_1179),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1591),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1594),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1596),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1577),
.Y(n_1708)
);

INVx3_ASAP7_75t_L g1709 ( 
.A(n_1514),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1585),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_1597),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1503),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1588),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1581),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1491),
.B(n_1179),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1495),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1501),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1581),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1554),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1554),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1581),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1554),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1554),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1554),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1491),
.B(n_1179),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1554),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1494),
.B(n_1060),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1547),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1495),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1547),
.Y(n_1730)
);

BUFx6f_ASAP7_75t_L g1731 ( 
.A(n_1495),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1554),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1554),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1554),
.B(n_1062),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1501),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1581),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1547),
.Y(n_1737)
);

CKINVDCx16_ASAP7_75t_R g1738 ( 
.A(n_1554),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1581),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1581),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1495),
.Y(n_1741)
);

CKINVDCx5p33_ASAP7_75t_R g1742 ( 
.A(n_1554),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_R g1743 ( 
.A(n_1554),
.B(n_1066),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1547),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1554),
.B(n_1072),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1554),
.B(n_1073),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1581),
.Y(n_1747)
);

BUFx6f_ASAP7_75t_L g1748 ( 
.A(n_1495),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1554),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1501),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_1554),
.Y(n_1751)
);

BUFx6f_ASAP7_75t_L g1752 ( 
.A(n_1495),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1554),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1554),
.B(n_1077),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_1501),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1547),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1510),
.B(n_1228),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1554),
.Y(n_1758)
);

AND2x6_ASAP7_75t_L g1759 ( 
.A(n_1510),
.B(n_1228),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1554),
.B(n_1015),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1554),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1581),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1581),
.Y(n_1763)
);

CKINVDCx20_ASAP7_75t_R g1764 ( 
.A(n_1501),
.Y(n_1764)
);

CKINVDCx20_ASAP7_75t_R g1765 ( 
.A(n_1501),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1547),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1554),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1581),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1581),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1547),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1501),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1581),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1554),
.B(n_1085),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1554),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1581),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1547),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1703),
.B(n_1179),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1713),
.A2(n_1090),
.B1(n_1096),
.B2(n_1091),
.Y(n_1778)
);

INVx4_ASAP7_75t_SL g1779 ( 
.A(n_1604),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1606),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1639),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1724),
.B(n_1343),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1657),
.B(n_1179),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1701),
.B(n_1386),
.Y(n_1784)
);

INVx5_ASAP7_75t_L g1785 ( 
.A(n_1738),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1642),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1611),
.B(n_1386),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1699),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1631),
.B(n_1099),
.Y(n_1789)
);

OAI22x1_ASAP7_75t_L g1790 ( 
.A1(n_1686),
.A2(n_1409),
.B1(n_1360),
.B2(n_1382),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1726),
.B(n_1093),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1653),
.Y(n_1792)
);

INVx4_ASAP7_75t_L g1793 ( 
.A(n_1732),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1626),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1612),
.B(n_1760),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1634),
.Y(n_1796)
);

INVx3_ASAP7_75t_L g1797 ( 
.A(n_1632),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1719),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1608),
.A2(n_1360),
.B1(n_1382),
.B2(n_1352),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1720),
.B(n_1352),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1749),
.B(n_1015),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1722),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1743),
.Y(n_1803)
);

INVx2_ASAP7_75t_SL g1804 ( 
.A(n_1648),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1676),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1649),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1645),
.B(n_1095),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1650),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1774),
.B(n_1652),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1629),
.B(n_1605),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1599),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_SL g1812 ( 
.A1(n_1648),
.A2(n_1102),
.B1(n_1103),
.B2(n_1101),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_SL g1813 ( 
.A(n_1688),
.B(n_1015),
.Y(n_1813)
);

INVx2_ASAP7_75t_SL g1814 ( 
.A(n_1604),
.Y(n_1814)
);

OAI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1614),
.A2(n_1387),
.B1(n_1061),
.B2(n_1067),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_L g1816 ( 
.A1(n_1637),
.A2(n_1167),
.B1(n_1168),
.B2(n_1166),
.Y(n_1816)
);

BUFx6f_ASAP7_75t_L g1817 ( 
.A(n_1723),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1733),
.Y(n_1818)
);

OR2x2_ASAP7_75t_SL g1819 ( 
.A(n_1638),
.B(n_983),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1607),
.B(n_1386),
.Y(n_1820)
);

OR2x6_ASAP7_75t_L g1821 ( 
.A(n_1633),
.B(n_1043),
.Y(n_1821)
);

AND2x6_ASAP7_75t_L g1822 ( 
.A(n_1641),
.B(n_1053),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1691),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1691),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1617),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_SL g1826 ( 
.A(n_1734),
.B(n_1084),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1745),
.B(n_1111),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1618),
.B(n_1386),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1621),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1742),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1751),
.Y(n_1831)
);

INVx1_ASAP7_75t_SL g1832 ( 
.A(n_1619),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_L g1833 ( 
.A(n_1696),
.B(n_1113),
.C(n_1112),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1746),
.B(n_1084),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1656),
.A2(n_1174),
.B1(n_1180),
.B2(n_1173),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1754),
.B(n_1115),
.Y(n_1836)
);

INVx3_ASAP7_75t_L g1837 ( 
.A(n_1756),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1654),
.B(n_1386),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1659),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1600),
.A2(n_1116),
.B1(n_1127),
.B2(n_1124),
.Y(n_1840)
);

INVx5_ASAP7_75t_L g1841 ( 
.A(n_1770),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1773),
.B(n_1139),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1658),
.B(n_1386),
.Y(n_1843)
);

BUFx6f_ASAP7_75t_L g1844 ( 
.A(n_1753),
.Y(n_1844)
);

CKINVDCx5p33_ASAP7_75t_R g1845 ( 
.A(n_1758),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1761),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1602),
.B(n_1640),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1666),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1601),
.B(n_1128),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1669),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1728),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1620),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1714),
.B(n_1131),
.Y(n_1853)
);

INVx5_ASAP7_75t_L g1854 ( 
.A(n_1759),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1667),
.B(n_1386),
.Y(n_1855)
);

AND2x6_ASAP7_75t_L g1856 ( 
.A(n_1709),
.B(n_1107),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1718),
.A2(n_1141),
.B1(n_1142),
.B2(n_1137),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1675),
.A2(n_1187),
.B1(n_1193),
.B2(n_1183),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1668),
.B(n_1481),
.Y(n_1859)
);

INVx3_ASAP7_75t_L g1860 ( 
.A(n_1730),
.Y(n_1860)
);

NAND2xp33_ASAP7_75t_SL g1861 ( 
.A(n_1767),
.B(n_1143),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1677),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1622),
.Y(n_1863)
);

INVx6_ASAP7_75t_L g1864 ( 
.A(n_1674),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1721),
.B(n_1150),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1736),
.B(n_1139),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1673),
.B(n_1481),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1739),
.A2(n_1145),
.B1(n_1151),
.B2(n_1148),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1685),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1740),
.B(n_1153),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1623),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1747),
.B(n_1144),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1683),
.B(n_1481),
.Y(n_1873)
);

AND2x6_ASAP7_75t_L g1874 ( 
.A(n_1684),
.B(n_1190),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1737),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1694),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1762),
.B(n_1065),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1744),
.Y(n_1878)
);

BUFx3_ASAP7_75t_L g1879 ( 
.A(n_1627),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1766),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1763),
.B(n_1768),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1692),
.B(n_1481),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1769),
.B(n_1068),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1698),
.B(n_1144),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1759),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1695),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1702),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1705),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1706),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1707),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1674),
.A2(n_1206),
.B1(n_1210),
.B2(n_1203),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1776),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1772),
.B(n_1775),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1757),
.Y(n_1894)
);

OR2x6_ASAP7_75t_L g1895 ( 
.A(n_1615),
.B(n_1265),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1610),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1630),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1727),
.B(n_1679),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1757),
.B(n_1481),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1693),
.B(n_1485),
.Y(n_1900)
);

BUFx2_ASAP7_75t_L g1901 ( 
.A(n_1636),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1704),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1613),
.Y(n_1903)
);

INVxp67_ASAP7_75t_SL g1904 ( 
.A(n_1616),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1715),
.B(n_1159),
.Y(n_1905)
);

INVx4_ASAP7_75t_L g1906 ( 
.A(n_1643),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1625),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1725),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1651),
.B(n_1144),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1664),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1665),
.B(n_1485),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1670),
.A2(n_1215),
.B1(n_1217),
.B2(n_1211),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1671),
.Y(n_1913)
);

INVx4_ASAP7_75t_L g1914 ( 
.A(n_1672),
.Y(n_1914)
);

INVx3_ASAP7_75t_L g1915 ( 
.A(n_1678),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1680),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1681),
.A2(n_1226),
.B1(n_1236),
.B2(n_1223),
.Y(n_1917)
);

NAND2xp33_ASAP7_75t_L g1918 ( 
.A(n_1655),
.B(n_1485),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1687),
.B(n_1161),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1644),
.Y(n_1920)
);

BUFx10_ASAP7_75t_L g1921 ( 
.A(n_1609),
.Y(n_1921)
);

NOR3xp33_ASAP7_75t_L g1922 ( 
.A(n_1700),
.B(n_1049),
.C(n_1227),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1710),
.B(n_1164),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1644),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1661),
.B(n_1485),
.Y(n_1925)
);

BUFx10_ASAP7_75t_L g1926 ( 
.A(n_1624),
.Y(n_1926)
);

BUFx6f_ASAP7_75t_L g1927 ( 
.A(n_1628),
.Y(n_1927)
);

INVxp67_ASAP7_75t_SL g1928 ( 
.A(n_1646),
.Y(n_1928)
);

INVx3_ASAP7_75t_L g1929 ( 
.A(n_1635),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1661),
.B(n_1485),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1647),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1660),
.B(n_1146),
.Y(n_1932)
);

BUFx6f_ASAP7_75t_L g1933 ( 
.A(n_1716),
.Y(n_1933)
);

BUFx4f_ASAP7_75t_L g1934 ( 
.A(n_1689),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1690),
.B(n_1171),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1662),
.Y(n_1936)
);

INVx4_ASAP7_75t_SL g1937 ( 
.A(n_1662),
.Y(n_1937)
);

AOI22xp33_ASAP7_75t_L g1938 ( 
.A1(n_1731),
.A2(n_1240),
.B1(n_1242),
.B2(n_1237),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1697),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_L g1940 ( 
.A1(n_1663),
.A2(n_1253),
.B1(n_1260),
.B2(n_1252),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1663),
.Y(n_1941)
);

NAND2xp33_ASAP7_75t_L g1942 ( 
.A(n_1682),
.B(n_1134),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1682),
.B(n_1172),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1682),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1729),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1708),
.B(n_1176),
.Y(n_1946)
);

OR2x2_ASAP7_75t_L g1947 ( 
.A(n_1711),
.B(n_1261),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1729),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1717),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1741),
.B(n_1146),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1741),
.Y(n_1951)
);

NAND3xp33_ASAP7_75t_SL g1952 ( 
.A(n_1735),
.B(n_1454),
.C(n_1442),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1750),
.B(n_1152),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1755),
.B(n_1181),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1748),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1748),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1752),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1764),
.A2(n_1186),
.B1(n_1194),
.B2(n_1185),
.Y(n_1958)
);

AND2x6_ASAP7_75t_L g1959 ( 
.A(n_1752),
.B(n_1192),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1771),
.B(n_1195),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1765),
.A2(n_1277),
.B1(n_1282),
.B2(n_1272),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1703),
.B(n_1200),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1606),
.Y(n_1963)
);

INVx4_ASAP7_75t_L g1964 ( 
.A(n_1603),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1760),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1703),
.B(n_1204),
.Y(n_1966)
);

INVx4_ASAP7_75t_SL g1967 ( 
.A(n_1604),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1642),
.Y(n_1968)
);

BUFx6f_ASAP7_75t_L g1969 ( 
.A(n_1603),
.Y(n_1969)
);

AO22x2_ASAP7_75t_L g1970 ( 
.A1(n_1703),
.A2(n_1482),
.B1(n_1375),
.B2(n_1403),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1703),
.B(n_1212),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1743),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1603),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1642),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1606),
.B(n_1152),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1642),
.Y(n_1976)
);

INVx3_ASAP7_75t_L g1977 ( 
.A(n_1632),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1603),
.Y(n_1978)
);

OAI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1606),
.A2(n_1461),
.B1(n_1122),
.B2(n_1175),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1603),
.Y(n_1980)
);

INVx5_ASAP7_75t_L g1981 ( 
.A(n_1738),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1632),
.Y(n_1982)
);

INVx1_ASAP7_75t_SL g1983 ( 
.A(n_1606),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1760),
.B(n_1221),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1642),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1760),
.B(n_1221),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1606),
.Y(n_1987)
);

AND2x4_ASAP7_75t_L g1988 ( 
.A(n_1603),
.B(n_983),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1642),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1642),
.Y(n_1990)
);

BUFx6f_ASAP7_75t_L g1991 ( 
.A(n_1603),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1703),
.A2(n_1243),
.B1(n_1244),
.B2(n_1238),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1760),
.B(n_1221),
.Y(n_1993)
);

AOI22xp33_ASAP7_75t_L g1994 ( 
.A1(n_1712),
.A2(n_1286),
.B1(n_1293),
.B2(n_1287),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1603),
.B(n_1122),
.Y(n_1995)
);

BUFx10_ASAP7_75t_L g1996 ( 
.A(n_1719),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1703),
.B(n_1247),
.Y(n_1997)
);

BUFx10_ASAP7_75t_L g1998 ( 
.A(n_1719),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1807),
.B(n_1248),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1780),
.B(n_1249),
.Y(n_2000)
);

BUFx3_ASAP7_75t_L g2001 ( 
.A(n_1785),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1805),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1822),
.A2(n_1366),
.B1(n_1224),
.B2(n_1254),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1807),
.B(n_1250),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1781),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1983),
.B(n_1258),
.Y(n_2006)
);

CKINVDCx14_ASAP7_75t_R g2007 ( 
.A(n_1863),
.Y(n_2007)
);

BUFx6f_ASAP7_75t_SL g2008 ( 
.A(n_1926),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1822),
.A2(n_1366),
.B1(n_1268),
.B2(n_1271),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_SL g2010 ( 
.A(n_1906),
.B(n_1175),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1962),
.B(n_1267),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1987),
.B(n_1963),
.Y(n_2012)
);

OR2x6_ASAP7_75t_L g2013 ( 
.A(n_1791),
.B(n_992),
.Y(n_2013)
);

OAI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1788),
.A2(n_1308),
.B(n_1307),
.Y(n_2014)
);

OR2x6_ASAP7_75t_L g2015 ( 
.A(n_1914),
.B(n_992),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1887),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1825),
.B(n_1178),
.Y(n_2017)
);

BUFx4f_ASAP7_75t_L g2018 ( 
.A(n_1798),
.Y(n_2018)
);

NAND2xp33_ASAP7_75t_L g2019 ( 
.A(n_1874),
.B(n_1279),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1969),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1971),
.B(n_1281),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1969),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1965),
.B(n_1292),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1779),
.B(n_991),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_SL g2025 ( 
.A(n_1854),
.B(n_1294),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1888),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1795),
.B(n_1295),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1865),
.B(n_1366),
.Y(n_2028)
);

CKINVDCx14_ASAP7_75t_R g2029 ( 
.A(n_1871),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_L g2030 ( 
.A(n_1919),
.B(n_1923),
.C(n_1836),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1822),
.A2(n_1301),
.B1(n_1304),
.B2(n_1300),
.Y(n_2031)
);

O2A1O1Ixp5_ASAP7_75t_L g2032 ( 
.A1(n_1911),
.A2(n_1230),
.B(n_1320),
.C(n_1199),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1975),
.B(n_1306),
.Y(n_2033)
);

AOI22xp5_ASAP7_75t_L g2034 ( 
.A1(n_1866),
.A2(n_1309),
.B1(n_1316),
.B2(n_1313),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1779),
.B(n_993),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1872),
.A2(n_1321),
.B1(n_1325),
.B2(n_1323),
.Y(n_2036)
);

INVx2_ASAP7_75t_SL g2037 ( 
.A(n_1978),
.Y(n_2037)
);

INVx2_ASAP7_75t_SL g2038 ( 
.A(n_1978),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1889),
.Y(n_2039)
);

BUFx2_ASAP7_75t_L g2040 ( 
.A(n_1973),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1992),
.A2(n_1330),
.B1(n_1334),
.B2(n_1332),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1890),
.Y(n_2042)
);

NOR2x1p5_ASAP7_75t_L g2043 ( 
.A(n_1952),
.B(n_1338),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1997),
.B(n_1476),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1777),
.B(n_1479),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1847),
.B(n_1342),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1810),
.B(n_1488),
.Y(n_2047)
);

NOR2xp33_ASAP7_75t_L g2048 ( 
.A(n_1881),
.B(n_1865),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1808),
.B(n_1345),
.Y(n_2049)
);

OAI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_1881),
.A2(n_1229),
.B1(n_1269),
.B2(n_1178),
.Y(n_2050)
);

O2A1O1Ixp33_ASAP7_75t_L g2051 ( 
.A1(n_1812),
.A2(n_1426),
.B(n_1456),
.C(n_1278),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1893),
.A2(n_1355),
.B1(n_1358),
.B2(n_1350),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1785),
.Y(n_2053)
);

INVx2_ASAP7_75t_SL g2054 ( 
.A(n_1980),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1789),
.B(n_1778),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1894),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1786),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1832),
.B(n_1229),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1792),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1968),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_1815),
.B(n_1475),
.C(n_1465),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1804),
.B(n_1365),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1874),
.A2(n_1372),
.B1(n_1373),
.B2(n_1370),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1974),
.Y(n_2064)
);

INVx2_ASAP7_75t_SL g2065 ( 
.A(n_1980),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1994),
.B(n_1378),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1976),
.Y(n_2067)
);

O2A1O1Ixp33_ASAP7_75t_L g2068 ( 
.A1(n_1840),
.A2(n_1319),
.B(n_1322),
.C(n_1310),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1985),
.B(n_1383),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1787),
.A2(n_1828),
.B(n_1820),
.Y(n_2070)
);

AND2x4_ASAP7_75t_L g2071 ( 
.A(n_1967),
.B(n_1884),
.Y(n_2071)
);

OAI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_1852),
.A2(n_1289),
.B1(n_1347),
.B2(n_1269),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1813),
.B(n_1384),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1981),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1989),
.B(n_1990),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1783),
.A2(n_1472),
.B(n_1421),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1784),
.A2(n_1472),
.B(n_1421),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1814),
.B(n_1885),
.Y(n_2078)
);

BUFx6f_ASAP7_75t_L g2079 ( 
.A(n_1959),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1799),
.B(n_1469),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1839),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1909),
.B(n_1390),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1801),
.B(n_1833),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1947),
.B(n_1470),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1829),
.B(n_1001),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1848),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1850),
.Y(n_2087)
);

NOR3xp33_ASAP7_75t_L g2088 ( 
.A(n_1979),
.B(n_1040),
.C(n_1006),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1991),
.Y(n_2089)
);

O2A1O1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1868),
.A2(n_1339),
.B(n_1340),
.C(n_1327),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_L g2091 ( 
.A(n_1984),
.B(n_1388),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1959),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1959),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_SL g2094 ( 
.A(n_1897),
.B(n_1289),
.Y(n_2094)
);

INVxp67_ASAP7_75t_L g2095 ( 
.A(n_1901),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1874),
.A2(n_1393),
.B1(n_1397),
.B2(n_1391),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_1931),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1862),
.B(n_1400),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1869),
.B(n_1402),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1876),
.Y(n_2100)
);

BUFx6f_ASAP7_75t_L g2101 ( 
.A(n_1927),
.Y(n_2101)
);

OAI22xp5_ASAP7_75t_L g2102 ( 
.A1(n_1891),
.A2(n_1347),
.B1(n_1064),
.B2(n_1069),
.Y(n_2102)
);

NOR2x1p5_ASAP7_75t_L g2103 ( 
.A(n_1797),
.B(n_1405),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_1991),
.Y(n_2104)
);

INVxp67_ASAP7_75t_L g2105 ( 
.A(n_1958),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1793),
.B(n_1450),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1886),
.B(n_1410),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1896),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1903),
.Y(n_2109)
);

NOR2xp33_ASAP7_75t_L g2110 ( 
.A(n_1986),
.B(n_1414),
.Y(n_2110)
);

AND2x4_ASAP7_75t_SL g2111 ( 
.A(n_1964),
.B(n_987),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1827),
.B(n_1816),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1857),
.B(n_1418),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_L g2114 ( 
.A1(n_1970),
.A2(n_1425),
.B1(n_1428),
.B2(n_1419),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1907),
.Y(n_2115)
);

INVxp67_ASAP7_75t_L g2116 ( 
.A(n_1800),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1892),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1898),
.B(n_1444),
.Y(n_2118)
);

OR2x6_ASAP7_75t_L g2119 ( 
.A(n_1821),
.B(n_1087),
.Y(n_2119)
);

BUFx8_ASAP7_75t_L g2120 ( 
.A(n_1798),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1993),
.B(n_1436),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1794),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1856),
.B(n_1437),
.Y(n_2123)
);

NOR2xp33_ASAP7_75t_SL g2124 ( 
.A(n_1879),
.B(n_1089),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1927),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_SL g2126 ( 
.A(n_1905),
.B(n_1449),
.Y(n_2126)
);

INVx2_ASAP7_75t_SL g2127 ( 
.A(n_1977),
.Y(n_2127)
);

NOR2xp33_ASAP7_75t_L g2128 ( 
.A(n_1864),
.B(n_1826),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1849),
.B(n_1438),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1853),
.B(n_1443),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_1970),
.A2(n_1447),
.B1(n_1452),
.B2(n_1445),
.Y(n_2131)
);

NOR2xp33_ASAP7_75t_L g2132 ( 
.A(n_1864),
.B(n_1453),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1899),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_1900),
.Y(n_2134)
);

AOI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_1870),
.A2(n_1463),
.B1(n_1467),
.B2(n_1458),
.Y(n_2135)
);

NOR3xp33_ASAP7_75t_L g2136 ( 
.A(n_1935),
.B(n_1130),
.C(n_1109),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1796),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_SL g2138 ( 
.A(n_1806),
.B(n_984),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_1834),
.B(n_1424),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1875),
.Y(n_2140)
);

NAND3xp33_ASAP7_75t_SL g2141 ( 
.A(n_1803),
.B(n_1232),
.C(n_1149),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1875),
.B(n_985),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1838),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_1878),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1835),
.B(n_1349),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_1831),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_1842),
.B(n_986),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1845),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1843),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1858),
.B(n_1480),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1823),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1824),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_1809),
.B(n_994),
.Y(n_2153)
);

AND2x6_ASAP7_75t_SL g2154 ( 
.A(n_1946),
.B(n_1003),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_SL g2155 ( 
.A(n_1972),
.B(n_1205),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1912),
.B(n_1474),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_1917),
.A2(n_1353),
.B1(n_1354),
.B2(n_1351),
.Y(n_2157)
);

BUFx6f_ASAP7_75t_L g2158 ( 
.A(n_1933),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1982),
.B(n_1205),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1922),
.A2(n_1359),
.B1(n_1361),
.B2(n_1357),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1895),
.A2(n_1002),
.B1(n_1004),
.B2(n_999),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1925),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1930),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_1904),
.A2(n_1473),
.B(n_1371),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_SL g2165 ( 
.A(n_1910),
.B(n_1011),
.Y(n_2165)
);

INVxp67_ASAP7_75t_SL g2166 ( 
.A(n_1915),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1913),
.B(n_1017),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1855),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_1877),
.A2(n_1376),
.B1(n_1381),
.B2(n_1367),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1859),
.B(n_1483),
.Y(n_2170)
);

AOI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_1867),
.A2(n_1473),
.B(n_1385),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_1873),
.B(n_1882),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1916),
.B(n_1021),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1851),
.B(n_1389),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_1943),
.Y(n_2175)
);

NOR2xp67_ASAP7_75t_L g2176 ( 
.A(n_1902),
.B(n_3),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1782),
.B(n_1027),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_1811),
.B(n_1028),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1908),
.B(n_1034),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1860),
.B(n_1464),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_1949),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1861),
.B(n_1047),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1880),
.B(n_1468),
.Y(n_2183)
);

AND2x4_ASAP7_75t_SL g2184 ( 
.A(n_1996),
.B(n_1205),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1940),
.B(n_1063),
.Y(n_2185)
);

INVxp33_ASAP7_75t_L g2186 ( 
.A(n_1954),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1837),
.B(n_1070),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_1932),
.B(n_1255),
.Y(n_2188)
);

AOI22xp33_ASAP7_75t_L g2189 ( 
.A1(n_1883),
.A2(n_1396),
.B1(n_1399),
.B2(n_1394),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1937),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1937),
.Y(n_2191)
);

INVx3_ASAP7_75t_L g2192 ( 
.A(n_1841),
.Y(n_2192)
);

INVxp67_ASAP7_75t_L g2193 ( 
.A(n_1953),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1950),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_1821),
.Y(n_2195)
);

NOR2xp33_ASAP7_75t_L g2196 ( 
.A(n_1895),
.B(n_1080),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1988),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1938),
.B(n_1079),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_1995),
.B(n_1082),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1918),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_1942),
.A2(n_1404),
.B(n_1401),
.Y(n_2201)
);

BUFx3_ASAP7_75t_L g2202 ( 
.A(n_1802),
.Y(n_2202)
);

INVx2_ASAP7_75t_SL g2203 ( 
.A(n_1802),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1819),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1929),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1846),
.Y(n_2206)
);

INVx2_ASAP7_75t_SL g2207 ( 
.A(n_1817),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1960),
.B(n_1415),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_1928),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1933),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1817),
.B(n_1086),
.Y(n_2211)
);

INVx3_ASAP7_75t_L g2212 ( 
.A(n_1955),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1818),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1818),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1790),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1830),
.Y(n_2216)
);

BUFx6f_ASAP7_75t_L g2217 ( 
.A(n_1956),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_SL g2218 ( 
.A(n_1844),
.B(n_1098),
.Y(n_2218)
);

A2O1A1Ixp33_ASAP7_75t_L g2219 ( 
.A1(n_1920),
.A2(n_1423),
.B(n_1427),
.C(n_1420),
.Y(n_2219)
);

INVx3_ASAP7_75t_L g2220 ( 
.A(n_1998),
.Y(n_2220)
);

AO221x1_ASAP7_75t_L g2221 ( 
.A1(n_1934),
.A2(n_1259),
.B1(n_1333),
.B2(n_1264),
.C(n_1222),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1924),
.Y(n_2222)
);

AND2x2_ASAP7_75t_SL g2223 ( 
.A(n_1921),
.B(n_1433),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1939),
.B(n_1255),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_1941),
.B(n_1105),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_1944),
.B(n_1457),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_1945),
.B(n_1106),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1951),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1936),
.Y(n_2229)
);

NOR2xp33_ASAP7_75t_L g2230 ( 
.A(n_1948),
.B(n_1119),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_1957),
.B(n_1255),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_1966),
.B(n_1120),
.Y(n_2232)
);

OR2x6_ASAP7_75t_L g2233 ( 
.A(n_1791),
.B(n_1087),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1887),
.Y(n_2234)
);

OAI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_1961),
.A2(n_1317),
.B1(n_1430),
.B2(n_1312),
.C(n_1262),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1966),
.B(n_1121),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1887),
.Y(n_2237)
);

NAND2x1_ASAP7_75t_L g2238 ( 
.A(n_1874),
.B(n_1222),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1966),
.B(n_1140),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1780),
.B(n_1256),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1780),
.B(n_1154),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_1780),
.B(n_1155),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_1822),
.A2(n_1259),
.B1(n_1264),
.B2(n_1222),
.Y(n_2243)
);

OR2x6_ASAP7_75t_L g2244 ( 
.A(n_1791),
.B(n_1163),
.Y(n_2244)
);

NAND2xp33_ASAP7_75t_L g2245 ( 
.A(n_1874),
.B(n_1134),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1807),
.B(n_1158),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_1780),
.B(n_1165),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_1966),
.B(n_1177),
.Y(n_2248)
);

AOI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_1979),
.A2(n_1024),
.B1(n_1025),
.B2(n_1009),
.C(n_1008),
.Y(n_2249)
);

OR2x2_ASAP7_75t_L g2250 ( 
.A(n_1780),
.B(n_1439),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_1966),
.B(n_1184),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1966),
.B(n_1188),
.Y(n_2252)
);

AND2x6_ASAP7_75t_SL g2253 ( 
.A(n_1935),
.B(n_1037),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1807),
.B(n_1197),
.Y(n_2254)
);

INVx3_ASAP7_75t_L g2255 ( 
.A(n_1875),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1887),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_SL g2257 ( 
.A(n_1906),
.B(n_1256),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1887),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1966),
.B(n_1198),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_1780),
.B(n_1208),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1966),
.B(n_1214),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_1785),
.Y(n_2262)
);

OAI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_1780),
.A2(n_1057),
.B1(n_1071),
.B2(n_1041),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1887),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1887),
.Y(n_2265)
);

NOR3xp33_ASAP7_75t_L g2266 ( 
.A(n_1952),
.B(n_1220),
.C(n_1216),
.Y(n_2266)
);

AOI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_1822),
.A2(n_1264),
.B1(n_1333),
.B2(n_1259),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1887),
.Y(n_2268)
);

AOI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_1780),
.A2(n_1233),
.B1(n_1234),
.B2(n_1231),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_SL g2270 ( 
.A1(n_1970),
.A2(n_1395),
.B1(n_1256),
.B2(n_1241),
.Y(n_2270)
);

NOR2xp33_ASAP7_75t_L g2271 ( 
.A(n_1807),
.B(n_1239),
.Y(n_2271)
);

AND2x6_ASAP7_75t_L g2272 ( 
.A(n_2079),
.B(n_1264),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2070),
.A2(n_1078),
.B(n_1074),
.Y(n_2273)
);

CKINVDCx10_ASAP7_75t_R g2274 ( 
.A(n_2008),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2048),
.B(n_2028),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1999),
.B(n_1245),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_2172),
.A2(n_1092),
.B(n_1081),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2016),
.Y(n_2278)
);

AND2x4_ASAP7_75t_L g2279 ( 
.A(n_2166),
.B(n_1094),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2026),
.Y(n_2280)
);

NOR2xp33_ASAP7_75t_L g2281 ( 
.A(n_2193),
.B(n_1246),
.Y(n_2281)
);

INVx3_ASAP7_75t_L g2282 ( 
.A(n_2079),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2075),
.A2(n_1257),
.B1(n_1270),
.B2(n_1251),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2004),
.B(n_1274),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_2008),
.Y(n_2285)
);

O2A1O1Ixp5_ASAP7_75t_SL g2286 ( 
.A1(n_2215),
.A2(n_1196),
.B(n_1202),
.C(n_1201),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2039),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2105),
.B(n_1283),
.Y(n_2288)
);

OAI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2112),
.A2(n_1285),
.B1(n_1291),
.B2(n_1284),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2055),
.A2(n_1275),
.B(n_1273),
.Y(n_2290)
);

AOI21xp5_ASAP7_75t_L g2291 ( 
.A1(n_2143),
.A2(n_1290),
.B(n_1280),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2012),
.B(n_1297),
.Y(n_2292)
);

CKINVDCx5p33_ASAP7_75t_R g2293 ( 
.A(n_2120),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2246),
.B(n_1395),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2047),
.B(n_1298),
.Y(n_2295)
);

NOR2xp67_ASAP7_75t_L g2296 ( 
.A(n_2095),
.B(n_1),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2014),
.A2(n_1303),
.B1(n_1305),
.B2(n_1302),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2116),
.B(n_1314),
.Y(n_2298)
);

OAI21xp33_ASAP7_75t_L g2299 ( 
.A1(n_2271),
.A2(n_1318),
.B(n_1315),
.Y(n_2299)
);

AND2x4_ASAP7_75t_L g2300 ( 
.A(n_2042),
.B(n_1296),
.Y(n_2300)
);

AND2x4_ASAP7_75t_L g2301 ( 
.A(n_2234),
.B(n_1299),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_SL g2302 ( 
.A(n_2257),
.B(n_1344),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2254),
.B(n_1346),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2171),
.A2(n_1329),
.B(n_1326),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2186),
.B(n_2188),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2082),
.B(n_2209),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2149),
.A2(n_1337),
.B(n_1331),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2168),
.A2(n_2045),
.B(n_2170),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2237),
.B(n_1348),
.Y(n_2309)
);

OAI21xp5_ASAP7_75t_L g2310 ( 
.A1(n_2076),
.A2(n_2077),
.B(n_2133),
.Y(n_2310)
);

OAI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2164),
.A2(n_1422),
.B(n_1417),
.Y(n_2311)
);

INVx4_ASAP7_75t_L g2312 ( 
.A(n_2018),
.Y(n_2312)
);

O2A1O1Ixp33_ASAP7_75t_L g2313 ( 
.A1(n_2208),
.A2(n_1448),
.B(n_1451),
.C(n_1441),
.Y(n_2313)
);

AOI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_2010),
.A2(n_1363),
.B1(n_1368),
.B2(n_1362),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2256),
.Y(n_2315)
);

INVx4_ASAP7_75t_L g2316 ( 
.A(n_2018),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2017),
.A2(n_1374),
.B1(n_1377),
.B2(n_1369),
.Y(n_2317)
);

OAI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2134),
.A2(n_1489),
.B(n_1209),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2258),
.B(n_1398),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2264),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2197),
.B(n_1407),
.Y(n_2321)
);

NOR2xp33_ASAP7_75t_L g2322 ( 
.A(n_2084),
.B(n_1408),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2265),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2268),
.B(n_1411),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2157),
.B(n_1412),
.Y(n_2325)
);

AO32x2_ASAP7_75t_L g2326 ( 
.A1(n_2263),
.A2(n_2221),
.A3(n_2195),
.B1(n_2131),
.B2(n_2114),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2057),
.Y(n_2327)
);

NOR2xp67_ASAP7_75t_L g2328 ( 
.A(n_2146),
.B(n_1),
.Y(n_2328)
);

O2A1O1Ixp5_ASAP7_75t_L g2329 ( 
.A1(n_2200),
.A2(n_1219),
.B(n_1288),
.C(n_1235),
.Y(n_2329)
);

NOR2xp33_ASAP7_75t_L g2330 ( 
.A(n_2139),
.B(n_1416),
.Y(n_2330)
);

A2O1A1Ixp33_ASAP7_75t_L g2331 ( 
.A1(n_2046),
.A2(n_2175),
.B(n_2030),
.C(n_2090),
.Y(n_2331)
);

NOR2x1_ASAP7_75t_L g2332 ( 
.A(n_2013),
.B(n_1406),
.Y(n_2332)
);

AOI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_2011),
.A2(n_1432),
.B(n_1429),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2027),
.B(n_1434),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2040),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2049),
.A2(n_1440),
.B1(n_1446),
.B2(n_1435),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2223),
.B(n_1484),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2059),
.Y(n_2338)
);

AOI21xp5_ASAP7_75t_L g2339 ( 
.A1(n_2021),
.A2(n_1460),
.B(n_1459),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_2181),
.B(n_2033),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2081),
.Y(n_2341)
);

OR2x6_ASAP7_75t_SL g2342 ( 
.A(n_2050),
.B(n_1477),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2060),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2058),
.B(n_1395),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2101),
.B(n_1156),
.Y(n_2345)
);

AOI33xp33_ASAP7_75t_L g2346 ( 
.A1(n_2169),
.A2(n_5),
.A3(n_7),
.B1(n_3),
.B2(n_4),
.B3(n_6),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2156),
.B(n_3),
.Y(n_2347)
);

CKINVDCx10_ASAP7_75t_R g2348 ( 
.A(n_2119),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2101),
.B(n_1156),
.Y(n_2349)
);

AOI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_2094),
.A2(n_1462),
.B1(n_1392),
.B2(n_6),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2092),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_2044),
.A2(n_2083),
.B(n_2126),
.Y(n_2352)
);

NOR3xp33_ASAP7_75t_L g2353 ( 
.A(n_2141),
.B(n_6),
.C(n_5),
.Y(n_2353)
);

NOR2xp67_ASAP7_75t_L g2354 ( 
.A(n_2148),
.B(n_4),
.Y(n_2354)
);

AOI21xp5_ASAP7_75t_L g2355 ( 
.A1(n_2069),
.A2(n_1462),
.B(n_1392),
.Y(n_2355)
);

NOR2x1_ASAP7_75t_L g2356 ( 
.A(n_2013),
.B(n_1392),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2064),
.Y(n_2357)
);

AOI211xp5_ASAP7_75t_L g2358 ( 
.A1(n_2072),
.A2(n_2051),
.B(n_2204),
.C(n_2235),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2087),
.Y(n_2359)
);

BUFx12f_ASAP7_75t_L g2360 ( 
.A(n_2120),
.Y(n_2360)
);

AOI21xp5_ASAP7_75t_L g2361 ( 
.A1(n_2098),
.A2(n_8),
.B(n_9),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_2125),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2099),
.A2(n_8),
.B(n_9),
.Y(n_2363)
);

BUFx12f_ASAP7_75t_L g2364 ( 
.A(n_2097),
.Y(n_2364)
);

HB1xp67_ASAP7_75t_L g2365 ( 
.A(n_2233),
.Y(n_2365)
);

NAND3xp33_ASAP7_75t_L g2366 ( 
.A(n_2270),
.B(n_9),
.C(n_10),
.Y(n_2366)
);

INVxp67_ASAP7_75t_L g2367 ( 
.A(n_2124),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2117),
.Y(n_2368)
);

AOI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2107),
.A2(n_10),
.B(n_11),
.Y(n_2369)
);

A2O1A1Ixp33_ASAP7_75t_L g2370 ( 
.A1(n_2068),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2189),
.B(n_12),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2227),
.A2(n_13),
.B(n_14),
.Y(n_2372)
);

AOI22xp33_ASAP7_75t_L g2373 ( 
.A1(n_2061),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2108),
.Y(n_2374)
);

AO21x1_ASAP7_75t_L g2375 ( 
.A1(n_2245),
.A2(n_710),
.B(n_709),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2145),
.B(n_15),
.Y(n_2376)
);

AOI21xp5_ASAP7_75t_L g2377 ( 
.A1(n_2222),
.A2(n_16),
.B(n_17),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2102),
.B(n_2250),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2150),
.B(n_18),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2125),
.B(n_2158),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2109),
.Y(n_2381)
);

O2A1O1Ixp33_ASAP7_75t_L g2382 ( 
.A1(n_2219),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_2382)
);

OAI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2067),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_2383)
);

AOI22xp33_ASAP7_75t_L g2384 ( 
.A1(n_2088),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_2384)
);

NOR3xp33_ASAP7_75t_L g2385 ( 
.A(n_2136),
.B(n_25),
.C(n_23),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2162),
.A2(n_22),
.B(n_23),
.Y(n_2386)
);

OR2x2_ASAP7_75t_SL g2387 ( 
.A(n_2080),
.B(n_22),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2086),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2034),
.B(n_26),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_2158),
.Y(n_2390)
);

HB1xp67_ASAP7_75t_L g2391 ( 
.A(n_2233),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2163),
.A2(n_26),
.B(n_27),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2100),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2115),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2122),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2240),
.B(n_27),
.Y(n_2396)
);

AOI22xp33_ASAP7_75t_L g2397 ( 
.A1(n_2153),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2118),
.A2(n_2130),
.B(n_2129),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2036),
.B(n_31),
.Y(n_2399)
);

AOI22xp33_ASAP7_75t_L g2400 ( 
.A1(n_2249),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_2400)
);

INVx4_ASAP7_75t_L g2401 ( 
.A(n_2244),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2228),
.A2(n_32),
.B(n_33),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2052),
.B(n_33),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2056),
.Y(n_2404)
);

AOI21xp5_ASAP7_75t_L g2405 ( 
.A1(n_2229),
.A2(n_35),
.B(n_36),
.Y(n_2405)
);

AOI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2151),
.A2(n_35),
.B(n_37),
.Y(n_2406)
);

AO21x1_ASAP7_75t_L g2407 ( 
.A1(n_2019),
.A2(n_712),
.B(n_711),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2266),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2408)
);

OAI21xp5_ASAP7_75t_L g2409 ( 
.A1(n_2226),
.A2(n_37),
.B(n_38),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2152),
.A2(n_38),
.B(n_39),
.Y(n_2410)
);

BUFx6f_ASAP7_75t_L g2411 ( 
.A(n_2158),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_SL g2412 ( 
.A(n_2002),
.B(n_41),
.Y(n_2412)
);

AOI21xp5_ASAP7_75t_L g2413 ( 
.A1(n_2232),
.A2(n_40),
.B(n_41),
.Y(n_2413)
);

CKINVDCx10_ASAP7_75t_R g2414 ( 
.A(n_2119),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2236),
.A2(n_40),
.B(n_41),
.Y(n_2415)
);

INVx2_ASAP7_75t_L g2416 ( 
.A(n_2137),
.Y(n_2416)
);

BUFx8_ASAP7_75t_SL g2417 ( 
.A(n_2244),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2066),
.B(n_2085),
.Y(n_2418)
);

NOR2xp33_ASAP7_75t_L g2419 ( 
.A(n_2177),
.B(n_40),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2085),
.B(n_42),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2063),
.B(n_43),
.Y(n_2421)
);

NOR2x1_ASAP7_75t_L g2422 ( 
.A(n_2001),
.B(n_44),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2174),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2239),
.A2(n_45),
.B(n_46),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2041),
.B(n_45),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2199),
.B(n_45),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2135),
.B(n_46),
.Y(n_2427)
);

AOI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2248),
.A2(n_2261),
.B(n_2259),
.Y(n_2428)
);

BUFx6f_ASAP7_75t_L g2429 ( 
.A(n_2093),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2031),
.B(n_47),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2180),
.Y(n_2431)
);

BUFx3_ASAP7_75t_L g2432 ( 
.A(n_2202),
.Y(n_2432)
);

AOI22x1_ASAP7_75t_L g2433 ( 
.A1(n_2201),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2113),
.B(n_49),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2160),
.B(n_50),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2000),
.B(n_52),
.Y(n_2436)
);

AOI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2251),
.A2(n_53),
.B(n_54),
.Y(n_2437)
);

AND2x6_ASAP7_75t_SL g2438 ( 
.A(n_2007),
.B(n_53),
.Y(n_2438)
);

AOI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2252),
.A2(n_54),
.B(n_55),
.Y(n_2439)
);

BUFx3_ASAP7_75t_L g2440 ( 
.A(n_2214),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2015),
.B(n_56),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2096),
.B(n_57),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2009),
.B(n_57),
.Y(n_2443)
);

NOR2xp33_ASAP7_75t_L g2444 ( 
.A(n_2006),
.B(n_58),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2140),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2183),
.B(n_59),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2269),
.B(n_61),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_2111),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2003),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_2449)
);

A2O1A1Ixp33_ASAP7_75t_L g2450 ( 
.A1(n_2023),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_2450)
);

AOI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2179),
.A2(n_63),
.B(n_64),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2231),
.B(n_64),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2155),
.B(n_66),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2073),
.B(n_67),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2194),
.Y(n_2455)
);

INVxp67_ASAP7_75t_L g2456 ( 
.A(n_2015),
.Y(n_2456)
);

OR2x2_ASAP7_75t_L g2457 ( 
.A(n_2104),
.B(n_68),
.Y(n_2457)
);

AOI21xp5_ASAP7_75t_L g2458 ( 
.A1(n_2078),
.A2(n_69),
.B(n_70),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2138),
.A2(n_69),
.B(n_70),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_SL g2460 ( 
.A(n_2093),
.B(n_72),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_SL g2461 ( 
.A(n_2161),
.B(n_72),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2091),
.B(n_2110),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_SL g2463 ( 
.A(n_2123),
.B(n_74),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2210),
.Y(n_2464)
);

OAI22xp5_ASAP7_75t_L g2465 ( 
.A1(n_2243),
.A2(n_2267),
.B1(n_2255),
.B2(n_2144),
.Y(n_2465)
);

OAI22xp5_ASAP7_75t_L g2466 ( 
.A1(n_2144),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2217),
.Y(n_2467)
);

BUFx8_ASAP7_75t_SL g2468 ( 
.A(n_2220),
.Y(n_2468)
);

OAI22xp5_ASAP7_75t_L g2469 ( 
.A1(n_2255),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_2165),
.A2(n_76),
.B(n_77),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2121),
.B(n_77),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2159),
.B(n_77),
.Y(n_2472)
);

BUFx4f_ASAP7_75t_L g2473 ( 
.A(n_2220),
.Y(n_2473)
);

A2O1A1Ixp33_ASAP7_75t_L g2474 ( 
.A1(n_2230),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_2474)
);

O2A1O1Ixp33_ASAP7_75t_L g2475 ( 
.A1(n_2185),
.A2(n_82),
.B(n_78),
.C(n_81),
.Y(n_2475)
);

AOI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_2167),
.A2(n_81),
.B(n_82),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2173),
.A2(n_81),
.B(n_82),
.Y(n_2477)
);

AOI21xp5_ASAP7_75t_L g2478 ( 
.A1(n_2225),
.A2(n_83),
.B(n_84),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2132),
.B(n_83),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_2190),
.Y(n_2480)
);

OAI22xp5_ASAP7_75t_L g2481 ( 
.A1(n_2062),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2103),
.B(n_84),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2224),
.B(n_85),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2196),
.B(n_86),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2217),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2241),
.B(n_86),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2242),
.B(n_88),
.Y(n_2487)
);

INVx11_ASAP7_75t_L g2488 ( 
.A(n_2029),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2198),
.A2(n_88),
.B(n_89),
.Y(n_2489)
);

NOR2xp33_ASAP7_75t_L g2490 ( 
.A(n_2247),
.B(n_89),
.Y(n_2490)
);

OAI21xp5_ASAP7_75t_L g2491 ( 
.A1(n_2147),
.A2(n_90),
.B(n_91),
.Y(n_2491)
);

NAND2x1_ASAP7_75t_L g2492 ( 
.A(n_2212),
.B(n_91),
.Y(n_2492)
);

AOI21xp5_ASAP7_75t_L g2493 ( 
.A1(n_2128),
.A2(n_92),
.B(n_93),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_2260),
.B(n_94),
.Y(n_2494)
);

NAND2x1p5_ASAP7_75t_L g2495 ( 
.A(n_2053),
.B(n_95),
.Y(n_2495)
);

AO21x1_ASAP7_75t_L g2496 ( 
.A1(n_2024),
.A2(n_715),
.B(n_714),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2106),
.B(n_96),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2071),
.B(n_96),
.Y(n_2498)
);

AO21x1_ASAP7_75t_L g2499 ( 
.A1(n_2024),
.A2(n_2035),
.B(n_2142),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2035),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2071),
.B(n_2020),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_2074),
.Y(n_2502)
);

OAI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2178),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2022),
.B(n_100),
.Y(n_2504)
);

O2A1O1Ixp33_ASAP7_75t_L g2505 ( 
.A1(n_2182),
.A2(n_103),
.B(n_101),
.C(n_102),
.Y(n_2505)
);

O2A1O1Ixp33_ASAP7_75t_L g2506 ( 
.A1(n_2211),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_2506)
);

O2A1O1Ixp33_ASAP7_75t_L g2507 ( 
.A1(n_2218),
.A2(n_105),
.B(n_102),
.C(n_103),
.Y(n_2507)
);

INVx2_ASAP7_75t_SL g2508 ( 
.A(n_2262),
.Y(n_2508)
);

OAI21x1_ASAP7_75t_L g2509 ( 
.A1(n_2191),
.A2(n_718),
.B(n_717),
.Y(n_2509)
);

OR2x2_ASAP7_75t_SL g2510 ( 
.A(n_2154),
.B(n_106),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2037),
.B(n_109),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2038),
.B(n_2054),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2212),
.Y(n_2513)
);

OAI21xp5_ASAP7_75t_L g2514 ( 
.A1(n_2025),
.A2(n_2187),
.B(n_2205),
.Y(n_2514)
);

NOR2xp33_ASAP7_75t_R g2515 ( 
.A(n_2203),
.B(n_110),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2065),
.B(n_111),
.Y(n_2516)
);

INVx3_ASAP7_75t_L g2517 ( 
.A(n_2192),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2089),
.B(n_116),
.Y(n_2518)
);

NAND2x1_ASAP7_75t_L g2519 ( 
.A(n_2192),
.B(n_114),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2206),
.Y(n_2520)
);

OAI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_2213),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2521)
);

OAI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_2216),
.A2(n_118),
.B(n_119),
.Y(n_2522)
);

BUFx3_ASAP7_75t_L g2523 ( 
.A(n_2207),
.Y(n_2523)
);

AOI21xp5_ASAP7_75t_L g2524 ( 
.A1(n_2127),
.A2(n_2184),
.B(n_2043),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2253),
.B(n_120),
.Y(n_2525)
);

OAI22xp5_ASAP7_75t_L g2526 ( 
.A1(n_2048),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2048),
.B(n_120),
.Y(n_2527)
);

AOI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2048),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2048),
.B(n_122),
.Y(n_2529)
);

BUFx6f_ASAP7_75t_L g2530 ( 
.A(n_2101),
.Y(n_2530)
);

INVx4_ASAP7_75t_L g2531 ( 
.A(n_2018),
.Y(n_2531)
);

AOI21xp5_ASAP7_75t_L g2532 ( 
.A1(n_2070),
.A2(n_123),
.B(n_124),
.Y(n_2532)
);

A2O1A1Ixp33_ASAP7_75t_L g2533 ( 
.A1(n_2112),
.A2(n_127),
.B(n_125),
.C(n_126),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2048),
.B(n_125),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2048),
.B(n_125),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2048),
.B(n_126),
.Y(n_2536)
);

AOI21xp5_ASAP7_75t_L g2537 ( 
.A1(n_2070),
.A2(n_128),
.B(n_129),
.Y(n_2537)
);

HB1xp67_ASAP7_75t_L g2538 ( 
.A(n_2012),
.Y(n_2538)
);

NAND3xp33_ASAP7_75t_L g2539 ( 
.A(n_2270),
.B(n_129),
.C(n_131),
.Y(n_2539)
);

AOI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2070),
.A2(n_131),
.B(n_132),
.Y(n_2540)
);

OAI21xp33_ASAP7_75t_L g2541 ( 
.A1(n_1999),
.A2(n_132),
.B(n_133),
.Y(n_2541)
);

INVx2_ASAP7_75t_SL g2542 ( 
.A(n_2120),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2016),
.Y(n_2543)
);

INVxp67_ASAP7_75t_L g2544 ( 
.A(n_2012),
.Y(n_2544)
);

NOR2x1_ASAP7_75t_L g2545 ( 
.A(n_2013),
.B(n_132),
.Y(n_2545)
);

AOI21xp5_ASAP7_75t_L g2546 ( 
.A1(n_2070),
.A2(n_133),
.B(n_134),
.Y(n_2546)
);

O2A1O1Ixp33_ASAP7_75t_L g2547 ( 
.A1(n_2112),
.A2(n_136),
.B(n_134),
.C(n_135),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2048),
.B(n_134),
.Y(n_2548)
);

AOI22xp5_ASAP7_75t_L g2549 ( 
.A1(n_2048),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2048),
.B(n_136),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2048),
.B(n_138),
.Y(n_2551)
);

AOI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2048),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2048),
.B(n_139),
.Y(n_2553)
);

BUFx4f_ASAP7_75t_L g2554 ( 
.A(n_2013),
.Y(n_2554)
);

INVx2_ASAP7_75t_SL g2555 ( 
.A(n_2120),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2070),
.A2(n_141),
.B(n_142),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2016),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2070),
.A2(n_141),
.B(n_142),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2016),
.Y(n_2559)
);

AOI21xp5_ASAP7_75t_L g2560 ( 
.A1(n_2070),
.A2(n_143),
.B(n_144),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2048),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_L g2562 ( 
.A(n_2193),
.B(n_143),
.Y(n_2562)
);

O2A1O1Ixp5_ASAP7_75t_L g2563 ( 
.A1(n_2032),
.A2(n_146),
.B(n_144),
.C(n_145),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2048),
.B(n_146),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_SL g2565 ( 
.A(n_2012),
.B(n_148),
.Y(n_2565)
);

NOR2xp67_ASAP7_75t_L g2566 ( 
.A(n_2095),
.B(n_147),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_2101),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2016),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2016),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2070),
.A2(n_149),
.B(n_150),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2048),
.B(n_149),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2048),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_2572)
);

AOI21xp5_ASAP7_75t_L g2573 ( 
.A1(n_2070),
.A2(n_150),
.B(n_151),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2101),
.Y(n_2574)
);

NAND2xp33_ASAP7_75t_L g2575 ( 
.A(n_2101),
.B(n_152),
.Y(n_2575)
);

OAI321xp33_ASAP7_75t_L g2576 ( 
.A1(n_2114),
.A2(n_153),
.A3(n_156),
.B1(n_151),
.B2(n_152),
.C(n_154),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2101),
.Y(n_2577)
);

AOI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_2048),
.A2(n_154),
.B1(n_152),
.B2(n_153),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2070),
.A2(n_153),
.B(n_154),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2193),
.B(n_157),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2048),
.B(n_157),
.Y(n_2581)
);

AOI21xp5_ASAP7_75t_L g2582 ( 
.A1(n_2070),
.A2(n_158),
.B(n_159),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2193),
.B(n_158),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2048),
.B(n_158),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2120),
.Y(n_2585)
);

HB1xp67_ASAP7_75t_L g2586 ( 
.A(n_2012),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2193),
.B(n_159),
.Y(n_2587)
);

NAND3xp33_ASAP7_75t_L g2588 ( 
.A(n_2270),
.B(n_160),
.C(n_161),
.Y(n_2588)
);

OAI22xp5_ASAP7_75t_L g2589 ( 
.A1(n_2048),
.A2(n_163),
.B1(n_161),
.B2(n_162),
.Y(n_2589)
);

OR2x2_ASAP7_75t_L g2590 ( 
.A(n_2050),
.B(n_162),
.Y(n_2590)
);

OAI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2048),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_2591)
);

NAND3xp33_ASAP7_75t_L g2592 ( 
.A(n_2270),
.B(n_164),
.C(n_165),
.Y(n_2592)
);

NOR2xp33_ASAP7_75t_L g2593 ( 
.A(n_2193),
.B(n_166),
.Y(n_2593)
);

CKINVDCx6p67_ASAP7_75t_R g2594 ( 
.A(n_2008),
.Y(n_2594)
);

AOI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2048),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2048),
.B(n_167),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2070),
.A2(n_168),
.B(n_169),
.Y(n_2597)
);

AOI21xp5_ASAP7_75t_L g2598 ( 
.A1(n_2070),
.A2(n_169),
.B(n_170),
.Y(n_2598)
);

A2O1A1Ixp33_ASAP7_75t_L g2599 ( 
.A1(n_2112),
.A2(n_172),
.B(n_170),
.C(n_171),
.Y(n_2599)
);

AO32x1_ASAP7_75t_L g2600 ( 
.A1(n_2221),
.A2(n_172),
.A3(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_2600)
);

AO32x1_ASAP7_75t_L g2601 ( 
.A1(n_2221),
.A2(n_173),
.A3(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2048),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2005),
.Y(n_2603)
);

AOI21xp5_ASAP7_75t_L g2604 ( 
.A1(n_2070),
.A2(n_175),
.B(n_177),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2016),
.Y(n_2605)
);

AOI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_2070),
.A2(n_178),
.B(n_179),
.Y(n_2606)
);

A2O1A1Ixp33_ASAP7_75t_L g2607 ( 
.A1(n_2112),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_2607)
);

O2A1O1Ixp33_ASAP7_75t_SL g2608 ( 
.A1(n_2238),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2070),
.A2(n_182),
.B(n_183),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2193),
.B(n_184),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2005),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2048),
.B(n_185),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2048),
.B(n_185),
.Y(n_2613)
);

A2O1A1Ixp33_ASAP7_75t_L g2614 ( 
.A1(n_2112),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_2614)
);

A2O1A1Ixp33_ASAP7_75t_L g2615 ( 
.A1(n_2112),
.A2(n_190),
.B(n_186),
.C(n_189),
.Y(n_2615)
);

INVx2_ASAP7_75t_L g2616 ( 
.A(n_2005),
.Y(n_2616)
);

AOI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2070),
.A2(n_189),
.B(n_190),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_2120),
.Y(n_2618)
);

AOI21xp5_ASAP7_75t_L g2619 ( 
.A1(n_2070),
.A2(n_189),
.B(n_190),
.Y(n_2619)
);

BUFx6f_ASAP7_75t_L g2620 ( 
.A(n_2101),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2048),
.B(n_191),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_2012),
.Y(n_2622)
);

OAI321xp33_ASAP7_75t_L g2623 ( 
.A1(n_2114),
.A2(n_194),
.A3(n_196),
.B1(n_191),
.B2(n_193),
.C(n_195),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2048),
.A2(n_196),
.B1(n_194),
.B2(n_195),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2016),
.Y(n_2625)
);

HB1xp67_ASAP7_75t_L g2626 ( 
.A(n_2012),
.Y(n_2626)
);

O2A1O1Ixp5_ASAP7_75t_L g2627 ( 
.A1(n_2032),
.A2(n_197),
.B(n_195),
.C(n_196),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2048),
.B(n_197),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2016),
.Y(n_2629)
);

OAI21x1_ASAP7_75t_L g2630 ( 
.A1(n_2005),
.A2(n_720),
.B(n_719),
.Y(n_2630)
);

OR2x6_ASAP7_75t_L g2631 ( 
.A(n_2013),
.B(n_198),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2048),
.B(n_199),
.Y(n_2632)
);

AND2x6_ASAP7_75t_SL g2633 ( 
.A(n_2119),
.B(n_200),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2048),
.B(n_201),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2048),
.B(n_201),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2048),
.A2(n_204),
.B1(n_202),
.B2(n_203),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2048),
.B(n_202),
.Y(n_2637)
);

AOI21xp5_ASAP7_75t_L g2638 ( 
.A1(n_2070),
.A2(n_204),
.B(n_205),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2016),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2048),
.B(n_205),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2193),
.B(n_205),
.Y(n_2641)
);

AND2x4_ASAP7_75t_L g2642 ( 
.A(n_2166),
.B(n_206),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_2193),
.B(n_206),
.Y(n_2643)
);

AOI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2048),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2048),
.B(n_207),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2008),
.Y(n_2646)
);

OAI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2048),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2647)
);

OAI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2048),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2016),
.Y(n_2649)
);

AOI21xp5_ASAP7_75t_L g2650 ( 
.A1(n_2070),
.A2(n_211),
.B(n_212),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2048),
.B(n_212),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2048),
.B(n_213),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2048),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2048),
.B(n_214),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2008),
.Y(n_2655)
);

AOI21xp5_ASAP7_75t_L g2656 ( 
.A1(n_2070),
.A2(n_215),
.B(n_216),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2193),
.B(n_216),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_SL g2658 ( 
.A(n_2012),
.B(n_218),
.Y(n_2658)
);

O2A1O1Ixp33_ASAP7_75t_L g2659 ( 
.A1(n_2112),
.A2(n_220),
.B(n_217),
.C(n_219),
.Y(n_2659)
);

AOI21xp5_ASAP7_75t_L g2660 ( 
.A1(n_2070),
.A2(n_217),
.B(n_220),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2048),
.B(n_221),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_SL g2662 ( 
.A(n_2012),
.B(n_222),
.Y(n_2662)
);

OAI22xp5_ASAP7_75t_L g2663 ( 
.A1(n_2048),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.Y(n_2663)
);

AO32x1_ASAP7_75t_L g2664 ( 
.A1(n_2221),
.A2(n_225),
.A3(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_2664)
);

OAI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2048),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2070),
.A2(n_227),
.B(n_228),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2193),
.B(n_229),
.Y(n_2667)
);

HB1xp67_ASAP7_75t_L g2668 ( 
.A(n_2012),
.Y(n_2668)
);

AOI21xp5_ASAP7_75t_L g2669 ( 
.A1(n_2070),
.A2(n_230),
.B(n_231),
.Y(n_2669)
);

AOI21x1_ASAP7_75t_L g2670 ( 
.A1(n_2176),
.A2(n_230),
.B(n_232),
.Y(n_2670)
);

AOI21xp5_ASAP7_75t_L g2671 ( 
.A1(n_2070),
.A2(n_232),
.B(n_233),
.Y(n_2671)
);

BUFx6f_ASAP7_75t_L g2672 ( 
.A(n_2101),
.Y(n_2672)
);

BUFx6f_ASAP7_75t_L g2673 ( 
.A(n_2101),
.Y(n_2673)
);

NOR2x1_ASAP7_75t_L g2674 ( 
.A(n_2013),
.B(n_233),
.Y(n_2674)
);

OAI22xp5_ASAP7_75t_L g2675 ( 
.A1(n_2048),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_2675)
);

AND2x2_ASAP7_75t_L g2676 ( 
.A(n_2048),
.B(n_236),
.Y(n_2676)
);

INVx1_ASAP7_75t_SL g2677 ( 
.A(n_2012),
.Y(n_2677)
);

AOI21xp5_ASAP7_75t_L g2678 ( 
.A1(n_2070),
.A2(n_238),
.B(n_239),
.Y(n_2678)
);

A2O1A1Ixp33_ASAP7_75t_L g2679 ( 
.A1(n_2112),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2679)
);

AOI21x1_ASAP7_75t_L g2680 ( 
.A1(n_2176),
.A2(n_240),
.B(n_241),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2016),
.Y(n_2681)
);

BUFx3_ASAP7_75t_L g2682 ( 
.A(n_2120),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2048),
.B(n_240),
.Y(n_2683)
);

NOR2xp67_ASAP7_75t_L g2684 ( 
.A(n_2095),
.B(n_241),
.Y(n_2684)
);

NAND3xp33_ASAP7_75t_L g2685 ( 
.A(n_2270),
.B(n_242),
.C(n_243),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_SL g2686 ( 
.A(n_2012),
.B(n_246),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2048),
.B(n_245),
.Y(n_2687)
);

NAND2xp5_ASAP7_75t_SL g2688 ( 
.A(n_2012),
.B(n_247),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2016),
.Y(n_2689)
);

A2O1A1Ixp33_ASAP7_75t_L g2690 ( 
.A1(n_2112),
.A2(n_251),
.B(n_248),
.C(n_250),
.Y(n_2690)
);

AOI21xp5_ASAP7_75t_L g2691 ( 
.A1(n_2070),
.A2(n_248),
.B(n_250),
.Y(n_2691)
);

OR2x2_ASAP7_75t_L g2692 ( 
.A(n_2050),
.B(n_250),
.Y(n_2692)
);

AOI21xp5_ASAP7_75t_L g2693 ( 
.A1(n_2070),
.A2(n_251),
.B(n_252),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2012),
.B(n_254),
.Y(n_2694)
);

AOI21x1_ASAP7_75t_L g2695 ( 
.A1(n_2176),
.A2(n_253),
.B(n_254),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2048),
.B(n_255),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2012),
.B(n_256),
.Y(n_2697)
);

AOI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2048),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_2698)
);

AOI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2070),
.A2(n_257),
.B(n_258),
.Y(n_2699)
);

OAI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2048),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_SL g2701 ( 
.A(n_2012),
.B(n_260),
.Y(n_2701)
);

A2O1A1Ixp33_ASAP7_75t_L g2702 ( 
.A1(n_2112),
.A2(n_261),
.B(n_258),
.C(n_260),
.Y(n_2702)
);

NOR2xp67_ASAP7_75t_L g2703 ( 
.A(n_2095),
.B(n_261),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2048),
.B(n_261),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2048),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2012),
.B(n_265),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2048),
.B(n_264),
.Y(n_2707)
);

OAI22xp5_ASAP7_75t_L g2708 ( 
.A1(n_2048),
.A2(n_267),
.B1(n_265),
.B2(n_266),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2012),
.B(n_268),
.Y(n_2709)
);

INVx1_ASAP7_75t_SL g2710 ( 
.A(n_2012),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2016),
.Y(n_2711)
);

BUFx2_ASAP7_75t_L g2712 ( 
.A(n_2012),
.Y(n_2712)
);

AOI21xp5_ASAP7_75t_L g2713 ( 
.A1(n_2070),
.A2(n_268),
.B(n_269),
.Y(n_2713)
);

INVx4_ASAP7_75t_L g2714 ( 
.A(n_2018),
.Y(n_2714)
);

AO32x1_ASAP7_75t_L g2715 ( 
.A1(n_2221),
.A2(n_271),
.A3(n_269),
.B1(n_270),
.B2(n_272),
.Y(n_2715)
);

AOI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2048),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_2716)
);

AOI21xp5_ASAP7_75t_L g2717 ( 
.A1(n_2070),
.A2(n_270),
.B(n_271),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2016),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2012),
.Y(n_2719)
);

AOI22xp5_ASAP7_75t_L g2720 ( 
.A1(n_2048),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2720)
);

INVx3_ASAP7_75t_SL g2721 ( 
.A(n_2013),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2048),
.B(n_275),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2048),
.B(n_275),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2048),
.B(n_276),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2048),
.B(n_276),
.Y(n_2725)
);

INVxp67_ASAP7_75t_SL g2726 ( 
.A(n_2050),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_2048),
.B(n_277),
.Y(n_2727)
);

OAI22xp5_ASAP7_75t_L g2728 ( 
.A1(n_2048),
.A2(n_279),
.B1(n_277),
.B2(n_278),
.Y(n_2728)
);

O2A1O1Ixp33_ASAP7_75t_L g2729 ( 
.A1(n_2112),
.A2(n_280),
.B(n_278),
.C(n_279),
.Y(n_2729)
);

AOI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2070),
.A2(n_282),
.B(n_283),
.Y(n_2730)
);

O2A1O1Ixp33_ASAP7_75t_L g2731 ( 
.A1(n_2112),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2016),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2101),
.Y(n_2733)
);

AOI21xp5_ASAP7_75t_L g2734 ( 
.A1(n_2070),
.A2(n_284),
.B(n_285),
.Y(n_2734)
);

NAND2x1p5_ASAP7_75t_L g2735 ( 
.A(n_2018),
.B(n_286),
.Y(n_2735)
);

O2A1O1Ixp33_ASAP7_75t_L g2736 ( 
.A1(n_2112),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_2736)
);

INVx4_ASAP7_75t_L g2737 ( 
.A(n_2018),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2048),
.B(n_287),
.Y(n_2738)
);

A2O1A1Ixp33_ASAP7_75t_L g2739 ( 
.A1(n_2112),
.A2(n_289),
.B(n_287),
.C(n_288),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_SL g2740 ( 
.A(n_2012),
.B(n_289),
.Y(n_2740)
);

AOI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2308),
.A2(n_288),
.B(n_289),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2341),
.Y(n_2742)
);

INVx4_ASAP7_75t_L g2743 ( 
.A(n_2360),
.Y(n_2743)
);

A2O1A1Ixp33_ASAP7_75t_L g2744 ( 
.A1(n_2428),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_2744)
);

OR2x2_ASAP7_75t_L g2745 ( 
.A(n_2677),
.B(n_290),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2275),
.B(n_291),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2710),
.B(n_292),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2538),
.B(n_2586),
.Y(n_2748)
);

NOR2x1_ASAP7_75t_L g2749 ( 
.A(n_2682),
.B(n_292),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2359),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_2274),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2726),
.B(n_293),
.Y(n_2752)
);

AOI21xp5_ASAP7_75t_L g2753 ( 
.A1(n_2398),
.A2(n_295),
.B(n_296),
.Y(n_2753)
);

OAI22xp5_ASAP7_75t_L g2754 ( 
.A1(n_2631),
.A2(n_2378),
.B1(n_2342),
.B2(n_2552),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2423),
.B(n_296),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_SL g2756 ( 
.A(n_2293),
.B(n_297),
.Y(n_2756)
);

AOI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2310),
.A2(n_297),
.B(n_298),
.Y(n_2757)
);

OAI21x1_ASAP7_75t_L g2758 ( 
.A1(n_2380),
.A2(n_299),
.B(n_300),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2431),
.B(n_299),
.Y(n_2759)
);

INVx5_ASAP7_75t_L g2760 ( 
.A(n_2631),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2622),
.B(n_301),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2626),
.B(n_301),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_2352),
.A2(n_302),
.B(n_303),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_SL g2764 ( 
.A(n_2554),
.B(n_720),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2278),
.Y(n_2765)
);

HB1xp67_ASAP7_75t_L g2766 ( 
.A(n_2631),
.Y(n_2766)
);

OAI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_2552),
.A2(n_305),
.B1(n_302),
.B2(n_304),
.Y(n_2767)
);

INVxp67_ASAP7_75t_L g2768 ( 
.A(n_2712),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2368),
.Y(n_2769)
);

OAI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2331),
.A2(n_304),
.B(n_305),
.Y(n_2770)
);

NAND3x1_ASAP7_75t_L g2771 ( 
.A(n_2545),
.B(n_305),
.C(n_306),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2280),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_SL g2773 ( 
.A1(n_2362),
.A2(n_307),
.B(n_308),
.Y(n_2773)
);

NAND3xp33_ASAP7_75t_L g2774 ( 
.A(n_2286),
.B(n_309),
.C(n_310),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2340),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2362),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2305),
.B(n_312),
.Y(n_2777)
);

OAI21xp5_ASAP7_75t_L g2778 ( 
.A1(n_2329),
.A2(n_313),
.B(n_315),
.Y(n_2778)
);

AOI21xp5_ASAP7_75t_L g2779 ( 
.A1(n_2355),
.A2(n_313),
.B(n_315),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2273),
.A2(n_316),
.B(n_317),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2668),
.B(n_317),
.Y(n_2781)
);

AOI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2529),
.A2(n_318),
.B(n_319),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2362),
.Y(n_2783)
);

OAI21x1_ASAP7_75t_L g2784 ( 
.A1(n_2630),
.A2(n_319),
.B(n_320),
.Y(n_2784)
);

AOI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2322),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_2785)
);

BUFx6f_ASAP7_75t_L g2786 ( 
.A(n_2390),
.Y(n_2786)
);

NOR2xp33_ASAP7_75t_SL g2787 ( 
.A(n_2554),
.B(n_321),
.Y(n_2787)
);

AND2x4_ASAP7_75t_L g2788 ( 
.A(n_2287),
.B(n_322),
.Y(n_2788)
);

AND2x4_ASAP7_75t_L g2789 ( 
.A(n_2315),
.B(n_322),
.Y(n_2789)
);

AOI21x1_ASAP7_75t_L g2790 ( 
.A1(n_2670),
.A2(n_323),
.B(n_324),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2535),
.A2(n_323),
.B(n_324),
.Y(n_2791)
);

AOI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2536),
.A2(n_324),
.B(n_325),
.Y(n_2792)
);

O2A1O1Ixp33_ASAP7_75t_SL g2793 ( 
.A1(n_2492),
.A2(n_327),
.B(n_325),
.C(n_326),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2548),
.A2(n_326),
.B(n_328),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2719),
.B(n_328),
.Y(n_2795)
);

AOI21x1_ASAP7_75t_L g2796 ( 
.A1(n_2680),
.A2(n_328),
.B(n_329),
.Y(n_2796)
);

NOR2xp33_ASAP7_75t_SL g2797 ( 
.A(n_2417),
.B(n_329),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2527),
.B(n_2534),
.Y(n_2798)
);

AND2x4_ASAP7_75t_L g2799 ( 
.A(n_2320),
.B(n_329),
.Y(n_2799)
);

OAI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2277),
.A2(n_330),
.B(n_331),
.Y(n_2800)
);

OAI21xp5_ASAP7_75t_L g2801 ( 
.A1(n_2291),
.A2(n_330),
.B(n_331),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2581),
.B(n_331),
.Y(n_2802)
);

AOI21xp5_ASAP7_75t_L g2803 ( 
.A1(n_2550),
.A2(n_332),
.B(n_333),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2323),
.Y(n_2804)
);

AOI21x1_ASAP7_75t_L g2805 ( 
.A1(n_2695),
.A2(n_334),
.B(n_335),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2551),
.A2(n_336),
.B(n_337),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2543),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2557),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_2634),
.B(n_337),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2559),
.Y(n_2810)
);

OR2x6_ASAP7_75t_L g2811 ( 
.A(n_2542),
.B(n_2555),
.Y(n_2811)
);

OAI21x1_ASAP7_75t_L g2812 ( 
.A1(n_2509),
.A2(n_338),
.B(n_339),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2568),
.Y(n_2813)
);

AOI221xp5_ASAP7_75t_L g2814 ( 
.A1(n_2313),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.C(n_341),
.Y(n_2814)
);

AOI21xp33_ASAP7_75t_L g2815 ( 
.A1(n_2553),
.A2(n_338),
.B(n_339),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2569),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_L g2817 ( 
.A(n_2637),
.B(n_340),
.Y(n_2817)
);

A2O1A1Ixp33_ASAP7_75t_L g2818 ( 
.A1(n_2541),
.A2(n_343),
.B(n_341),
.C(n_342),
.Y(n_2818)
);

AOI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2564),
.A2(n_344),
.B(n_345),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2401),
.B(n_721),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2544),
.B(n_344),
.Y(n_2821)
);

OR2x2_ASAP7_75t_L g2822 ( 
.A(n_2721),
.B(n_346),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2651),
.B(n_346),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2605),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2571),
.A2(n_347),
.B(n_348),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2661),
.B(n_348),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2676),
.B(n_349),
.Y(n_2827)
);

OAI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2561),
.A2(n_2636),
.B1(n_2716),
.B2(n_2698),
.Y(n_2828)
);

NAND2x1p5_ASAP7_75t_L g2829 ( 
.A(n_2312),
.B(n_350),
.Y(n_2829)
);

BUFx2_ASAP7_75t_L g2830 ( 
.A(n_2335),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2683),
.B(n_351),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_2707),
.B(n_351),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2625),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2723),
.B(n_351),
.Y(n_2834)
);

A2O1A1Ixp33_ASAP7_75t_L g2835 ( 
.A1(n_2491),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_2835)
);

NOR2xp33_ASAP7_75t_L g2836 ( 
.A(n_2462),
.B(n_352),
.Y(n_2836)
);

BUFx6f_ASAP7_75t_L g2837 ( 
.A(n_2390),
.Y(n_2837)
);

OR2x6_ASAP7_75t_L g2838 ( 
.A(n_2585),
.B(n_353),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2629),
.B(n_2639),
.Y(n_2839)
);

AOI21xp5_ASAP7_75t_SL g2840 ( 
.A1(n_2390),
.A2(n_355),
.B(n_356),
.Y(n_2840)
);

AO21x1_ASAP7_75t_L g2841 ( 
.A1(n_2547),
.A2(n_723),
.B(n_722),
.Y(n_2841)
);

NOR2xp33_ASAP7_75t_L g2842 ( 
.A(n_2337),
.B(n_355),
.Y(n_2842)
);

NOR2xp33_ASAP7_75t_SL g2843 ( 
.A(n_2401),
.B(n_355),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2411),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2649),
.Y(n_2845)
);

OAI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2307),
.A2(n_356),
.B(n_357),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2681),
.Y(n_2847)
);

AOI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2330),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2274),
.Y(n_2849)
);

OAI22xp5_ASAP7_75t_L g2850 ( 
.A1(n_2561),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2689),
.B(n_2711),
.Y(n_2851)
);

NOR2x1_ASAP7_75t_L g2852 ( 
.A(n_2312),
.B(n_359),
.Y(n_2852)
);

NOR2xp33_ASAP7_75t_L g2853 ( 
.A(n_2456),
.B(n_359),
.Y(n_2853)
);

OAI21x1_ASAP7_75t_L g2854 ( 
.A1(n_2345),
.A2(n_360),
.B(n_361),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2718),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2732),
.B(n_360),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2358),
.B(n_361),
.Y(n_2857)
);

AND2x4_ASAP7_75t_L g2858 ( 
.A(n_2356),
.B(n_361),
.Y(n_2858)
);

AOI21xp5_ASAP7_75t_L g2859 ( 
.A1(n_2584),
.A2(n_362),
.B(n_363),
.Y(n_2859)
);

INVx4_ASAP7_75t_L g2860 ( 
.A(n_2594),
.Y(n_2860)
);

OAI21xp5_ASAP7_75t_L g2861 ( 
.A1(n_2563),
.A2(n_362),
.B(n_363),
.Y(n_2861)
);

NAND2x1p5_ASAP7_75t_L g2862 ( 
.A(n_2316),
.B(n_364),
.Y(n_2862)
);

OAI21x1_ASAP7_75t_L g2863 ( 
.A1(n_2349),
.A2(n_365),
.B(n_366),
.Y(n_2863)
);

BUFx3_ASAP7_75t_L g2864 ( 
.A(n_2618),
.Y(n_2864)
);

BUFx2_ASAP7_75t_SL g2865 ( 
.A(n_2316),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2418),
.B(n_365),
.Y(n_2866)
);

AND2x2_ASAP7_75t_L g2867 ( 
.A(n_2525),
.B(n_367),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2327),
.Y(n_2868)
);

NOR2x1_ASAP7_75t_SL g2869 ( 
.A(n_2411),
.B(n_367),
.Y(n_2869)
);

CKINVDCx5p33_ASAP7_75t_R g2870 ( 
.A(n_2348),
.Y(n_2870)
);

AOI21xp5_ASAP7_75t_L g2871 ( 
.A1(n_2596),
.A2(n_367),
.B(n_368),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2435),
.B(n_368),
.Y(n_2872)
);

BUFx4f_ASAP7_75t_L g2873 ( 
.A(n_2364),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2612),
.A2(n_369),
.B(n_370),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2338),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2441),
.B(n_369),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2343),
.B(n_370),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2357),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2613),
.A2(n_370),
.B(n_371),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2388),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2395),
.Y(n_2881)
);

INVx3_ASAP7_75t_L g2882 ( 
.A(n_2411),
.Y(n_2882)
);

BUFx6f_ASAP7_75t_L g2883 ( 
.A(n_2530),
.Y(n_2883)
);

AO31x2_ASAP7_75t_L g2884 ( 
.A1(n_2375),
.A2(n_373),
.A3(n_371),
.B(n_372),
.Y(n_2884)
);

OAI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2627),
.A2(n_374),
.B(n_375),
.Y(n_2885)
);

INVx3_ASAP7_75t_L g2886 ( 
.A(n_2530),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2416),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2621),
.A2(n_374),
.B(n_375),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_SL g2889 ( 
.A(n_2367),
.B(n_724),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2393),
.B(n_376),
.Y(n_2890)
);

OAI21x1_ASAP7_75t_L g2891 ( 
.A1(n_2603),
.A2(n_376),
.B(n_377),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2404),
.B(n_376),
.Y(n_2892)
);

INVx3_ASAP7_75t_L g2893 ( 
.A(n_2530),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2628),
.A2(n_377),
.B(n_378),
.Y(n_2894)
);

NOR2x1_ASAP7_75t_SL g2895 ( 
.A(n_2567),
.B(n_377),
.Y(n_2895)
);

AND2x4_ASAP7_75t_L g2896 ( 
.A(n_2531),
.B(n_378),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2567),
.Y(n_2897)
);

AOI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2288),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_2898)
);

OR2x6_ASAP7_75t_L g2899 ( 
.A(n_2735),
.B(n_379),
.Y(n_2899)
);

BUFx6f_ASAP7_75t_L g2900 ( 
.A(n_2567),
.Y(n_2900)
);

INVx3_ASAP7_75t_L g2901 ( 
.A(n_2574),
.Y(n_2901)
);

INVx2_ASAP7_75t_SL g2902 ( 
.A(n_2348),
.Y(n_2902)
);

A2O1A1Ixp33_ASAP7_75t_L g2903 ( 
.A1(n_2413),
.A2(n_381),
.B(n_379),
.C(n_380),
.Y(n_2903)
);

NOR3xp33_ASAP7_75t_L g2904 ( 
.A(n_2366),
.B(n_380),
.C(n_382),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2611),
.Y(n_2905)
);

OAI21x1_ASAP7_75t_L g2906 ( 
.A1(n_2616),
.A2(n_382),
.B(n_383),
.Y(n_2906)
);

AO31x2_ASAP7_75t_L g2907 ( 
.A1(n_2407),
.A2(n_384),
.A3(n_382),
.B(n_383),
.Y(n_2907)
);

OAI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2290),
.A2(n_383),
.B(n_384),
.Y(n_2908)
);

AND2x4_ASAP7_75t_L g2909 ( 
.A(n_2531),
.B(n_384),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2414),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2346),
.Y(n_2911)
);

AOI21x1_ASAP7_75t_SL g2912 ( 
.A1(n_2479),
.A2(n_385),
.B(n_387),
.Y(n_2912)
);

INVx1_ASAP7_75t_SL g2913 ( 
.A(n_2414),
.Y(n_2913)
);

OAI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2636),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_2914)
);

O2A1O1Ixp5_ASAP7_75t_L g2915 ( 
.A1(n_2499),
.A2(n_390),
.B(n_388),
.C(n_389),
.Y(n_2915)
);

INVx2_ASAP7_75t_SL g2916 ( 
.A(n_2473),
.Y(n_2916)
);

OAI21x1_ASAP7_75t_SL g2917 ( 
.A1(n_2409),
.A2(n_388),
.B(n_389),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2632),
.A2(n_389),
.B(n_390),
.Y(n_2918)
);

OAI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2318),
.A2(n_391),
.B(n_392),
.Y(n_2919)
);

OAI21x1_ASAP7_75t_L g2920 ( 
.A1(n_2465),
.A2(n_391),
.B(n_392),
.Y(n_2920)
);

OAI22x1_ASAP7_75t_L g2921 ( 
.A1(n_2698),
.A2(n_395),
.B1(n_391),
.B2(n_393),
.Y(n_2921)
);

AOI21xp33_ASAP7_75t_L g2922 ( 
.A1(n_2635),
.A2(n_393),
.B(n_395),
.Y(n_2922)
);

INVx4_ASAP7_75t_L g2923 ( 
.A(n_2714),
.Y(n_2923)
);

AOI22xp33_ASAP7_75t_SL g2924 ( 
.A1(n_2515),
.A2(n_397),
.B1(n_393),
.B2(n_396),
.Y(n_2924)
);

OAI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2640),
.A2(n_396),
.B(n_398),
.Y(n_2925)
);

A2O1A1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2415),
.A2(n_399),
.B(n_396),
.C(n_398),
.Y(n_2926)
);

AND2x4_ASAP7_75t_L g2927 ( 
.A(n_2714),
.B(n_398),
.Y(n_2927)
);

OAI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2645),
.A2(n_400),
.B(n_401),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_SL g2929 ( 
.A1(n_2574),
.A2(n_2620),
.B(n_2577),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2652),
.A2(n_400),
.B(n_401),
.Y(n_2930)
);

OAI21x1_ASAP7_75t_L g2931 ( 
.A1(n_2282),
.A2(n_400),
.B(n_401),
.Y(n_2931)
);

INVx4_ASAP7_75t_L g2932 ( 
.A(n_2737),
.Y(n_2932)
);

BUFx12f_ASAP7_75t_L g2933 ( 
.A(n_2285),
.Y(n_2933)
);

AOI21xp33_ASAP7_75t_L g2934 ( 
.A1(n_2654),
.A2(n_402),
.B(n_403),
.Y(n_2934)
);

CKINVDCx20_ASAP7_75t_R g2935 ( 
.A(n_2468),
.Y(n_2935)
);

OAI22x1_ASAP7_75t_L g2936 ( 
.A1(n_2716),
.A2(n_404),
.B1(n_402),
.B2(n_403),
.Y(n_2936)
);

AO31x2_ASAP7_75t_L g2937 ( 
.A1(n_2496),
.A2(n_408),
.A3(n_406),
.B(n_407),
.Y(n_2937)
);

INVx3_ASAP7_75t_L g2938 ( 
.A(n_2574),
.Y(n_2938)
);

NOR2xp67_ASAP7_75t_L g2939 ( 
.A(n_2737),
.B(n_409),
.Y(n_2939)
);

NAND2x1p5_ASAP7_75t_L g2940 ( 
.A(n_2473),
.B(n_2432),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2687),
.A2(n_409),
.B(n_410),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_L g2942 ( 
.A(n_2365),
.B(n_411),
.Y(n_2942)
);

AO221x2_ASAP7_75t_L g2943 ( 
.A1(n_2526),
.A2(n_414),
.B1(n_411),
.B2(n_413),
.C(n_415),
.Y(n_2943)
);

AOI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2696),
.A2(n_413),
.B(n_414),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2425),
.B(n_413),
.Y(n_2945)
);

AOI22xp5_ASAP7_75t_L g2946 ( 
.A1(n_2642),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_2946)
);

OAI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2704),
.A2(n_416),
.B(n_417),
.Y(n_2947)
);

INVxp67_ASAP7_75t_SL g2948 ( 
.A(n_2577),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2455),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2457),
.Y(n_2950)
);

OR2x2_ASAP7_75t_L g2951 ( 
.A(n_2292),
.B(n_418),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2520),
.Y(n_2952)
);

BUFx3_ASAP7_75t_L g2953 ( 
.A(n_2440),
.Y(n_2953)
);

HB1xp67_ASAP7_75t_L g2954 ( 
.A(n_2391),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_SL g2955 ( 
.A1(n_2577),
.A2(n_419),
.B(n_420),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2722),
.A2(n_2725),
.B(n_2724),
.Y(n_2956)
);

OAI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2727),
.A2(n_419),
.B(n_421),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2738),
.A2(n_421),
.B(n_422),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2374),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2381),
.Y(n_2960)
);

AO31x2_ASAP7_75t_L g2961 ( 
.A1(n_2533),
.A2(n_423),
.A3(n_421),
.B(n_422),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2394),
.Y(n_2962)
);

HB1xp67_ASAP7_75t_L g2963 ( 
.A(n_2498),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2344),
.B(n_424),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2562),
.B(n_424),
.Y(n_2965)
);

INVx5_ASAP7_75t_L g2966 ( 
.A(n_2272),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2580),
.B(n_425),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2306),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2583),
.B(n_427),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2587),
.B(n_428),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2420),
.Y(n_2971)
);

OAI21x1_ASAP7_75t_L g2972 ( 
.A1(n_2351),
.A2(n_429),
.B(n_430),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2593),
.B(n_431),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2610),
.B(n_431),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_2276),
.B(n_431),
.Y(n_2975)
);

AOI21xp5_ASAP7_75t_L g2976 ( 
.A1(n_2434),
.A2(n_432),
.B(n_433),
.Y(n_2976)
);

BUFx2_ASAP7_75t_L g2977 ( 
.A(n_2502),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_SL g2978 ( 
.A(n_2296),
.B(n_725),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2641),
.B(n_434),
.Y(n_2979)
);

OR2x2_ASAP7_75t_L g2980 ( 
.A(n_2590),
.B(n_435),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2643),
.B(n_436),
.Y(n_2981)
);

AOI21x1_ASAP7_75t_SL g2982 ( 
.A1(n_2454),
.A2(n_436),
.B(n_437),
.Y(n_2982)
);

AOI21xp5_ASAP7_75t_L g2983 ( 
.A1(n_2304),
.A2(n_438),
.B(n_439),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2657),
.B(n_439),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2667),
.B(n_440),
.Y(n_2985)
);

A2O1A1Ixp33_ASAP7_75t_L g2986 ( 
.A1(n_2424),
.A2(n_442),
.B(n_440),
.C(n_441),
.Y(n_2986)
);

INVx3_ASAP7_75t_SL g2987 ( 
.A(n_2646),
.Y(n_2987)
);

NOR2xp33_ASAP7_75t_L g2988 ( 
.A(n_2284),
.B(n_443),
.Y(n_2988)
);

AO31x2_ASAP7_75t_L g2989 ( 
.A1(n_2599),
.A2(n_445),
.A3(n_443),
.B(n_444),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2294),
.B(n_445),
.Y(n_2990)
);

OAI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2311),
.A2(n_446),
.B(n_447),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2300),
.B(n_446),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_2300),
.B(n_447),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2504),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2692),
.B(n_2674),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2498),
.B(n_449),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2301),
.B(n_450),
.Y(n_2997)
);

AOI21xp5_ASAP7_75t_L g2998 ( 
.A1(n_2347),
.A2(n_452),
.B(n_453),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2301),
.B(n_452),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2523),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2303),
.B(n_454),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2376),
.A2(n_455),
.B(n_456),
.Y(n_3002)
);

OAI21xp5_ASAP7_75t_L g3003 ( 
.A1(n_2471),
.A2(n_455),
.B(n_456),
.Y(n_3003)
);

BUFx3_ASAP7_75t_L g3004 ( 
.A(n_2655),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2433),
.Y(n_3005)
);

INVxp67_ASAP7_75t_L g3006 ( 
.A(n_2332),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2500),
.B(n_457),
.Y(n_3007)
);

INVx3_ASAP7_75t_L g3008 ( 
.A(n_2620),
.Y(n_3008)
);

OR2x6_ASAP7_75t_L g3009 ( 
.A(n_2495),
.B(n_457),
.Y(n_3009)
);

OR2x2_ASAP7_75t_L g3010 ( 
.A(n_2387),
.B(n_458),
.Y(n_3010)
);

OAI22x1_ASAP7_75t_L g3011 ( 
.A1(n_2720),
.A2(n_460),
.B1(n_458),
.B2(n_459),
.Y(n_3011)
);

AOI21xp5_ASAP7_75t_L g3012 ( 
.A1(n_2379),
.A2(n_460),
.B(n_461),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2511),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2396),
.B(n_460),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2371),
.B(n_462),
.Y(n_3015)
);

INVx3_ASAP7_75t_L g3016 ( 
.A(n_2620),
.Y(n_3016)
);

INVx4_ASAP7_75t_L g3017 ( 
.A(n_2488),
.Y(n_3017)
);

OR2x6_ASAP7_75t_L g3018 ( 
.A(n_2524),
.B(n_462),
.Y(n_3018)
);

CKINVDCx20_ASAP7_75t_R g3019 ( 
.A(n_2448),
.Y(n_3019)
);

AO31x2_ASAP7_75t_L g3020 ( 
.A1(n_2607),
.A2(n_465),
.A3(n_463),
.B(n_464),
.Y(n_3020)
);

AOI21xp33_ASAP7_75t_L g3021 ( 
.A1(n_2419),
.A2(n_463),
.B(n_464),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2426),
.B(n_466),
.Y(n_3022)
);

AOI21xp5_ASAP7_75t_L g3023 ( 
.A1(n_2446),
.A2(n_466),
.B(n_467),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2516),
.Y(n_3024)
);

AO31x2_ASAP7_75t_L g3025 ( 
.A1(n_2614),
.A2(n_469),
.A3(n_466),
.B(n_468),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2521),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2389),
.B(n_470),
.Y(n_3027)
);

OAI21x1_ASAP7_75t_L g3028 ( 
.A1(n_2532),
.A2(n_471),
.B(n_472),
.Y(n_3028)
);

AND2x4_ASAP7_75t_L g3029 ( 
.A(n_2514),
.B(n_471),
.Y(n_3029)
);

OAI21xp5_ASAP7_75t_L g3030 ( 
.A1(n_2452),
.A2(n_472),
.B(n_473),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2399),
.B(n_472),
.Y(n_3031)
);

OAI21xp5_ASAP7_75t_L g3032 ( 
.A1(n_2472),
.A2(n_473),
.B(n_474),
.Y(n_3032)
);

AO31x2_ASAP7_75t_L g3033 ( 
.A1(n_2615),
.A2(n_475),
.A3(n_473),
.B(n_474),
.Y(n_3033)
);

AND2x6_ASAP7_75t_L g3034 ( 
.A(n_2672),
.B(n_474),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2720),
.Y(n_3035)
);

AOI22xp5_ASAP7_75t_L g3036 ( 
.A1(n_2281),
.A2(n_477),
.B1(n_475),
.B2(n_476),
.Y(n_3036)
);

BUFx2_ASAP7_75t_L g3037 ( 
.A(n_2633),
.Y(n_3037)
);

NOR2xp33_ASAP7_75t_SL g3038 ( 
.A(n_2272),
.B(n_475),
.Y(n_3038)
);

AOI21xp5_ASAP7_75t_L g3039 ( 
.A1(n_2575),
.A2(n_476),
.B(n_477),
.Y(n_3039)
);

AND2x4_ASAP7_75t_L g3040 ( 
.A(n_2517),
.B(n_476),
.Y(n_3040)
);

AND2x2_ASAP7_75t_L g3041 ( 
.A(n_2385),
.B(n_477),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2403),
.B(n_478),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_L g3043 ( 
.A(n_2483),
.B(n_478),
.Y(n_3043)
);

OAI22xp5_ASAP7_75t_L g3044 ( 
.A1(n_2528),
.A2(n_480),
.B1(n_478),
.B2(n_479),
.Y(n_3044)
);

AOI22xp5_ASAP7_75t_L g3045 ( 
.A1(n_2297),
.A2(n_481),
.B1(n_479),
.B2(n_480),
.Y(n_3045)
);

OAI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2333),
.A2(n_2339),
.B(n_2295),
.Y(n_3046)
);

OAI21x1_ASAP7_75t_L g3047 ( 
.A1(n_2537),
.A2(n_479),
.B(n_481),
.Y(n_3047)
);

OAI21x1_ASAP7_75t_L g3048 ( 
.A1(n_2540),
.A2(n_482),
.B(n_483),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2466),
.Y(n_3049)
);

BUFx4f_ASAP7_75t_SL g3050 ( 
.A(n_2508),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_L g3051 ( 
.A1(n_2546),
.A2(n_482),
.B(n_483),
.Y(n_3051)
);

OAI21xp5_ASAP7_75t_L g3052 ( 
.A1(n_2427),
.A2(n_482),
.B(n_484),
.Y(n_3052)
);

AOI21xp5_ASAP7_75t_L g3053 ( 
.A1(n_2556),
.A2(n_485),
.B(n_486),
.Y(n_3053)
);

OAI21x1_ASAP7_75t_L g3054 ( 
.A1(n_2558),
.A2(n_485),
.B(n_486),
.Y(n_3054)
);

NAND2x1p5_ASAP7_75t_L g3055 ( 
.A(n_2672),
.B(n_485),
.Y(n_3055)
);

AOI21x1_ASAP7_75t_SL g3056 ( 
.A1(n_2484),
.A2(n_486),
.B(n_487),
.Y(n_3056)
);

OAI21xp5_ASAP7_75t_L g3057 ( 
.A1(n_2430),
.A2(n_487),
.B(n_488),
.Y(n_3057)
);

INVx4_ASAP7_75t_L g3058 ( 
.A(n_2272),
.Y(n_3058)
);

NAND2xp33_ASAP7_75t_L g3059 ( 
.A(n_2272),
.B(n_488),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2325),
.B(n_488),
.Y(n_3060)
);

AND2x2_ASAP7_75t_L g3061 ( 
.A(n_2279),
.B(n_489),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2279),
.B(n_489),
.Y(n_3062)
);

OAI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2442),
.A2(n_490),
.B(n_491),
.Y(n_3063)
);

BUFx3_ASAP7_75t_L g3064 ( 
.A(n_2512),
.Y(n_3064)
);

INVx2_ASAP7_75t_SL g3065 ( 
.A(n_2501),
.Y(n_3065)
);

OAI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2443),
.A2(n_490),
.B(n_491),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2560),
.A2(n_490),
.B(n_491),
.Y(n_3067)
);

A2O1A1Ixp33_ASAP7_75t_L g3068 ( 
.A1(n_2437),
.A2(n_494),
.B(n_492),
.C(n_493),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2400),
.B(n_494),
.Y(n_3069)
);

AOI21x1_ASAP7_75t_SL g3070 ( 
.A1(n_2482),
.A2(n_495),
.B(n_496),
.Y(n_3070)
);

AOI21xp5_ASAP7_75t_L g3071 ( 
.A1(n_2570),
.A2(n_495),
.B(n_496),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2740),
.B(n_495),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2334),
.B(n_497),
.Y(n_3073)
);

AOI21xp5_ASAP7_75t_L g3074 ( 
.A1(n_2573),
.A2(n_497),
.B(n_498),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2565),
.B(n_497),
.Y(n_3075)
);

O2A1O1Ixp5_ASAP7_75t_L g3076 ( 
.A1(n_2463),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2658),
.B(n_498),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2662),
.B(n_499),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2579),
.A2(n_499),
.B(n_500),
.Y(n_3079)
);

AOI21xp5_ASAP7_75t_L g3080 ( 
.A1(n_2582),
.A2(n_500),
.B(n_501),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2686),
.B(n_501),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2688),
.B(n_502),
.Y(n_3082)
);

AOI21x1_ASAP7_75t_L g3083 ( 
.A1(n_2460),
.A2(n_502),
.B(n_503),
.Y(n_3083)
);

BUFx4f_ASAP7_75t_L g3084 ( 
.A(n_2673),
.Y(n_3084)
);

OAI22xp5_ASAP7_75t_L g3085 ( 
.A1(n_2549),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_3085)
);

INVx3_ASAP7_75t_L g3086 ( 
.A(n_2673),
.Y(n_3086)
);

INVxp67_ASAP7_75t_L g3087 ( 
.A(n_2436),
.Y(n_3087)
);

OAI21xp5_ASAP7_75t_L g3088 ( 
.A1(n_2421),
.A2(n_503),
.B(n_504),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2694),
.B(n_505),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2697),
.B(n_505),
.Y(n_3090)
);

OAI21x1_ASAP7_75t_L g3091 ( 
.A1(n_2597),
.A2(n_505),
.B(n_506),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2701),
.B(n_506),
.Y(n_3092)
);

OAI21x1_ASAP7_75t_L g3093 ( 
.A1(n_2598),
.A2(n_506),
.B(n_507),
.Y(n_3093)
);

HB1xp67_ASAP7_75t_L g3094 ( 
.A(n_2566),
.Y(n_3094)
);

BUFx2_ASAP7_75t_L g3095 ( 
.A(n_2438),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2733),
.Y(n_3096)
);

CKINVDCx20_ASAP7_75t_R g3097 ( 
.A(n_2510),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2706),
.B(n_507),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_L g3099 ( 
.A(n_2709),
.B(n_2289),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2461),
.B(n_508),
.Y(n_3100)
);

BUFx8_ASAP7_75t_L g3101 ( 
.A(n_2326),
.Y(n_3101)
);

OAI21xp5_ASAP7_75t_L g3102 ( 
.A1(n_2361),
.A2(n_508),
.B(n_509),
.Y(n_3102)
);

OAI21xp5_ASAP7_75t_L g3103 ( 
.A1(n_2363),
.A2(n_510),
.B(n_511),
.Y(n_3103)
);

BUFx3_ASAP7_75t_L g3104 ( 
.A(n_2517),
.Y(n_3104)
);

AOI21x1_ASAP7_75t_L g3105 ( 
.A1(n_2604),
.A2(n_510),
.B(n_511),
.Y(n_3105)
);

OAI21x1_ASAP7_75t_L g3106 ( 
.A1(n_2606),
.A2(n_510),
.B(n_511),
.Y(n_3106)
);

NAND2x1p5_ASAP7_75t_L g3107 ( 
.A(n_2733),
.B(n_512),
.Y(n_3107)
);

AOI21x1_ASAP7_75t_L g3108 ( 
.A1(n_2609),
.A2(n_512),
.B(n_513),
.Y(n_3108)
);

OAI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2369),
.A2(n_514),
.B(n_515),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2384),
.B(n_514),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_SL g3111 ( 
.A(n_2684),
.B(n_726),
.Y(n_3111)
);

OAI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_2578),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.Y(n_3112)
);

INVx5_ASAP7_75t_L g3113 ( 
.A(n_2733),
.Y(n_3113)
);

A2O1A1Ixp33_ASAP7_75t_L g3114 ( 
.A1(n_2439),
.A2(n_519),
.B(n_516),
.C(n_518),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2617),
.A2(n_519),
.B(n_520),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2469),
.Y(n_3116)
);

AOI21x1_ASAP7_75t_SL g3117 ( 
.A1(n_2309),
.A2(n_2324),
.B(n_2319),
.Y(n_3117)
);

NOR2xp33_ASAP7_75t_L g3118 ( 
.A(n_2299),
.B(n_519),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_2619),
.A2(n_520),
.B(n_521),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2373),
.B(n_522),
.Y(n_3120)
);

INVx3_ASAP7_75t_L g3121 ( 
.A(n_2429),
.Y(n_3121)
);

AOI221xp5_ASAP7_75t_L g3122 ( 
.A1(n_2572),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.C(n_528),
.Y(n_3122)
);

AND2x4_ASAP7_75t_L g3123 ( 
.A(n_2480),
.B(n_527),
.Y(n_3123)
);

OAI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2372),
.A2(n_527),
.B(n_529),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2444),
.B(n_529),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2589),
.Y(n_3126)
);

OAI22xp5_ASAP7_75t_L g3127 ( 
.A1(n_2595),
.A2(n_532),
.B1(n_530),
.B2(n_531),
.Y(n_3127)
);

AND2x2_ASAP7_75t_SL g3128 ( 
.A(n_2353),
.B(n_530),
.Y(n_3128)
);

BUFx2_ASAP7_75t_SL g3129 ( 
.A(n_2703),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_2480),
.B(n_533),
.Y(n_3130)
);

A2O1A1Ixp33_ASAP7_75t_L g3131 ( 
.A1(n_2638),
.A2(n_2656),
.B(n_2660),
.C(n_2650),
.Y(n_3131)
);

INVx2_ASAP7_75t_SL g3132 ( 
.A(n_2519),
.Y(n_3132)
);

OAI21x1_ASAP7_75t_L g3133 ( 
.A1(n_2666),
.A2(n_534),
.B(n_535),
.Y(n_3133)
);

AOI21xp33_ASAP7_75t_L g3134 ( 
.A1(n_2659),
.A2(n_537),
.B(n_538),
.Y(n_3134)
);

AOI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_2669),
.A2(n_538),
.B(n_539),
.Y(n_3135)
);

AO31x2_ASAP7_75t_L g3136 ( 
.A1(n_2679),
.A2(n_2702),
.A3(n_2690),
.B(n_2739),
.Y(n_3136)
);

AOI221xp5_ASAP7_75t_SL g3137 ( 
.A1(n_2478),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.C(n_542),
.Y(n_3137)
);

BUFx2_ASAP7_75t_L g3138 ( 
.A(n_2467),
.Y(n_3138)
);

AND3x2_ASAP7_75t_L g3139 ( 
.A(n_2486),
.B(n_540),
.C(n_541),
.Y(n_3139)
);

AOI21xp5_ASAP7_75t_L g3140 ( 
.A1(n_2671),
.A2(n_541),
.B(n_542),
.Y(n_3140)
);

AO31x2_ASAP7_75t_L g3141 ( 
.A1(n_2678),
.A2(n_545),
.A3(n_543),
.B(n_544),
.Y(n_3141)
);

BUFx4f_ASAP7_75t_L g3142 ( 
.A(n_2429),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2591),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2497),
.B(n_546),
.Y(n_3144)
);

AOI21xp5_ASAP7_75t_SL g3145 ( 
.A1(n_2429),
.A2(n_546),
.B(n_547),
.Y(n_3145)
);

A2O1A1Ixp33_ASAP7_75t_L g3146 ( 
.A1(n_2691),
.A2(n_548),
.B(n_546),
.C(n_547),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2487),
.B(n_549),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2602),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_2314),
.B(n_2317),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2283),
.B(n_550),
.Y(n_3150)
);

BUFx2_ASAP7_75t_L g3151 ( 
.A(n_2467),
.Y(n_3151)
);

A2O1A1Ixp33_ASAP7_75t_L g3152 ( 
.A1(n_2693),
.A2(n_552),
.B(n_550),
.C(n_551),
.Y(n_3152)
);

AOI211x1_ASAP7_75t_L g3153 ( 
.A1(n_2522),
.A2(n_553),
.B(n_551),
.C(n_552),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2467),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2490),
.B(n_553),
.Y(n_3155)
);

OA22x2_ASAP7_75t_L g3156 ( 
.A1(n_2644),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2494),
.B(n_554),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2370),
.B(n_554),
.Y(n_3158)
);

A2O1A1Ixp33_ASAP7_75t_L g3159 ( 
.A1(n_2699),
.A2(n_557),
.B(n_555),
.C(n_556),
.Y(n_3159)
);

AO31x2_ASAP7_75t_L g3160 ( 
.A1(n_2713),
.A2(n_557),
.A3(n_555),
.B(n_556),
.Y(n_3160)
);

OAI21xp5_ASAP7_75t_L g3161 ( 
.A1(n_2717),
.A2(n_556),
.B(n_558),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2336),
.B(n_558),
.Y(n_3162)
);

NAND2x1_ASAP7_75t_L g3163 ( 
.A(n_2485),
.B(n_559),
.Y(n_3163)
);

AO31x2_ASAP7_75t_L g3164 ( 
.A1(n_2730),
.A2(n_562),
.A3(n_560),
.B(n_561),
.Y(n_3164)
);

NAND3xp33_ASAP7_75t_L g3165 ( 
.A(n_2539),
.B(n_560),
.C(n_561),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2397),
.B(n_562),
.Y(n_3166)
);

OAI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2734),
.A2(n_563),
.B(n_564),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2447),
.B(n_563),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2321),
.B(n_564),
.Y(n_3169)
);

AND2x4_ASAP7_75t_L g3170 ( 
.A(n_2513),
.B(n_565),
.Y(n_3170)
);

BUFx3_ASAP7_75t_L g3171 ( 
.A(n_2464),
.Y(n_3171)
);

OAI22x1_ASAP7_75t_L g3172 ( 
.A1(n_2422),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_2445),
.Y(n_3173)
);

AOI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2754),
.A2(n_2828),
.B1(n_2787),
.B2(n_3035),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2911),
.B(n_2624),
.Y(n_3175)
);

AOI22xp5_ASAP7_75t_L g3176 ( 
.A1(n_2843),
.A2(n_2588),
.B1(n_2685),
.B2(n_2592),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2748),
.B(n_2647),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_3061),
.B(n_3062),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2765),
.Y(n_3179)
);

AOI22xp5_ASAP7_75t_L g3180 ( 
.A1(n_2995),
.A2(n_2298),
.B1(n_2449),
.B2(n_2453),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2772),
.Y(n_3181)
);

AOI22xp33_ASAP7_75t_L g3182 ( 
.A1(n_3128),
.A2(n_2481),
.B1(n_2503),
.B2(n_2648),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2798),
.B(n_2653),
.Y(n_3183)
);

AOI22xp33_ASAP7_75t_L g3184 ( 
.A1(n_2943),
.A2(n_2665),
.B1(n_2675),
.B2(n_2663),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2956),
.A2(n_2601),
.B(n_2600),
.Y(n_3185)
);

AND2x4_ASAP7_75t_L g3186 ( 
.A(n_2760),
.B(n_2518),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2777),
.B(n_2700),
.Y(n_3187)
);

BUFx12f_ASAP7_75t_L g3188 ( 
.A(n_2743),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3126),
.B(n_2705),
.Y(n_3189)
);

AND2x4_ASAP7_75t_L g3190 ( 
.A(n_2760),
.B(n_2386),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2807),
.Y(n_3191)
);

CKINVDCx5p33_ASAP7_75t_R g3192 ( 
.A(n_2751),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2945),
.B(n_2328),
.Y(n_3193)
);

OR2x2_ASAP7_75t_L g3194 ( 
.A(n_2980),
.B(n_2708),
.Y(n_3194)
);

BUFx2_ASAP7_75t_L g3195 ( 
.A(n_3034),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2808),
.Y(n_3196)
);

INVx1_ASAP7_75t_SL g3197 ( 
.A(n_3019),
.Y(n_3197)
);

AND2x4_ASAP7_75t_L g3198 ( 
.A(n_2760),
.B(n_2392),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3143),
.B(n_2728),
.Y(n_3199)
);

HB1xp67_ASAP7_75t_L g3200 ( 
.A(n_2830),
.Y(n_3200)
);

CKINVDCx20_ASAP7_75t_R g3201 ( 
.A(n_2935),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_L g3202 ( 
.A(n_2766),
.B(n_2412),
.Y(n_3202)
);

AOI21xp5_ASAP7_75t_L g3203 ( 
.A1(n_3131),
.A2(n_2715),
.B(n_2664),
.Y(n_3203)
);

AOI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_3005),
.A2(n_2715),
.B(n_2664),
.Y(n_3204)
);

INVx2_ASAP7_75t_L g3205 ( 
.A(n_2810),
.Y(n_3205)
);

BUFx6f_ASAP7_75t_L g3206 ( 
.A(n_2953),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2804),
.Y(n_3207)
);

AND2x4_ASAP7_75t_L g3208 ( 
.A(n_3017),
.B(n_2354),
.Y(n_3208)
);

OAI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_2963),
.A2(n_2350),
.B1(n_2408),
.B2(n_2450),
.Y(n_3209)
);

INVx2_ASAP7_75t_SL g3210 ( 
.A(n_3050),
.Y(n_3210)
);

INVx2_ASAP7_75t_SL g3211 ( 
.A(n_2743),
.Y(n_3211)
);

CKINVDCx5p33_ASAP7_75t_R g3212 ( 
.A(n_2849),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_2923),
.Y(n_3213)
);

NAND2x1p5_ASAP7_75t_L g3214 ( 
.A(n_2860),
.B(n_2302),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3148),
.B(n_2493),
.Y(n_3215)
);

INVx4_ASAP7_75t_L g3216 ( 
.A(n_2860),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2813),
.Y(n_3217)
);

OAI22xp33_ASAP7_75t_L g3218 ( 
.A1(n_3009),
.A2(n_2576),
.B1(n_2623),
.B2(n_2383),
.Y(n_3218)
);

INVx8_ASAP7_75t_L g3219 ( 
.A(n_2838),
.Y(n_3219)
);

INVx3_ASAP7_75t_L g3220 ( 
.A(n_2923),
.Y(n_3220)
);

INVx1_ASAP7_75t_SL g3221 ( 
.A(n_3000),
.Y(n_3221)
);

INVx3_ASAP7_75t_L g3222 ( 
.A(n_2932),
.Y(n_3222)
);

INVx4_ASAP7_75t_L g3223 ( 
.A(n_2870),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2816),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2833),
.B(n_2847),
.Y(n_3225)
);

INVx2_ASAP7_75t_SL g3226 ( 
.A(n_2873),
.Y(n_3226)
);

INVxp67_ASAP7_75t_L g3227 ( 
.A(n_2756),
.Y(n_3227)
);

BUFx2_ASAP7_75t_L g3228 ( 
.A(n_3034),
.Y(n_3228)
);

CKINVDCx6p67_ASAP7_75t_R g3229 ( 
.A(n_2987),
.Y(n_3229)
);

O2A1O1Ixp33_ASAP7_75t_L g3230 ( 
.A1(n_3149),
.A2(n_2474),
.B(n_2382),
.C(n_2729),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2824),
.Y(n_3231)
);

BUFx8_ASAP7_75t_SL g3232 ( 
.A(n_2933),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2845),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3009),
.A2(n_2736),
.B1(n_2731),
.B2(n_2507),
.Y(n_3234)
);

OAI21xp33_ASAP7_75t_L g3235 ( 
.A1(n_2924),
.A2(n_2476),
.B(n_2470),
.Y(n_3235)
);

OAI22xp5_ASAP7_75t_L g3236 ( 
.A1(n_2899),
.A2(n_2506),
.B1(n_2406),
.B2(n_2410),
.Y(n_3236)
);

CKINVDCx9p33_ASAP7_75t_R g3237 ( 
.A(n_3037),
.Y(n_3237)
);

OR2x6_ASAP7_75t_L g3238 ( 
.A(n_2902),
.B(n_2477),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_3084),
.Y(n_3239)
);

CKINVDCx5p33_ASAP7_75t_R g3240 ( 
.A(n_2913),
.Y(n_3240)
);

AND2x2_ASAP7_75t_L g3241 ( 
.A(n_2996),
.B(n_567),
.Y(n_3241)
);

O2A1O1Ixp33_ASAP7_75t_L g3242 ( 
.A1(n_3087),
.A2(n_2505),
.B(n_2475),
.C(n_2608),
.Y(n_3242)
);

CKINVDCx20_ASAP7_75t_R g3243 ( 
.A(n_2910),
.Y(n_3243)
);

INVx4_ASAP7_75t_L g3244 ( 
.A(n_3017),
.Y(n_3244)
);

OAI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2899),
.A2(n_2402),
.B1(n_2405),
.B2(n_2377),
.Y(n_3245)
);

BUFx4f_ASAP7_75t_L g3246 ( 
.A(n_2838),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2855),
.B(n_2451),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2868),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_2864),
.B(n_2459),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2875),
.Y(n_3250)
);

INVx1_ASAP7_75t_L g3251 ( 
.A(n_2878),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_2742),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2880),
.B(n_2489),
.Y(n_3253)
);

BUFx6f_ASAP7_75t_L g3254 ( 
.A(n_3084),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_2932),
.B(n_2458),
.Y(n_3255)
);

OR2x6_ASAP7_75t_L g3256 ( 
.A(n_2865),
.B(n_568),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_2836),
.B(n_568),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2839),
.B(n_569),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2952),
.Y(n_3259)
);

BUFx6f_ASAP7_75t_SL g3260 ( 
.A(n_3004),
.Y(n_3260)
);

BUFx6f_ASAP7_75t_L g3261 ( 
.A(n_3113),
.Y(n_3261)
);

INVx5_ASAP7_75t_L g3262 ( 
.A(n_3034),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2876),
.B(n_2747),
.Y(n_3263)
);

BUFx2_ASAP7_75t_L g3264 ( 
.A(n_3058),
.Y(n_3264)
);

AOI22xp33_ASAP7_75t_L g3265 ( 
.A1(n_3029),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3265)
);

O2A1O1Ixp33_ASAP7_75t_L g3266 ( 
.A1(n_2857),
.A2(n_572),
.B(n_570),
.C(n_571),
.Y(n_3266)
);

OAI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_2946),
.A2(n_576),
.B1(n_573),
.B2(n_575),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2851),
.B(n_575),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2971),
.B(n_576),
.Y(n_3269)
);

CKINVDCx16_ASAP7_75t_R g3270 ( 
.A(n_2797),
.Y(n_3270)
);

AOI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_3059),
.A2(n_576),
.B(n_577),
.Y(n_3271)
);

O2A1O1Ixp5_ASAP7_75t_L g3272 ( 
.A1(n_2861),
.A2(n_579),
.B(n_577),
.C(n_578),
.Y(n_3272)
);

AOI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3097),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_3273)
);

BUFx3_ASAP7_75t_L g3274 ( 
.A(n_2811),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_2867),
.B(n_578),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_SL g3276 ( 
.A(n_3038),
.B(n_579),
.Y(n_3276)
);

NOR2x1p5_ASAP7_75t_L g3277 ( 
.A(n_3010),
.B(n_581),
.Y(n_3277)
);

O2A1O1Ixp5_ASAP7_75t_SL g3278 ( 
.A1(n_3094),
.A2(n_728),
.B(n_729),
.C(n_727),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2872),
.B(n_581),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_2788),
.B(n_581),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_2750),
.Y(n_3281)
);

AOI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_2929),
.A2(n_582),
.B(n_583),
.Y(n_3282)
);

INVx2_ASAP7_75t_L g3283 ( 
.A(n_2769),
.Y(n_3283)
);

INVxp67_ASAP7_75t_L g3284 ( 
.A(n_2977),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_2788),
.B(n_582),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_2789),
.B(n_583),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_SL g3287 ( 
.A(n_2966),
.B(n_3058),
.Y(n_3287)
);

BUFx6f_ASAP7_75t_L g3288 ( 
.A(n_3113),
.Y(n_3288)
);

OR2x2_ASAP7_75t_L g3289 ( 
.A(n_2745),
.B(n_583),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_L g3290 ( 
.A(n_2768),
.B(n_584),
.Y(n_3290)
);

NAND2x1p5_ASAP7_75t_L g3291 ( 
.A(n_2966),
.B(n_584),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_2789),
.B(n_585),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_2949),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_2990),
.B(n_585),
.Y(n_3294)
);

AOI22xp5_ASAP7_75t_L g3295 ( 
.A1(n_3041),
.A2(n_587),
.B1(n_585),
.B2(n_586),
.Y(n_3295)
);

INVx3_ASAP7_75t_SL g3296 ( 
.A(n_2811),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2799),
.Y(n_3297)
);

BUFx12f_ASAP7_75t_L g3298 ( 
.A(n_3095),
.Y(n_3298)
);

INVx6_ASAP7_75t_L g3299 ( 
.A(n_3064),
.Y(n_3299)
);

AOI22xp5_ASAP7_75t_L g3300 ( 
.A1(n_2975),
.A2(n_588),
.B1(n_586),
.B2(n_587),
.Y(n_3300)
);

INVxp67_ASAP7_75t_L g3301 ( 
.A(n_2942),
.Y(n_3301)
);

BUFx10_ASAP7_75t_L g3302 ( 
.A(n_2896),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_2940),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2799),
.Y(n_3304)
);

HB1xp67_ASAP7_75t_L g3305 ( 
.A(n_3040),
.Y(n_3305)
);

NAND2x1p5_ASAP7_75t_L g3306 ( 
.A(n_2966),
.B(n_588),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3007),
.Y(n_3307)
);

OR2x6_ASAP7_75t_SL g3308 ( 
.A(n_2822),
.B(n_589),
.Y(n_3308)
);

HB1xp67_ASAP7_75t_L g3309 ( 
.A(n_3040),
.Y(n_3309)
);

A2O1A1Ixp33_ASAP7_75t_L g3310 ( 
.A1(n_2919),
.A2(n_592),
.B(n_590),
.C(n_591),
.Y(n_3310)
);

HB1xp67_ASAP7_75t_L g3311 ( 
.A(n_3123),
.Y(n_3311)
);

BUFx3_ASAP7_75t_L g3312 ( 
.A(n_2916),
.Y(n_3312)
);

INVx3_ASAP7_75t_L g3313 ( 
.A(n_3104),
.Y(n_3313)
);

BUFx3_ASAP7_75t_L g3314 ( 
.A(n_3171),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_2764),
.B(n_592),
.Y(n_3315)
);

AND2x4_ASAP7_75t_L g3316 ( 
.A(n_2896),
.B(n_592),
.Y(n_3316)
);

AOI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_2988),
.A2(n_595),
.B1(n_593),
.B2(n_594),
.Y(n_3317)
);

BUFx6f_ASAP7_75t_L g3318 ( 
.A(n_3113),
.Y(n_3318)
);

AOI22xp33_ASAP7_75t_L g3319 ( 
.A1(n_2904),
.A2(n_3026),
.B1(n_3116),
.B2(n_3049),
.Y(n_3319)
);

INVx3_ASAP7_75t_L g3320 ( 
.A(n_3123),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_L g3321 ( 
.A(n_3006),
.B(n_595),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2881),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_2885),
.A2(n_595),
.B(n_596),
.Y(n_3323)
);

OR2x6_ASAP7_75t_L g3324 ( 
.A(n_2829),
.B(n_596),
.Y(n_3324)
);

INVx2_ASAP7_75t_SL g3325 ( 
.A(n_2909),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_2950),
.B(n_2821),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_2746),
.B(n_597),
.Y(n_3327)
);

AND2x2_ASAP7_75t_SL g3328 ( 
.A(n_2858),
.B(n_597),
.Y(n_3328)
);

A2O1A1Ixp33_ASAP7_75t_SL g3329 ( 
.A1(n_3001),
.A2(n_3073),
.B(n_3118),
.C(n_3003),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_3007),
.Y(n_3330)
);

INVx1_ASAP7_75t_SL g3331 ( 
.A(n_2954),
.Y(n_3331)
);

O2A1O1Ixp33_ASAP7_75t_L g3332 ( 
.A1(n_3169),
.A2(n_600),
.B(n_598),
.C(n_599),
.Y(n_3332)
);

CKINVDCx6p67_ASAP7_75t_R g3333 ( 
.A(n_2909),
.Y(n_3333)
);

BUFx12f_ASAP7_75t_L g3334 ( 
.A(n_2927),
.Y(n_3334)
);

INVx5_ASAP7_75t_L g3335 ( 
.A(n_2783),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_2887),
.Y(n_3336)
);

CKINVDCx16_ASAP7_75t_R g3337 ( 
.A(n_2927),
.Y(n_3337)
);

AOI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_2767),
.A2(n_600),
.B1(n_598),
.B2(n_599),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2761),
.Y(n_3339)
);

INVx3_ASAP7_75t_L g3340 ( 
.A(n_3130),
.Y(n_3340)
);

INVx4_ASAP7_75t_L g3341 ( 
.A(n_2862),
.Y(n_3341)
);

BUFx3_ASAP7_75t_L g3342 ( 
.A(n_3173),
.Y(n_3342)
);

INVx1_ASAP7_75t_SL g3343 ( 
.A(n_3130),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_2964),
.B(n_599),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2866),
.B(n_601),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_L g3346 ( 
.A1(n_3156),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_3346)
);

INVxp67_ASAP7_75t_SL g3347 ( 
.A(n_3170),
.Y(n_3347)
);

AOI22xp33_ASAP7_75t_L g3348 ( 
.A1(n_2850),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2752),
.B(n_2755),
.Y(n_3349)
);

NOR2xp67_ASAP7_75t_L g3350 ( 
.A(n_2921),
.B(n_602),
.Y(n_3350)
);

OAI321xp33_ASAP7_75t_L g3351 ( 
.A1(n_2770),
.A2(n_732),
.A3(n_730),
.B1(n_733),
.B2(n_731),
.C(n_729),
.Y(n_3351)
);

OAI22xp5_ASAP7_75t_L g3352 ( 
.A1(n_3018),
.A2(n_605),
.B1(n_603),
.B2(n_604),
.Y(n_3352)
);

NAND3xp33_ASAP7_75t_L g3353 ( 
.A(n_2774),
.B(n_605),
.C(n_606),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3170),
.B(n_606),
.Y(n_3354)
);

INVxp67_ASAP7_75t_SL g3355 ( 
.A(n_2783),
.Y(n_3355)
);

NOR2xp33_ASAP7_75t_L g3356 ( 
.A(n_2992),
.B(n_606),
.Y(n_3356)
);

OR2x2_ASAP7_75t_L g3357 ( 
.A(n_2993),
.B(n_607),
.Y(n_3357)
);

OAI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3018),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.Y(n_3358)
);

AND2x2_ASAP7_75t_L g3359 ( 
.A(n_3065),
.B(n_608),
.Y(n_3359)
);

NOR3xp33_ASAP7_75t_L g3360 ( 
.A(n_2820),
.B(n_609),
.C(n_610),
.Y(n_3360)
);

INVx3_ASAP7_75t_L g3361 ( 
.A(n_2858),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2762),
.Y(n_3362)
);

OR2x2_ASAP7_75t_L g3363 ( 
.A(n_2997),
.B(n_611),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_2905),
.Y(n_3364)
);

AOI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_2914),
.A2(n_613),
.B1(n_611),
.B2(n_612),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_2781),
.Y(n_3366)
);

NOR2xp33_ASAP7_75t_L g3367 ( 
.A(n_2999),
.B(n_611),
.Y(n_3367)
);

AOI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_2778),
.A2(n_612),
.B(n_613),
.Y(n_3368)
);

BUFx24_ASAP7_75t_SL g3369 ( 
.A(n_2785),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_2991),
.A2(n_615),
.B1(n_612),
.B2(n_614),
.Y(n_3370)
);

INVx5_ASAP7_75t_L g3371 ( 
.A(n_2786),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_3142),
.Y(n_3372)
);

NAND3xp33_ASAP7_75t_L g3373 ( 
.A(n_3153),
.B(n_614),
.C(n_615),
.Y(n_3373)
);

CKINVDCx8_ASAP7_75t_R g3374 ( 
.A(n_3129),
.Y(n_3374)
);

NAND3xp33_ASAP7_75t_L g3375 ( 
.A(n_3137),
.B(n_615),
.C(n_616),
.Y(n_3375)
);

AOI21xp5_ASAP7_75t_L g3376 ( 
.A1(n_2757),
.A2(n_616),
.B(n_617),
.Y(n_3376)
);

O2A1O1Ixp33_ASAP7_75t_L g3377 ( 
.A1(n_3046),
.A2(n_618),
.B(n_616),
.C(n_617),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_2749),
.B(n_617),
.Y(n_3378)
);

AND2x4_ASAP7_75t_L g3379 ( 
.A(n_3132),
.B(n_618),
.Y(n_3379)
);

BUFx12f_ASAP7_75t_L g3380 ( 
.A(n_3055),
.Y(n_3380)
);

AOI22xp33_ASAP7_75t_L g3381 ( 
.A1(n_3044),
.A2(n_3112),
.B1(n_3127),
.B2(n_3085),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_2959),
.Y(n_3382)
);

INVx2_ASAP7_75t_L g3383 ( 
.A(n_2960),
.Y(n_3383)
);

OR2x2_ASAP7_75t_SL g3384 ( 
.A(n_3150),
.B(n_619),
.Y(n_3384)
);

NOR2xp33_ASAP7_75t_L g3385 ( 
.A(n_2951),
.B(n_619),
.Y(n_3385)
);

BUFx3_ASAP7_75t_L g3386 ( 
.A(n_3142),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2795),
.Y(n_3387)
);

AOI21xp5_ASAP7_75t_L g3388 ( 
.A1(n_2948),
.A2(n_620),
.B(n_621),
.Y(n_3388)
);

NAND2x1p5_ASAP7_75t_L g3389 ( 
.A(n_2939),
.B(n_620),
.Y(n_3389)
);

AND2x4_ASAP7_75t_L g3390 ( 
.A(n_2852),
.B(n_621),
.Y(n_3390)
);

O2A1O1Ixp33_ASAP7_75t_L g3391 ( 
.A1(n_3099),
.A2(n_624),
.B(n_622),
.C(n_623),
.Y(n_3391)
);

AND2x4_ASAP7_75t_L g3392 ( 
.A(n_2994),
.B(n_622),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_2842),
.A2(n_2814),
.B1(n_3011),
.B2(n_2936),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2759),
.B(n_3013),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_3014),
.B(n_624),
.Y(n_3395)
);

INVx2_ASAP7_75t_SL g3396 ( 
.A(n_2962),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_L g3397 ( 
.A(n_2853),
.B(n_624),
.Y(n_3397)
);

BUFx2_ASAP7_75t_L g3398 ( 
.A(n_3101),
.Y(n_3398)
);

A2O1A1Ixp33_ASAP7_75t_L g3399 ( 
.A1(n_2800),
.A2(n_627),
.B(n_625),
.C(n_626),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3024),
.B(n_625),
.Y(n_3400)
);

AOI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_3021),
.A2(n_627),
.B1(n_625),
.B2(n_626),
.Y(n_3401)
);

INVx3_ASAP7_75t_L g3402 ( 
.A(n_2771),
.Y(n_3402)
);

AOI22xp5_ASAP7_75t_L g3403 ( 
.A1(n_3110),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3022),
.B(n_628),
.Y(n_3404)
);

CKINVDCx20_ASAP7_75t_R g3405 ( 
.A(n_3138),
.Y(n_3405)
);

AO21x2_ASAP7_75t_L g3406 ( 
.A1(n_2917),
.A2(n_629),
.B(n_630),
.Y(n_3406)
);

AND2x2_ASAP7_75t_L g3407 ( 
.A(n_2775),
.B(n_630),
.Y(n_3407)
);

CKINVDCx5p33_ASAP7_75t_R g3408 ( 
.A(n_3172),
.Y(n_3408)
);

NAND2x1p5_ASAP7_75t_L g3409 ( 
.A(n_2786),
.B(n_630),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2856),
.Y(n_3410)
);

O2A1O1Ixp33_ASAP7_75t_L g3411 ( 
.A1(n_3144),
.A2(n_3147),
.B(n_3155),
.C(n_3125),
.Y(n_3411)
);

OAI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_2835),
.A2(n_633),
.B1(n_631),
.B2(n_632),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_2891),
.Y(n_3413)
);

NOR2xp67_ASAP7_75t_L g3414 ( 
.A(n_2848),
.B(n_633),
.Y(n_3414)
);

BUFx2_ASAP7_75t_L g3415 ( 
.A(n_3101),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2877),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_2890),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_2802),
.B(n_634),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_2892),
.Y(n_3419)
);

INVx3_ASAP7_75t_L g3420 ( 
.A(n_3107),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3141),
.Y(n_3421)
);

CKINVDCx5p33_ASAP7_75t_R g3422 ( 
.A(n_2968),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3141),
.Y(n_3423)
);

AOI22xp5_ASAP7_75t_L g3424 ( 
.A1(n_3120),
.A2(n_636),
.B1(n_634),
.B2(n_635),
.Y(n_3424)
);

O2A1O1Ixp5_ASAP7_75t_SL g3425 ( 
.A1(n_2978),
.A2(n_733),
.B(n_734),
.C(n_732),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_2801),
.A2(n_637),
.B(n_635),
.C(n_636),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_2906),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3141),
.Y(n_3428)
);

O2A1O1Ixp33_ASAP7_75t_L g3429 ( 
.A1(n_3157),
.A2(n_2967),
.B(n_2969),
.C(n_2965),
.Y(n_3429)
);

INVx3_ASAP7_75t_L g3430 ( 
.A(n_2837),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2970),
.B(n_637),
.Y(n_3431)
);

BUFx3_ASAP7_75t_L g3432 ( 
.A(n_3151),
.Y(n_3432)
);

INVx3_ASAP7_75t_L g3433 ( 
.A(n_2837),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3160),
.Y(n_3434)
);

AND2x6_ASAP7_75t_L g3435 ( 
.A(n_2837),
.B(n_638),
.Y(n_3435)
);

OR2x6_ASAP7_75t_L g3436 ( 
.A(n_2773),
.B(n_639),
.Y(n_3436)
);

OAI22xp5_ASAP7_75t_L g3437 ( 
.A1(n_3045),
.A2(n_641),
.B1(n_639),
.B2(n_640),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_2883),
.Y(n_3438)
);

AND2x4_ASAP7_75t_L g3439 ( 
.A(n_2776),
.B(n_640),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3160),
.Y(n_3440)
);

BUFx3_ASAP7_75t_L g3441 ( 
.A(n_2883),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_3164),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2973),
.B(n_642),
.Y(n_3443)
);

AND2x4_ASAP7_75t_L g3444 ( 
.A(n_2776),
.B(n_643),
.Y(n_3444)
);

NAND2x1p5_ASAP7_75t_L g3445 ( 
.A(n_2883),
.B(n_643),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_2809),
.B(n_643),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3122),
.A2(n_646),
.B1(n_644),
.B2(n_645),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_2974),
.B(n_645),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3164),
.Y(n_3449)
);

OR2x2_ASAP7_75t_L g3450 ( 
.A(n_2817),
.B(n_645),
.Y(n_3450)
);

INVx2_ASAP7_75t_SL g3451 ( 
.A(n_3139),
.Y(n_3451)
);

OR2x2_ASAP7_75t_L g3452 ( 
.A(n_2823),
.B(n_646),
.Y(n_3452)
);

NAND2x1p5_ASAP7_75t_L g3453 ( 
.A(n_2900),
.B(n_646),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3164),
.Y(n_3454)
);

HB1xp67_ASAP7_75t_L g3455 ( 
.A(n_2826),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_2979),
.B(n_647),
.Y(n_3456)
);

CKINVDCx20_ASAP7_75t_R g3457 ( 
.A(n_3036),
.Y(n_3457)
);

AND2x4_ASAP7_75t_L g3458 ( 
.A(n_2844),
.B(n_648),
.Y(n_3458)
);

OR2x2_ASAP7_75t_L g3459 ( 
.A(n_2827),
.B(n_648),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_2931),
.Y(n_3460)
);

NAND3xp33_ASAP7_75t_L g3461 ( 
.A(n_2744),
.B(n_648),
.C(n_649),
.Y(n_3461)
);

INVx2_ASAP7_75t_SL g3462 ( 
.A(n_2900),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_2981),
.B(n_649),
.Y(n_3463)
);

AND2x4_ASAP7_75t_L g3464 ( 
.A(n_2846),
.B(n_649),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_2898),
.A2(n_652),
.B1(n_650),
.B2(n_651),
.Y(n_3465)
);

AOI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_2741),
.A2(n_650),
.B(n_651),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_2984),
.B(n_2985),
.Y(n_3467)
);

CKINVDCx5p33_ASAP7_75t_R g3468 ( 
.A(n_2840),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_2908),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_3469)
);

NOR2x1_ASAP7_75t_L g3470 ( 
.A(n_2955),
.B(n_654),
.Y(n_3470)
);

AND2x4_ASAP7_75t_L g3471 ( 
.A(n_2869),
.B(n_654),
.Y(n_3471)
);

AOI22xp5_ASAP7_75t_L g3472 ( 
.A1(n_3069),
.A2(n_657),
.B1(n_655),
.B2(n_656),
.Y(n_3472)
);

INVxp67_ASAP7_75t_L g3473 ( 
.A(n_2831),
.Y(n_3473)
);

BUFx2_ASAP7_75t_L g3474 ( 
.A(n_2900),
.Y(n_3474)
);

BUFx2_ASAP7_75t_R g3475 ( 
.A(n_3162),
.Y(n_3475)
);

OR2x6_ASAP7_75t_L g3476 ( 
.A(n_3145),
.B(n_656),
.Y(n_3476)
);

INVx2_ASAP7_75t_SL g3477 ( 
.A(n_2844),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_2832),
.B(n_657),
.Y(n_3478)
);

INVx3_ASAP7_75t_L g3479 ( 
.A(n_2882),
.Y(n_3479)
);

INVx3_ASAP7_75t_L g3480 ( 
.A(n_2882),
.Y(n_3480)
);

OAI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_2925),
.A2(n_659),
.B1(n_657),
.B2(n_658),
.Y(n_3481)
);

AND2x4_ASAP7_75t_L g3482 ( 
.A(n_2895),
.B(n_659),
.Y(n_3482)
);

NAND3xp33_ASAP7_75t_L g3483 ( 
.A(n_2915),
.B(n_2922),
.C(n_2815),
.Y(n_3483)
);

CKINVDCx8_ASAP7_75t_R g3484 ( 
.A(n_3070),
.Y(n_3484)
);

INVx3_ASAP7_75t_L g3485 ( 
.A(n_2886),
.Y(n_3485)
);

INVx3_ASAP7_75t_L g3486 ( 
.A(n_2886),
.Y(n_3486)
);

NOR2xp33_ASAP7_75t_L g3487 ( 
.A(n_2834),
.B(n_660),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_SL g3488 ( 
.A(n_2928),
.B(n_661),
.Y(n_3488)
);

INVx3_ASAP7_75t_L g3489 ( 
.A(n_2893),
.Y(n_3489)
);

OR2x6_ASAP7_75t_SL g3490 ( 
.A(n_3165),
.B(n_661),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3027),
.B(n_661),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_2972),
.Y(n_3492)
);

BUFx2_ASAP7_75t_L g3493 ( 
.A(n_2893),
.Y(n_3493)
);

AND2x4_ASAP7_75t_L g3494 ( 
.A(n_3111),
.B(n_662),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_L g3495 ( 
.A(n_3031),
.B(n_663),
.Y(n_3495)
);

NAND2x1p5_ASAP7_75t_L g3496 ( 
.A(n_2897),
.B(n_664),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_SL g3497 ( 
.A1(n_2818),
.A2(n_665),
.B(n_666),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3060),
.B(n_666),
.Y(n_3498)
);

INVx2_ASAP7_75t_SL g3499 ( 
.A(n_2897),
.Y(n_3499)
);

OAI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3030),
.A2(n_3032),
.B1(n_2947),
.B2(n_2957),
.Y(n_3500)
);

BUFx2_ASAP7_75t_L g3501 ( 
.A(n_2901),
.Y(n_3501)
);

CKINVDCx20_ASAP7_75t_R g3502 ( 
.A(n_2889),
.Y(n_3502)
);

BUFx6f_ASAP7_75t_L g3503 ( 
.A(n_2901),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3042),
.B(n_667),
.Y(n_3504)
);

AND2x6_ASAP7_75t_L g3505 ( 
.A(n_2938),
.B(n_667),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3015),
.B(n_668),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3043),
.B(n_668),
.Y(n_3507)
);

INVx3_ASAP7_75t_L g3508 ( 
.A(n_2938),
.Y(n_3508)
);

OAI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3166),
.A2(n_672),
.B1(n_670),
.B2(n_671),
.Y(n_3509)
);

O2A1O1Ixp5_ASAP7_75t_L g3510 ( 
.A1(n_2841),
.A2(n_673),
.B(n_671),
.C(n_672),
.Y(n_3510)
);

CKINVDCx20_ASAP7_75t_R g3511 ( 
.A(n_3072),
.Y(n_3511)
);

O2A1O1Ixp33_ASAP7_75t_SL g3512 ( 
.A1(n_3146),
.A2(n_674),
.B(n_672),
.C(n_673),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3075),
.B(n_673),
.Y(n_3513)
);

AND2x2_ASAP7_75t_L g3514 ( 
.A(n_3077),
.B(n_675),
.Y(n_3514)
);

CKINVDCx11_ASAP7_75t_R g3515 ( 
.A(n_3154),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3078),
.B(n_675),
.Y(n_3516)
);

AO21x2_ASAP7_75t_L g3517 ( 
.A1(n_2920),
.A2(n_675),
.B(n_676),
.Y(n_3517)
);

INVx5_ASAP7_75t_L g3518 ( 
.A(n_3008),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3081),
.B(n_676),
.Y(n_3519)
);

INVxp67_ASAP7_75t_L g3520 ( 
.A(n_3082),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3089),
.B(n_3090),
.Y(n_3521)
);

CKINVDCx20_ASAP7_75t_R g3522 ( 
.A(n_3092),
.Y(n_3522)
);

AND2x2_ASAP7_75t_L g3523 ( 
.A(n_3098),
.B(n_677),
.Y(n_3523)
);

NAND2xp5_ASAP7_75t_L g3524 ( 
.A(n_3088),
.B(n_677),
.Y(n_3524)
);

BUFx12f_ASAP7_75t_L g3525 ( 
.A(n_3056),
.Y(n_3525)
);

NOR2x1_ASAP7_75t_L g3526 ( 
.A(n_3052),
.B(n_679),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_3100),
.B(n_3057),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_2782),
.B(n_679),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_2791),
.B(n_680),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_3008),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2792),
.B(n_680),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2794),
.B(n_680),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_3016),
.Y(n_3533)
);

AND2x2_ASAP7_75t_SL g3534 ( 
.A(n_3158),
.B(n_681),
.Y(n_3534)
);

INVx4_ASAP7_75t_SL g3535 ( 
.A(n_2937),
.Y(n_3535)
);

AOI22xp5_ASAP7_75t_L g3536 ( 
.A1(n_3168),
.A2(n_684),
.B1(n_681),
.B2(n_683),
.Y(n_3536)
);

BUFx2_ASAP7_75t_L g3537 ( 
.A(n_3016),
.Y(n_3537)
);

OAI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3063),
.A2(n_684),
.B1(n_681),
.B2(n_683),
.Y(n_3538)
);

O2A1O1Ixp33_ASAP7_75t_L g3539 ( 
.A1(n_3134),
.A2(n_685),
.B(n_683),
.C(n_684),
.Y(n_3539)
);

OAI22xp5_ASAP7_75t_L g3540 ( 
.A1(n_3066),
.A2(n_688),
.B1(n_686),
.B2(n_687),
.Y(n_3540)
);

INVx2_ASAP7_75t_SL g3541 ( 
.A(n_3086),
.Y(n_3541)
);

INVx1_ASAP7_75t_L g3542 ( 
.A(n_2937),
.Y(n_3542)
);

O2A1O1Ixp5_ASAP7_75t_SL g3543 ( 
.A1(n_2934),
.A2(n_736),
.B(n_737),
.C(n_735),
.Y(n_3543)
);

BUFx6f_ASAP7_75t_L g3544 ( 
.A(n_3086),
.Y(n_3544)
);

INVxp67_ASAP7_75t_L g3545 ( 
.A(n_2983),
.Y(n_3545)
);

BUFx3_ASAP7_75t_L g3546 ( 
.A(n_3096),
.Y(n_3546)
);

AND2x4_ASAP7_75t_L g3547 ( 
.A(n_3096),
.B(n_686),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_L g3548 ( 
.A1(n_2753),
.A2(n_687),
.B(n_688),
.Y(n_3548)
);

INVx4_ASAP7_75t_L g3549 ( 
.A(n_3121),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_2803),
.B(n_687),
.Y(n_3550)
);

BUFx12f_ASAP7_75t_L g3551 ( 
.A(n_2982),
.Y(n_3551)
);

BUFx3_ASAP7_75t_L g3552 ( 
.A(n_3163),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3102),
.B(n_691),
.Y(n_3553)
);

BUFx6f_ASAP7_75t_L g3554 ( 
.A(n_2758),
.Y(n_3554)
);

BUFx12f_ASAP7_75t_L g3555 ( 
.A(n_2912),
.Y(n_3555)
);

INVx1_ASAP7_75t_SL g3556 ( 
.A(n_2806),
.Y(n_3556)
);

AND2x4_ASAP7_75t_L g3557 ( 
.A(n_3103),
.B(n_691),
.Y(n_3557)
);

AOI22x1_ASAP7_75t_L g3558 ( 
.A1(n_2779),
.A2(n_694),
.B1(n_692),
.B2(n_693),
.Y(n_3558)
);

OAI22xp5_ASAP7_75t_L g3559 ( 
.A1(n_3161),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.Y(n_3559)
);

INVx5_ASAP7_75t_L g3560 ( 
.A(n_2793),
.Y(n_3560)
);

AND2x4_ASAP7_75t_L g3561 ( 
.A(n_3167),
.B(n_696),
.Y(n_3561)
);

BUFx2_ASAP7_75t_L g3562 ( 
.A(n_2784),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3109),
.B(n_697),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_2819),
.B(n_697),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_2825),
.B(n_698),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_2790),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3028),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_2859),
.B(n_698),
.Y(n_3568)
);

O2A1O1Ixp33_ASAP7_75t_SL g3569 ( 
.A1(n_3152),
.A2(n_701),
.B(n_699),
.C(n_700),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3047),
.Y(n_3570)
);

AND2x6_ASAP7_75t_L g3571 ( 
.A(n_3117),
.B(n_699),
.Y(n_3571)
);

INVx5_ASAP7_75t_L g3572 ( 
.A(n_3039),
.Y(n_3572)
);

AND2x4_ASAP7_75t_L g3573 ( 
.A(n_3124),
.B(n_699),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_2871),
.B(n_700),
.Y(n_3574)
);

AOI21xp5_ASAP7_75t_L g3575 ( 
.A1(n_2763),
.A2(n_702),
.B(n_703),
.Y(n_3575)
);

AOI22xp33_ASAP7_75t_SL g3576 ( 
.A1(n_2812),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_3576)
);

INVx3_ASAP7_75t_L g3577 ( 
.A(n_3083),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3048),
.Y(n_3578)
);

INVx4_ASAP7_75t_L g3579 ( 
.A(n_3076),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3054),
.Y(n_3580)
);

AND2x2_ASAP7_75t_L g3581 ( 
.A(n_2874),
.B(n_702),
.Y(n_3581)
);

HB1xp67_ASAP7_75t_L g3582 ( 
.A(n_2854),
.Y(n_3582)
);

INVx1_ASAP7_75t_SL g3583 ( 
.A(n_2879),
.Y(n_3583)
);

OR2x2_ASAP7_75t_SL g3584 ( 
.A(n_2961),
.B(n_703),
.Y(n_3584)
);

AO32x2_ASAP7_75t_L g3585 ( 
.A1(n_2907),
.A2(n_706),
.A3(n_704),
.B1(n_705),
.B2(n_707),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_2796),
.Y(n_3586)
);

AND2x2_ASAP7_75t_L g3587 ( 
.A(n_2888),
.B(n_706),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_2894),
.B(n_706),
.Y(n_3588)
);

NAND2xp33_ASAP7_75t_L g3589 ( 
.A(n_3159),
.B(n_708),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_2918),
.B(n_708),
.Y(n_3590)
);

AND2x4_ASAP7_75t_L g3591 ( 
.A(n_3091),
.B(n_736),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3093),
.Y(n_3592)
);

AND2x4_ASAP7_75t_L g3593 ( 
.A(n_2903),
.B(n_738),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_2930),
.A2(n_743),
.B1(n_739),
.B2(n_742),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_2941),
.B(n_2944),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_2805),
.Y(n_3596)
);

INVx8_ASAP7_75t_L g3597 ( 
.A(n_2926),
.Y(n_3597)
);

BUFx2_ASAP7_75t_L g3598 ( 
.A(n_3136),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_3105),
.Y(n_3599)
);

INVx2_ASAP7_75t_L g3600 ( 
.A(n_3108),
.Y(n_3600)
);

AND2x4_ASAP7_75t_L g3601 ( 
.A(n_2986),
.B(n_978),
.Y(n_3601)
);

OR2x6_ASAP7_75t_L g3602 ( 
.A(n_2958),
.B(n_746),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3023),
.B(n_2976),
.Y(n_3603)
);

INVxp67_ASAP7_75t_L g3604 ( 
.A(n_2998),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3002),
.B(n_977),
.Y(n_3605)
);

INVx2_ASAP7_75t_SL g3606 ( 
.A(n_2961),
.Y(n_3606)
);

BUFx3_ASAP7_75t_L g3607 ( 
.A(n_2863),
.Y(n_3607)
);

INVx5_ASAP7_75t_L g3608 ( 
.A(n_3068),
.Y(n_3608)
);

AND2x6_ASAP7_75t_L g3609 ( 
.A(n_3136),
.B(n_3106),
.Y(n_3609)
);

BUFx2_ASAP7_75t_L g3610 ( 
.A(n_3136),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3012),
.B(n_977),
.Y(n_3611)
);

BUFx4f_ASAP7_75t_L g3612 ( 
.A(n_3219),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3179),
.Y(n_3613)
);

CKINVDCx20_ASAP7_75t_R g3614 ( 
.A(n_3201),
.Y(n_3614)
);

BUFx2_ASAP7_75t_L g3615 ( 
.A(n_3333),
.Y(n_3615)
);

INVx1_ASAP7_75t_SL g3616 ( 
.A(n_3221),
.Y(n_3616)
);

HB1xp67_ASAP7_75t_L g3617 ( 
.A(n_3200),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3181),
.Y(n_3618)
);

BUFx2_ASAP7_75t_L g3619 ( 
.A(n_3405),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3207),
.Y(n_3620)
);

BUFx2_ASAP7_75t_R g3621 ( 
.A(n_3232),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3227),
.B(n_3114),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_SL g3623 ( 
.A1(n_3195),
.A2(n_3228),
.B(n_3174),
.Y(n_3623)
);

AOI22xp5_ASAP7_75t_L g3624 ( 
.A1(n_3328),
.A2(n_2780),
.B1(n_3053),
.B2(n_3051),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3597),
.A2(n_3071),
.B1(n_3074),
.B2(n_3067),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3217),
.Y(n_3626)
);

BUFx2_ASAP7_75t_R g3627 ( 
.A(n_3192),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3252),
.Y(n_3628)
);

OAI22xp33_ASAP7_75t_L g3629 ( 
.A1(n_3337),
.A2(n_3080),
.B1(n_3115),
.B2(n_3079),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3224),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3248),
.Y(n_3631)
);

BUFx6f_ASAP7_75t_L g3632 ( 
.A(n_3261),
.Y(n_3632)
);

AOI22xp5_ASAP7_75t_SL g3633 ( 
.A1(n_3270),
.A2(n_3135),
.B1(n_3140),
.B2(n_3119),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3250),
.Y(n_3634)
);

BUFx6f_ASAP7_75t_L g3635 ( 
.A(n_3261),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3251),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3259),
.Y(n_3637)
);

BUFx2_ASAP7_75t_L g3638 ( 
.A(n_3334),
.Y(n_3638)
);

HB1xp67_ASAP7_75t_L g3639 ( 
.A(n_3331),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3293),
.Y(n_3640)
);

CKINVDCx16_ASAP7_75t_R g3641 ( 
.A(n_3188),
.Y(n_3641)
);

INVx4_ASAP7_75t_L g3642 ( 
.A(n_3262),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3225),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3191),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3196),
.Y(n_3645)
);

CKINVDCx11_ASAP7_75t_R g3646 ( 
.A(n_3243),
.Y(n_3646)
);

HB1xp67_ASAP7_75t_L g3647 ( 
.A(n_3311),
.Y(n_3647)
);

AND2x4_ASAP7_75t_L g3648 ( 
.A(n_3262),
.B(n_2961),
.Y(n_3648)
);

NAND2x1p5_ASAP7_75t_L g3649 ( 
.A(n_3246),
.B(n_3133),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3205),
.Y(n_3650)
);

AO21x2_ASAP7_75t_L g3651 ( 
.A1(n_3204),
.A2(n_3586),
.B(n_3566),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3263),
.B(n_752),
.Y(n_3652)
);

INVx4_ASAP7_75t_SL g3653 ( 
.A(n_3435),
.Y(n_3653)
);

INVx2_ASAP7_75t_L g3654 ( 
.A(n_3281),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3283),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_3475),
.B(n_753),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3326),
.B(n_3339),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3322),
.Y(n_3658)
);

INVx1_ASAP7_75t_SL g3659 ( 
.A(n_3296),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3231),
.Y(n_3660)
);

AOI22xp5_ASAP7_75t_L g3661 ( 
.A1(n_3457),
.A2(n_3422),
.B1(n_3414),
.B2(n_3277),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3233),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3336),
.Y(n_3663)
);

NAND2x1p5_ASAP7_75t_L g3664 ( 
.A(n_3216),
.B(n_754),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3364),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3382),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3383),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3396),
.Y(n_3668)
);

AOI21x1_ASAP7_75t_L g3669 ( 
.A1(n_3185),
.A2(n_2884),
.B(n_2907),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3379),
.Y(n_3670)
);

BUFx2_ASAP7_75t_R g3671 ( 
.A(n_3212),
.Y(n_3671)
);

BUFx2_ASAP7_75t_L g3672 ( 
.A(n_3432),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3362),
.B(n_2989),
.Y(n_3673)
);

OA21x2_ASAP7_75t_L g3674 ( 
.A1(n_3203),
.A2(n_2884),
.B(n_2989),
.Y(n_3674)
);

BUFx2_ASAP7_75t_R g3675 ( 
.A(n_3308),
.Y(n_3675)
);

HB1xp67_ASAP7_75t_L g3676 ( 
.A(n_3305),
.Y(n_3676)
);

INVx11_ASAP7_75t_L g3677 ( 
.A(n_3298),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3379),
.Y(n_3678)
);

AO21x2_ASAP7_75t_L g3679 ( 
.A1(n_3596),
.A2(n_3025),
.B(n_3020),
.Y(n_3679)
);

INVx2_ASAP7_75t_SL g3680 ( 
.A(n_3206),
.Y(n_3680)
);

NAND2x1_ASAP7_75t_L g3681 ( 
.A(n_3228),
.B(n_3025),
.Y(n_3681)
);

OAI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3384),
.A2(n_3184),
.B1(n_3324),
.B2(n_3534),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3297),
.Y(n_3683)
);

BUFx3_ASAP7_75t_L g3684 ( 
.A(n_3206),
.Y(n_3684)
);

BUFx2_ASAP7_75t_R g3685 ( 
.A(n_3240),
.Y(n_3685)
);

BUFx4f_ASAP7_75t_L g3686 ( 
.A(n_3229),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3366),
.B(n_3033),
.Y(n_3687)
);

INVx4_ASAP7_75t_L g3688 ( 
.A(n_3262),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3591),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3591),
.Y(n_3690)
);

CKINVDCx5p33_ASAP7_75t_R g3691 ( 
.A(n_3237),
.Y(n_3691)
);

HB1xp67_ASAP7_75t_L g3692 ( 
.A(n_3309),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3381),
.A2(n_759),
.B1(n_755),
.B2(n_757),
.Y(n_3693)
);

OAI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3272),
.A2(n_755),
.B(n_760),
.Y(n_3694)
);

OAI22xp33_ASAP7_75t_L g3695 ( 
.A1(n_3256),
.A2(n_3324),
.B1(n_3451),
.B2(n_3350),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3304),
.Y(n_3696)
);

CKINVDCx5p33_ASAP7_75t_R g3697 ( 
.A(n_3260),
.Y(n_3697)
);

INVx1_ASAP7_75t_L g3698 ( 
.A(n_3387),
.Y(n_3698)
);

AOI22xp5_ASAP7_75t_L g3699 ( 
.A1(n_3256),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_SL g3700 ( 
.A(n_3341),
.B(n_3244),
.Y(n_3700)
);

CKINVDCx14_ASAP7_75t_R g3701 ( 
.A(n_3223),
.Y(n_3701)
);

NAND2x1_ASAP7_75t_L g3702 ( 
.A(n_3562),
.B(n_3609),
.Y(n_3702)
);

AOI22xp5_ASAP7_75t_L g3703 ( 
.A1(n_3467),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3319),
.B(n_3455),
.Y(n_3704)
);

INVx3_ASAP7_75t_L g3705 ( 
.A(n_3288),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3359),
.Y(n_3706)
);

CKINVDCx6p67_ASAP7_75t_R g3707 ( 
.A(n_3274),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3307),
.Y(n_3708)
);

INVx1_ASAP7_75t_L g3709 ( 
.A(n_3330),
.Y(n_3709)
);

INVx3_ASAP7_75t_L g3710 ( 
.A(n_3213),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3400),
.Y(n_3711)
);

OA21x2_ASAP7_75t_L g3712 ( 
.A1(n_3542),
.A2(n_766),
.B(n_767),
.Y(n_3712)
);

BUFx6f_ASAP7_75t_L g3713 ( 
.A(n_3318),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3410),
.B(n_768),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3354),
.Y(n_3715)
);

BUFx6f_ASAP7_75t_L g3716 ( 
.A(n_3318),
.Y(n_3716)
);

CKINVDCx5p33_ASAP7_75t_R g3717 ( 
.A(n_3226),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3269),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3394),
.Y(n_3719)
);

CKINVDCx5p33_ASAP7_75t_R g3720 ( 
.A(n_3211),
.Y(n_3720)
);

AOI22xp33_ASAP7_75t_SL g3721 ( 
.A1(n_3402),
.A2(n_772),
.B1(n_770),
.B2(n_771),
.Y(n_3721)
);

INVx4_ASAP7_75t_L g3722 ( 
.A(n_3220),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3416),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3417),
.Y(n_3724)
);

AND2x2_ASAP7_75t_L g3725 ( 
.A(n_3178),
.B(n_976),
.Y(n_3725)
);

OR2x2_ASAP7_75t_L g3726 ( 
.A(n_3289),
.B(n_774),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3419),
.Y(n_3727)
);

INVx1_ASAP7_75t_L g3728 ( 
.A(n_3439),
.Y(n_3728)
);

BUFx2_ASAP7_75t_SL g3729 ( 
.A(n_3435),
.Y(n_3729)
);

BUFx2_ASAP7_75t_L g3730 ( 
.A(n_3222),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3439),
.Y(n_3731)
);

INVxp67_ASAP7_75t_L g3732 ( 
.A(n_3314),
.Y(n_3732)
);

AO21x1_ASAP7_75t_SL g3733 ( 
.A1(n_3460),
.A2(n_775),
.B(n_776),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3444),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3444),
.Y(n_3735)
);

INVx2_ASAP7_75t_L g3736 ( 
.A(n_3458),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_L g3737 ( 
.A1(n_3561),
.A2(n_780),
.B1(n_777),
.B2(n_778),
.Y(n_3737)
);

HB1xp67_ASAP7_75t_L g3738 ( 
.A(n_3343),
.Y(n_3738)
);

AO21x1_ASAP7_75t_L g3739 ( 
.A1(n_3352),
.A2(n_778),
.B(n_780),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3458),
.Y(n_3740)
);

OR2x2_ASAP7_75t_L g3741 ( 
.A(n_3398),
.B(n_781),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3547),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3547),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3247),
.Y(n_3744)
);

BUFx2_ASAP7_75t_L g3745 ( 
.A(n_3264),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3194),
.B(n_781),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_3342),
.Y(n_3747)
);

AOI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3397),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3585),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3584),
.Y(n_3750)
);

AOI22xp33_ASAP7_75t_SL g3751 ( 
.A1(n_3435),
.A2(n_786),
.B1(n_784),
.B2(n_785),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3585),
.Y(n_3752)
);

INVx3_ASAP7_75t_L g3753 ( 
.A(n_3335),
.Y(n_3753)
);

BUFx6f_ASAP7_75t_L g3754 ( 
.A(n_3515),
.Y(n_3754)
);

NAND2xp5_ASAP7_75t_L g3755 ( 
.A(n_3177),
.B(n_788),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3585),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3253),
.Y(n_3757)
);

BUFx12f_ASAP7_75t_L g3758 ( 
.A(n_3210),
.Y(n_3758)
);

CKINVDCx6p67_ASAP7_75t_R g3759 ( 
.A(n_3197),
.Y(n_3759)
);

AOI22xp33_ASAP7_75t_L g3760 ( 
.A1(n_3593),
.A2(n_790),
.B1(n_788),
.B2(n_789),
.Y(n_3760)
);

INVx2_ASAP7_75t_SL g3761 ( 
.A(n_3299),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3373),
.Y(n_3762)
);

HB1xp67_ASAP7_75t_SL g3763 ( 
.A(n_3374),
.Y(n_3763)
);

BUFx3_ASAP7_75t_L g3764 ( 
.A(n_3299),
.Y(n_3764)
);

INVx2_ASAP7_75t_SL g3765 ( 
.A(n_3302),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3392),
.Y(n_3766)
);

AOI22xp33_ASAP7_75t_L g3767 ( 
.A1(n_3601),
.A2(n_791),
.B1(n_789),
.B2(n_790),
.Y(n_3767)
);

AND2x4_ASAP7_75t_L g3768 ( 
.A(n_3398),
.B(n_791),
.Y(n_3768)
);

HB1xp67_ASAP7_75t_L g3769 ( 
.A(n_3284),
.Y(n_3769)
);

INVx2_ASAP7_75t_SL g3770 ( 
.A(n_3303),
.Y(n_3770)
);

HB1xp67_ASAP7_75t_L g3771 ( 
.A(n_3325),
.Y(n_3771)
);

OAI22xp5_ASAP7_75t_L g3772 ( 
.A1(n_3182),
.A2(n_794),
.B1(n_792),
.B2(n_793),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3258),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_L g3774 ( 
.A1(n_3500),
.A2(n_794),
.B1(n_792),
.B2(n_793),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3517),
.Y(n_3775)
);

CKINVDCx20_ASAP7_75t_R g3776 ( 
.A(n_3511),
.Y(n_3776)
);

BUFx2_ASAP7_75t_SL g3777 ( 
.A(n_3264),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3189),
.B(n_795),
.Y(n_3778)
);

AOI22xp33_ASAP7_75t_L g3779 ( 
.A1(n_3608),
.A2(n_3573),
.B1(n_3557),
.B2(n_3464),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3199),
.B(n_795),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3441),
.Y(n_3781)
);

AOI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_3608),
.A2(n_3360),
.B1(n_3234),
.B2(n_3602),
.Y(n_3782)
);

BUFx6f_ASAP7_75t_L g3783 ( 
.A(n_3239),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3473),
.B(n_796),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3599),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3600),
.Y(n_3786)
);

HB1xp67_ASAP7_75t_L g3787 ( 
.A(n_3347),
.Y(n_3787)
);

INVx3_ASAP7_75t_L g3788 ( 
.A(n_3386),
.Y(n_3788)
);

AOI22xp33_ASAP7_75t_SL g3789 ( 
.A1(n_3415),
.A2(n_800),
.B1(n_798),
.B2(n_799),
.Y(n_3789)
);

AOI22xp33_ASAP7_75t_L g3790 ( 
.A1(n_3608),
.A2(n_801),
.B1(n_798),
.B2(n_800),
.Y(n_3790)
);

AOI22xp33_ASAP7_75t_L g3791 ( 
.A1(n_3602),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3268),
.Y(n_3792)
);

INVx3_ASAP7_75t_L g3793 ( 
.A(n_3335),
.Y(n_3793)
);

NAND2x1p5_ASAP7_75t_L g3794 ( 
.A(n_3239),
.B(n_802),
.Y(n_3794)
);

AND2x2_ASAP7_75t_L g3795 ( 
.A(n_3275),
.B(n_3241),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3280),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_L g3797 ( 
.A(n_3254),
.Y(n_3797)
);

BUFx6f_ASAP7_75t_L g3798 ( 
.A(n_3254),
.Y(n_3798)
);

AND2x4_ASAP7_75t_L g3799 ( 
.A(n_3415),
.B(n_803),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_3183),
.B(n_804),
.Y(n_3800)
);

AO21x1_ASAP7_75t_SL g3801 ( 
.A1(n_3492),
.A2(n_805),
.B(n_806),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3285),
.Y(n_3802)
);

AOI22xp33_ASAP7_75t_L g3803 ( 
.A1(n_3589),
.A2(n_3218),
.B1(n_3407),
.B2(n_3393),
.Y(n_3803)
);

INVx1_ASAP7_75t_L g3804 ( 
.A(n_3286),
.Y(n_3804)
);

HB1xp67_ASAP7_75t_L g3805 ( 
.A(n_3320),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3292),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3505),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3553),
.A2(n_811),
.B1(n_808),
.B2(n_810),
.Y(n_3808)
);

INVx6_ASAP7_75t_L g3809 ( 
.A(n_3380),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3335),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3371),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3505),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3371),
.Y(n_3813)
);

AOI22xp33_ASAP7_75t_SL g3814 ( 
.A1(n_3408),
.A2(n_817),
.B1(n_815),
.B2(n_816),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3563),
.A2(n_818),
.B1(n_815),
.B2(n_817),
.Y(n_3815)
);

AOI22xp33_ASAP7_75t_L g3816 ( 
.A1(n_3238),
.A2(n_3209),
.B1(n_3476),
.B2(n_3436),
.Y(n_3816)
);

OAI21x1_ASAP7_75t_L g3817 ( 
.A1(n_3577),
.A2(n_818),
.B(n_821),
.Y(n_3817)
);

HB1xp67_ASAP7_75t_L g3818 ( 
.A(n_3340),
.Y(n_3818)
);

BUFx2_ASAP7_75t_L g3819 ( 
.A(n_3313),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3505),
.Y(n_3820)
);

OR2x2_ASAP7_75t_L g3821 ( 
.A(n_3344),
.B(n_821),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3421),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3423),
.Y(n_3823)
);

AOI22xp33_ASAP7_75t_L g3824 ( 
.A1(n_3238),
.A2(n_824),
.B1(n_822),
.B2(n_823),
.Y(n_3824)
);

CKINVDCx20_ASAP7_75t_R g3825 ( 
.A(n_3522),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3371),
.Y(n_3826)
);

HB1xp67_ASAP7_75t_L g3827 ( 
.A(n_3493),
.Y(n_3827)
);

CKINVDCx6p67_ASAP7_75t_R g3828 ( 
.A(n_3312),
.Y(n_3828)
);

AND2x2_ASAP7_75t_L g3829 ( 
.A(n_3316),
.B(n_825),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3503),
.Y(n_3830)
);

NAND2x1_ASAP7_75t_L g3831 ( 
.A(n_3609),
.B(n_826),
.Y(n_3831)
);

NAND2x1p5_ASAP7_75t_L g3832 ( 
.A(n_3372),
.B(n_827),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3503),
.Y(n_3833)
);

AOI22xp33_ASAP7_75t_L g3834 ( 
.A1(n_3436),
.A2(n_3476),
.B1(n_3187),
.B2(n_3526),
.Y(n_3834)
);

INVx8_ASAP7_75t_L g3835 ( 
.A(n_3208),
.Y(n_3835)
);

BUFx10_ASAP7_75t_L g3836 ( 
.A(n_3390),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3428),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3434),
.Y(n_3838)
);

INVx4_ASAP7_75t_L g3839 ( 
.A(n_3291),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3544),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3440),
.Y(n_3841)
);

OAI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_3273),
.A2(n_830),
.B1(n_828),
.B2(n_829),
.Y(n_3842)
);

HB1xp67_ASAP7_75t_L g3843 ( 
.A(n_3493),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3442),
.Y(n_3844)
);

INVx2_ASAP7_75t_L g3845 ( 
.A(n_3544),
.Y(n_3845)
);

OAI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_3490),
.A2(n_831),
.B1(n_828),
.B2(n_830),
.Y(n_3846)
);

AOI22xp33_ASAP7_75t_L g3847 ( 
.A1(n_3193),
.A2(n_833),
.B1(n_831),
.B2(n_832),
.Y(n_3847)
);

BUFx12f_ASAP7_75t_L g3848 ( 
.A(n_3214),
.Y(n_3848)
);

CKINVDCx11_ASAP7_75t_R g3849 ( 
.A(n_3502),
.Y(n_3849)
);

AOI22xp33_ASAP7_75t_L g3850 ( 
.A1(n_3249),
.A2(n_835),
.B1(n_832),
.B2(n_834),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3449),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3462),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3454),
.Y(n_3853)
);

INVx4_ASAP7_75t_L g3854 ( 
.A(n_3306),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3430),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3433),
.Y(n_3856)
);

BUFx2_ASAP7_75t_L g3857 ( 
.A(n_3549),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3349),
.B(n_837),
.Y(n_3858)
);

AND2x4_ASAP7_75t_L g3859 ( 
.A(n_3501),
.B(n_837),
.Y(n_3859)
);

HB1xp67_ASAP7_75t_L g3860 ( 
.A(n_3501),
.Y(n_3860)
);

BUFx6f_ASAP7_75t_L g3861 ( 
.A(n_3438),
.Y(n_3861)
);

AND2x2_ASAP7_75t_L g3862 ( 
.A(n_3378),
.B(n_838),
.Y(n_3862)
);

CKINVDCx6p67_ASAP7_75t_R g3863 ( 
.A(n_3471),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3438),
.Y(n_3864)
);

BUFx2_ASAP7_75t_L g3865 ( 
.A(n_3530),
.Y(n_3865)
);

BUFx3_ASAP7_75t_L g3866 ( 
.A(n_3546),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3406),
.Y(n_3867)
);

HB1xp67_ASAP7_75t_L g3868 ( 
.A(n_3537),
.Y(n_3868)
);

HB1xp67_ASAP7_75t_L g3869 ( 
.A(n_3537),
.Y(n_3869)
);

INVx1_ASAP7_75t_L g3870 ( 
.A(n_3446),
.Y(n_3870)
);

HB1xp67_ASAP7_75t_L g3871 ( 
.A(n_3361),
.Y(n_3871)
);

OAI22xp5_ASAP7_75t_L g3872 ( 
.A1(n_3265),
.A2(n_840),
.B1(n_838),
.B2(n_839),
.Y(n_3872)
);

HB1xp67_ASAP7_75t_L g3873 ( 
.A(n_3474),
.Y(n_3873)
);

BUFx8_ASAP7_75t_L g3874 ( 
.A(n_3482),
.Y(n_3874)
);

NOR2xp33_ASAP7_75t_L g3875 ( 
.A(n_3301),
.B(n_839),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3450),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3474),
.Y(n_3877)
);

AOI22xp33_ASAP7_75t_SL g3878 ( 
.A1(n_3560),
.A2(n_843),
.B1(n_840),
.B2(n_841),
.Y(n_3878)
);

HB1xp67_ASAP7_75t_L g3879 ( 
.A(n_3477),
.Y(n_3879)
);

INVx3_ASAP7_75t_L g3880 ( 
.A(n_3420),
.Y(n_3880)
);

NAND2x1p5_ASAP7_75t_L g3881 ( 
.A(n_3518),
.B(n_844),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_3287),
.B(n_845),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3567),
.Y(n_3883)
);

BUFx2_ASAP7_75t_L g3884 ( 
.A(n_3355),
.Y(n_3884)
);

INVx2_ASAP7_75t_L g3885 ( 
.A(n_3570),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3452),
.Y(n_3886)
);

INVx8_ASAP7_75t_L g3887 ( 
.A(n_3518),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3459),
.Y(n_3888)
);

INVx3_ASAP7_75t_L g3889 ( 
.A(n_3496),
.Y(n_3889)
);

INVx2_ASAP7_75t_SL g3890 ( 
.A(n_3389),
.Y(n_3890)
);

OR2x6_ASAP7_75t_L g3891 ( 
.A(n_3271),
.B(n_845),
.Y(n_3891)
);

INVx3_ASAP7_75t_L g3892 ( 
.A(n_3186),
.Y(n_3892)
);

BUFx2_ASAP7_75t_SL g3893 ( 
.A(n_3560),
.Y(n_3893)
);

AOI22xp5_ASAP7_75t_L g3894 ( 
.A1(n_3180),
.A2(n_848),
.B1(n_846),
.B2(n_847),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3375),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3357),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3578),
.Y(n_3897)
);

INVx6_ASAP7_75t_L g3898 ( 
.A(n_3255),
.Y(n_3898)
);

AOI22xp33_ASAP7_75t_L g3899 ( 
.A1(n_3465),
.A2(n_850),
.B1(n_848),
.B2(n_849),
.Y(n_3899)
);

AOI22xp33_ASAP7_75t_L g3900 ( 
.A1(n_3488),
.A2(n_853),
.B1(n_851),
.B2(n_852),
.Y(n_3900)
);

CKINVDCx20_ASAP7_75t_R g3901 ( 
.A(n_3468),
.Y(n_3901)
);

BUFx3_ASAP7_75t_L g3902 ( 
.A(n_3479),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_L g3903 ( 
.A(n_3520),
.B(n_854),
.Y(n_3903)
);

BUFx2_ASAP7_75t_L g3904 ( 
.A(n_3480),
.Y(n_3904)
);

AND2x2_ASAP7_75t_L g3905 ( 
.A(n_3418),
.B(n_857),
.Y(n_3905)
);

INVx3_ASAP7_75t_L g3906 ( 
.A(n_3186),
.Y(n_3906)
);

OAI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3346),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_3363),
.Y(n_3908)
);

INVx2_ASAP7_75t_SL g3909 ( 
.A(n_3485),
.Y(n_3909)
);

HB1xp67_ASAP7_75t_L g3910 ( 
.A(n_3499),
.Y(n_3910)
);

INVx4_ASAP7_75t_L g3911 ( 
.A(n_3560),
.Y(n_3911)
);

AOI22xp33_ASAP7_75t_SL g3912 ( 
.A1(n_3525),
.A2(n_860),
.B1(n_858),
.B2(n_859),
.Y(n_3912)
);

INVx1_ASAP7_75t_L g3913 ( 
.A(n_3215),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3385),
.B(n_860),
.Y(n_3914)
);

INVx2_ASAP7_75t_SL g3915 ( 
.A(n_3486),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3551),
.Y(n_3916)
);

INVx2_ASAP7_75t_L g3917 ( 
.A(n_3580),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3592),
.Y(n_3918)
);

OAI22xp5_ASAP7_75t_L g3919 ( 
.A1(n_3469),
.A2(n_863),
.B1(n_861),
.B2(n_862),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3555),
.Y(n_3920)
);

AOI22xp33_ASAP7_75t_L g3921 ( 
.A1(n_3463),
.A2(n_863),
.B1(n_861),
.B2(n_862),
.Y(n_3921)
);

BUFx5_ASAP7_75t_L g3922 ( 
.A(n_3571),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3484),
.Y(n_3923)
);

INVx3_ASAP7_75t_L g3924 ( 
.A(n_3489),
.Y(n_3924)
);

BUFx2_ASAP7_75t_L g3925 ( 
.A(n_3508),
.Y(n_3925)
);

BUFx6f_ASAP7_75t_L g3926 ( 
.A(n_3190),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3606),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_L g3928 ( 
.A(n_3395),
.B(n_866),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3514),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3516),
.B(n_866),
.Y(n_3930)
);

INVx3_ASAP7_75t_L g3931 ( 
.A(n_3552),
.Y(n_3931)
);

HB1xp67_ASAP7_75t_L g3932 ( 
.A(n_3541),
.Y(n_3932)
);

INVx2_ASAP7_75t_L g3933 ( 
.A(n_3574),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3519),
.B(n_867),
.Y(n_3934)
);

INVx1_ASAP7_75t_SL g3935 ( 
.A(n_3523),
.Y(n_3935)
);

INVx2_ASAP7_75t_SL g3936 ( 
.A(n_3533),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3491),
.Y(n_3937)
);

AO21x1_ASAP7_75t_L g3938 ( 
.A1(n_3358),
.A2(n_868),
.B(n_869),
.Y(n_3938)
);

OR2x6_ASAP7_75t_L g3939 ( 
.A(n_3276),
.B(n_869),
.Y(n_3939)
);

AOI22xp33_ASAP7_75t_L g3940 ( 
.A1(n_3267),
.A2(n_872),
.B1(n_870),
.B2(n_871),
.Y(n_3940)
);

INVx1_ASAP7_75t_L g3941 ( 
.A(n_3495),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3504),
.Y(n_3942)
);

BUFx6f_ASAP7_75t_L g3943 ( 
.A(n_3190),
.Y(n_3943)
);

OR2x2_ASAP7_75t_L g3944 ( 
.A(n_3279),
.B(n_870),
.Y(n_3944)
);

CKINVDCx11_ASAP7_75t_R g3945 ( 
.A(n_3494),
.Y(n_3945)
);

CKINVDCx11_ASAP7_75t_R g3946 ( 
.A(n_3556),
.Y(n_3946)
);

CKINVDCx20_ASAP7_75t_R g3947 ( 
.A(n_3290),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3581),
.Y(n_3948)
);

BUFx2_ASAP7_75t_L g3949 ( 
.A(n_3409),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3587),
.Y(n_3950)
);

AOI22xp33_ASAP7_75t_L g3951 ( 
.A1(n_3483),
.A2(n_873),
.B1(n_871),
.B2(n_872),
.Y(n_3951)
);

INVx11_ASAP7_75t_L g3952 ( 
.A(n_3571),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3590),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3535),
.Y(n_3954)
);

BUFx8_ASAP7_75t_L g3955 ( 
.A(n_3198),
.Y(n_3955)
);

BUFx2_ASAP7_75t_R g3956 ( 
.A(n_3294),
.Y(n_3956)
);

BUFx2_ASAP7_75t_R g3957 ( 
.A(n_3521),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3506),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3356),
.B(n_873),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3437),
.A2(n_3235),
.B1(n_3245),
.B2(n_3559),
.Y(n_3960)
);

BUFx2_ASAP7_75t_R g3961 ( 
.A(n_3513),
.Y(n_3961)
);

AOI21xp33_ASAP7_75t_L g3962 ( 
.A1(n_3329),
.A2(n_3411),
.B(n_3230),
.Y(n_3962)
);

BUFx6f_ASAP7_75t_L g3963 ( 
.A(n_3198),
.Y(n_3963)
);

INVx3_ASAP7_75t_L g3964 ( 
.A(n_3445),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3321),
.B(n_976),
.Y(n_3965)
);

INVx3_ASAP7_75t_L g3966 ( 
.A(n_3453),
.Y(n_3966)
);

NAND2x1p5_ASAP7_75t_L g3967 ( 
.A(n_3470),
.B(n_874),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3367),
.B(n_874),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3535),
.Y(n_3969)
);

INVx3_ASAP7_75t_L g3970 ( 
.A(n_3571),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3413),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3478),
.B(n_975),
.Y(n_3972)
);

NAND2x1p5_ASAP7_75t_L g3973 ( 
.A(n_3338),
.B(n_875),
.Y(n_3973)
);

BUFx10_ASAP7_75t_L g3974 ( 
.A(n_3202),
.Y(n_3974)
);

AND2x2_ASAP7_75t_L g3975 ( 
.A(n_3487),
.B(n_3295),
.Y(n_3975)
);

AND2x2_ASAP7_75t_L g3976 ( 
.A(n_3327),
.B(n_975),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3427),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3507),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3524),
.Y(n_3979)
);

INVx2_ASAP7_75t_SL g3980 ( 
.A(n_3257),
.Y(n_3980)
);

BUFx10_ASAP7_75t_L g3981 ( 
.A(n_3315),
.Y(n_3981)
);

BUFx3_ASAP7_75t_L g3982 ( 
.A(n_3528),
.Y(n_3982)
);

CKINVDCx20_ASAP7_75t_R g3983 ( 
.A(n_3536),
.Y(n_3983)
);

CKINVDCx20_ASAP7_75t_R g3984 ( 
.A(n_3300),
.Y(n_3984)
);

BUFx4f_ASAP7_75t_L g3985 ( 
.A(n_3527),
.Y(n_3985)
);

AOI22xp5_ASAP7_75t_L g3986 ( 
.A1(n_3176),
.A2(n_3369),
.B1(n_3365),
.B2(n_3236),
.Y(n_3986)
);

CKINVDCx11_ASAP7_75t_R g3987 ( 
.A(n_3583),
.Y(n_3987)
);

OAI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_3510),
.A2(n_875),
.B(n_876),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3431),
.B(n_3443),
.Y(n_3989)
);

BUFx2_ASAP7_75t_L g3990 ( 
.A(n_3607),
.Y(n_3990)
);

AOI22xp33_ASAP7_75t_L g3991 ( 
.A1(n_3538),
.A2(n_878),
.B1(n_876),
.B2(n_877),
.Y(n_3991)
);

AND2x4_ASAP7_75t_L g3992 ( 
.A(n_3598),
.B(n_3610),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3448),
.Y(n_3993)
);

INVx11_ASAP7_75t_L g3994 ( 
.A(n_3609),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3628),
.Y(n_3995)
);

INVx2_ASAP7_75t_L g3996 ( 
.A(n_3654),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3613),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3795),
.B(n_3598),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3655),
.Y(n_3999)
);

OR2x6_ASAP7_75t_L g4000 ( 
.A(n_3729),
.B(n_3282),
.Y(n_4000)
);

INVx2_ASAP7_75t_L g4001 ( 
.A(n_3658),
.Y(n_4001)
);

BUFx4f_ASAP7_75t_L g4002 ( 
.A(n_3754),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3618),
.Y(n_4003)
);

BUFx3_ASAP7_75t_L g4004 ( 
.A(n_3809),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3620),
.Y(n_4005)
);

NAND3x1_ASAP7_75t_L g4006 ( 
.A(n_3661),
.B(n_3317),
.C(n_3403),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3626),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3630),
.Y(n_4008)
);

INVx1_ASAP7_75t_L g4009 ( 
.A(n_3631),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3634),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3822),
.Y(n_4011)
);

INVx2_ASAP7_75t_SL g4012 ( 
.A(n_3809),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3823),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3837),
.Y(n_4014)
);

INVx2_ASAP7_75t_L g4015 ( 
.A(n_3665),
.Y(n_4015)
);

HB1xp67_ASAP7_75t_L g4016 ( 
.A(n_3639),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3838),
.Y(n_4017)
);

AND2x4_ASAP7_75t_L g4018 ( 
.A(n_3653),
.B(n_3610),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3841),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3644),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3796),
.B(n_3545),
.Y(n_4021)
);

INVx1_ASAP7_75t_L g4022 ( 
.A(n_3844),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3645),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3636),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3650),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3637),
.Y(n_4026)
);

OAI211xp5_ASAP7_75t_L g4027 ( 
.A1(n_3816),
.A2(n_3472),
.B(n_3424),
.C(n_3401),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3640),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3723),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3660),
.Y(n_4030)
);

OR2x2_ASAP7_75t_L g4031 ( 
.A(n_3617),
.B(n_3456),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3724),
.Y(n_4032)
);

INVx3_ASAP7_75t_L g4033 ( 
.A(n_3722),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3662),
.Y(n_4034)
);

INVx1_ASAP7_75t_SL g4035 ( 
.A(n_3828),
.Y(n_4035)
);

AND2x2_ASAP7_75t_L g4036 ( 
.A(n_3802),
.B(n_3804),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3727),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3663),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3698),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3643),
.Y(n_4040)
);

INVx3_ASAP7_75t_L g4041 ( 
.A(n_3722),
.Y(n_4041)
);

AND2x4_ASAP7_75t_L g4042 ( 
.A(n_3653),
.B(n_3572),
.Y(n_4042)
);

BUFx3_ASAP7_75t_L g4043 ( 
.A(n_3747),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_L g4044 ( 
.A(n_3719),
.B(n_3704),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3806),
.B(n_3604),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3683),
.Y(n_4046)
);

OAI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_3962),
.A2(n_3543),
.B(n_3351),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3696),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3666),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3667),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_3708),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3709),
.Y(n_4052)
);

INVx3_ASAP7_75t_L g4053 ( 
.A(n_3848),
.Y(n_4053)
);

OR2x6_ASAP7_75t_L g4054 ( 
.A(n_3729),
.B(n_3497),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_3884),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3647),
.Y(n_4056)
);

BUFx12f_ASAP7_75t_L g4057 ( 
.A(n_3646),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3948),
.B(n_3404),
.Y(n_4058)
);

HB1xp67_ASAP7_75t_L g4059 ( 
.A(n_3787),
.Y(n_4059)
);

BUFx2_ASAP7_75t_L g4060 ( 
.A(n_3745),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3676),
.Y(n_4061)
);

BUFx2_ASAP7_75t_L g4062 ( 
.A(n_3990),
.Y(n_4062)
);

INVx3_ASAP7_75t_L g4063 ( 
.A(n_3686),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3692),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3689),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3690),
.Y(n_4066)
);

BUFx2_ASAP7_75t_L g4067 ( 
.A(n_3827),
.Y(n_4067)
);

HB1xp67_ASAP7_75t_L g4068 ( 
.A(n_3843),
.Y(n_4068)
);

BUFx2_ASAP7_75t_SL g4069 ( 
.A(n_3839),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3769),
.Y(n_4070)
);

HB1xp67_ASAP7_75t_L g4071 ( 
.A(n_3860),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3668),
.Y(n_4072)
);

OR2x6_ASAP7_75t_L g4073 ( 
.A(n_3835),
.B(n_3323),
.Y(n_4073)
);

OAI21x1_ASAP7_75t_L g4074 ( 
.A1(n_3669),
.A2(n_3278),
.B(n_3425),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_3738),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3785),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_3715),
.B(n_3582),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3786),
.Y(n_4078)
);

BUFx3_ASAP7_75t_L g4079 ( 
.A(n_3754),
.Y(n_4079)
);

AOI22xp33_ASAP7_75t_SL g4080 ( 
.A1(n_3682),
.A2(n_3572),
.B1(n_3540),
.B2(n_3370),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_3935),
.B(n_3579),
.Y(n_4081)
);

BUFx6f_ASAP7_75t_L g4082 ( 
.A(n_3632),
.Y(n_4082)
);

NAND2x1p5_ASAP7_75t_L g4083 ( 
.A(n_3612),
.B(n_3558),
.Y(n_4083)
);

AND2x4_ASAP7_75t_L g4084 ( 
.A(n_3992),
.B(n_3572),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3864),
.Y(n_4085)
);

INVx2_ASAP7_75t_SL g4086 ( 
.A(n_3754),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3730),
.Y(n_4087)
);

OAI22xp5_ASAP7_75t_L g4088 ( 
.A1(n_3779),
.A2(n_3426),
.B1(n_3399),
.B2(n_3310),
.Y(n_4088)
);

BUFx2_ASAP7_75t_L g4089 ( 
.A(n_3868),
.Y(n_4089)
);

HB1xp67_ASAP7_75t_L g4090 ( 
.A(n_3869),
.Y(n_4090)
);

NAND2x1p5_ASAP7_75t_L g4091 ( 
.A(n_3638),
.B(n_3594),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3851),
.Y(n_4092)
);

AO21x1_ASAP7_75t_SL g4093 ( 
.A1(n_3782),
.A2(n_3595),
.B(n_3603),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3853),
.Y(n_4094)
);

HB1xp67_ASAP7_75t_L g4095 ( 
.A(n_3672),
.Y(n_4095)
);

BUFx2_ASAP7_75t_L g4096 ( 
.A(n_3955),
.Y(n_4096)
);

OR2x6_ASAP7_75t_L g4097 ( 
.A(n_3835),
.B(n_3377),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3657),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3744),
.Y(n_4099)
);

OR2x2_ASAP7_75t_L g4100 ( 
.A(n_3933),
.B(n_3950),
.Y(n_4100)
);

INVx2_ASAP7_75t_L g4101 ( 
.A(n_3877),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3757),
.Y(n_4102)
);

BUFx3_ASAP7_75t_L g4103 ( 
.A(n_3684),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3913),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_3652),
.B(n_3554),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_L g4106 ( 
.A(n_3857),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3670),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3870),
.B(n_3429),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3678),
.Y(n_4109)
);

INVx4_ASAP7_75t_L g4110 ( 
.A(n_3887),
.Y(n_4110)
);

AND2x4_ASAP7_75t_L g4111 ( 
.A(n_3992),
.B(n_3353),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3876),
.Y(n_4112)
);

OR2x6_ASAP7_75t_L g4113 ( 
.A(n_3893),
.B(n_3368),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_3725),
.B(n_3576),
.Y(n_4114)
);

NOR2xp33_ASAP7_75t_L g4115 ( 
.A(n_3616),
.B(n_3498),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3886),
.B(n_3345),
.Y(n_4116)
);

AND2x2_ASAP7_75t_L g4117 ( 
.A(n_3929),
.B(n_878),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3888),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_3771),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3883),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3879),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3896),
.B(n_3509),
.Y(n_4122)
);

INVx1_ASAP7_75t_L g4123 ( 
.A(n_3910),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_3908),
.B(n_879),
.Y(n_4124)
);

INVx2_ASAP7_75t_L g4125 ( 
.A(n_3885),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_3706),
.B(n_879),
.Y(n_4126)
);

INVx2_ASAP7_75t_L g4127 ( 
.A(n_3897),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3932),
.Y(n_4128)
);

INVx1_ASAP7_75t_L g4129 ( 
.A(n_3871),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3805),
.Y(n_4130)
);

INVx3_ASAP7_75t_L g4131 ( 
.A(n_3641),
.Y(n_4131)
);

HB1xp67_ASAP7_75t_L g4132 ( 
.A(n_3873),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_3818),
.Y(n_4133)
);

INVx5_ASAP7_75t_L g4134 ( 
.A(n_3887),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_3953),
.B(n_880),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3766),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3979),
.B(n_3481),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_3773),
.B(n_3175),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_3777),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3917),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_3865),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_3918),
.Y(n_4142)
);

BUFx3_ASAP7_75t_L g4143 ( 
.A(n_3720),
.Y(n_4143)
);

OR2x6_ASAP7_75t_L g4144 ( 
.A(n_3893),
.B(n_3388),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_3792),
.B(n_3266),
.Y(n_4145)
);

INVx3_ASAP7_75t_L g4146 ( 
.A(n_3866),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3777),
.Y(n_4147)
);

HB1xp67_ASAP7_75t_L g4148 ( 
.A(n_3819),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_3741),
.Y(n_4149)
);

HB1xp67_ASAP7_75t_L g4150 ( 
.A(n_3859),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3615),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3711),
.B(n_3348),
.Y(n_4152)
);

HB1xp67_ASAP7_75t_L g4153 ( 
.A(n_3859),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_3861),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_3985),
.B(n_3980),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3993),
.Y(n_4156)
);

HB1xp67_ASAP7_75t_L g4157 ( 
.A(n_3904),
.Y(n_4157)
);

CKINVDCx20_ASAP7_75t_R g4158 ( 
.A(n_3614),
.Y(n_4158)
);

HB1xp67_ASAP7_75t_L g4159 ( 
.A(n_3925),
.Y(n_4159)
);

BUFx2_ASAP7_75t_L g4160 ( 
.A(n_3955),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3673),
.Y(n_4161)
);

HB1xp67_ASAP7_75t_L g4162 ( 
.A(n_3861),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3687),
.Y(n_4163)
);

NAND2xp5_ASAP7_75t_L g4164 ( 
.A(n_3718),
.B(n_3391),
.Y(n_4164)
);

AND2x2_ASAP7_75t_L g4165 ( 
.A(n_3750),
.B(n_880),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_3905),
.B(n_881),
.Y(n_4166)
);

INVx2_ASAP7_75t_SL g4167 ( 
.A(n_3764),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_3862),
.B(n_882),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3937),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_3941),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3942),
.Y(n_4171)
);

CKINVDCx16_ASAP7_75t_R g4172 ( 
.A(n_3763),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_3728),
.B(n_882),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3958),
.Y(n_4174)
);

BUFx3_ASAP7_75t_L g4175 ( 
.A(n_3619),
.Y(n_4175)
);

BUFx3_ASAP7_75t_L g4176 ( 
.A(n_3758),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_3861),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3978),
.Y(n_4178)
);

INVx2_ASAP7_75t_SL g4179 ( 
.A(n_3680),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3731),
.B(n_883),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3867),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3734),
.Y(n_4182)
);

INVx1_ASAP7_75t_L g4183 ( 
.A(n_3735),
.Y(n_4183)
);

OR2x6_ASAP7_75t_L g4184 ( 
.A(n_3768),
.B(n_3376),
.Y(n_4184)
);

BUFx2_ASAP7_75t_L g4185 ( 
.A(n_3926),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3740),
.Y(n_4186)
);

NOR2xp33_ASAP7_75t_L g4187 ( 
.A(n_3732),
.B(n_3945),
.Y(n_4187)
);

INVx2_ASAP7_75t_L g4188 ( 
.A(n_3852),
.Y(n_4188)
);

HB1xp67_ASAP7_75t_L g4189 ( 
.A(n_3982),
.Y(n_4189)
);

INVx2_ASAP7_75t_L g4190 ( 
.A(n_3651),
.Y(n_4190)
);

AND2x2_ASAP7_75t_L g4191 ( 
.A(n_3742),
.B(n_883),
.Y(n_4191)
);

AND2x4_ASAP7_75t_L g4192 ( 
.A(n_3926),
.B(n_3461),
.Y(n_4192)
);

BUFx3_ASAP7_75t_L g4193 ( 
.A(n_3717),
.Y(n_4193)
);

AND2x2_ASAP7_75t_L g4194 ( 
.A(n_3743),
.B(n_884),
.Y(n_4194)
);

INVx5_ASAP7_75t_SL g4195 ( 
.A(n_3677),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_3807),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_3821),
.B(n_3529),
.Y(n_4197)
);

OR2x6_ASAP7_75t_L g4198 ( 
.A(n_3768),
.B(n_3332),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_3812),
.Y(n_4199)
);

OAI21x1_ASAP7_75t_L g4200 ( 
.A1(n_3831),
.A2(n_3702),
.B(n_3775),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_3820),
.Y(n_4201)
);

OR2x6_ASAP7_75t_L g4202 ( 
.A(n_3799),
.B(n_3466),
.Y(n_4202)
);

HB1xp67_ASAP7_75t_L g4203 ( 
.A(n_3931),
.Y(n_4203)
);

BUFx3_ASAP7_75t_L g4204 ( 
.A(n_3707),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3749),
.Y(n_4205)
);

AOI222xp33_ASAP7_75t_L g4206 ( 
.A1(n_3695),
.A2(n_3412),
.B1(n_3550),
.B2(n_3588),
.C1(n_3532),
.C2(n_3568),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_3736),
.B(n_3930),
.Y(n_4207)
);

BUFx2_ASAP7_75t_L g4208 ( 
.A(n_3926),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_3989),
.B(n_3781),
.Y(n_4209)
);

OR2x2_ASAP7_75t_L g4210 ( 
.A(n_3726),
.B(n_3531),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3752),
.Y(n_4211)
);

INVx1_ASAP7_75t_SL g4212 ( 
.A(n_3849),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3756),
.Y(n_4213)
);

OAI21xp33_ASAP7_75t_SL g4214 ( 
.A1(n_3952),
.A2(n_3447),
.B(n_3605),
.Y(n_4214)
);

NOR2xp67_ASAP7_75t_SL g4215 ( 
.A(n_3970),
.B(n_3611),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3714),
.Y(n_4216)
);

AND2x2_ASAP7_75t_L g4217 ( 
.A(n_3863),
.B(n_884),
.Y(n_4217)
);

INVx2_ASAP7_75t_SL g4218 ( 
.A(n_3635),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3799),
.Y(n_4219)
);

BUFx2_ASAP7_75t_L g4220 ( 
.A(n_3943),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3931),
.Y(n_4221)
);

BUFx3_ASAP7_75t_L g4222 ( 
.A(n_3788),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3710),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_3829),
.B(n_885),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3855),
.Y(n_4225)
);

HB1xp67_ASAP7_75t_L g4226 ( 
.A(n_3810),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3784),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_3856),
.Y(n_4228)
);

INVx2_ASAP7_75t_SL g4229 ( 
.A(n_3713),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3712),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3712),
.Y(n_4231)
);

HB1xp67_ASAP7_75t_L g4232 ( 
.A(n_3811),
.Y(n_4232)
);

CKINVDCx5p33_ASAP7_75t_R g4233 ( 
.A(n_3621),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_3997),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_4003),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4055),
.Y(n_4236)
);

AND2x4_ASAP7_75t_L g4237 ( 
.A(n_4062),
.B(n_3954),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4011),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4011),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4013),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_3995),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_4013),
.Y(n_4242)
);

AND2x4_ASAP7_75t_L g4243 ( 
.A(n_4062),
.B(n_3969),
.Y(n_4243)
);

AND2x2_ASAP7_75t_L g4244 ( 
.A(n_3998),
.B(n_3974),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4014),
.Y(n_4245)
);

OR2x2_ASAP7_75t_L g4246 ( 
.A(n_4059),
.B(n_3623),
.Y(n_4246)
);

AND2x2_ASAP7_75t_L g4247 ( 
.A(n_4209),
.B(n_3974),
.Y(n_4247)
);

HB1xp67_ASAP7_75t_L g4248 ( 
.A(n_4106),
.Y(n_4248)
);

AND2x4_ASAP7_75t_L g4249 ( 
.A(n_4060),
.B(n_3648),
.Y(n_4249)
);

AND2x2_ASAP7_75t_L g4250 ( 
.A(n_4226),
.B(n_3943),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_4232),
.B(n_3943),
.Y(n_4251)
);

BUFx3_ASAP7_75t_L g4252 ( 
.A(n_4043),
.Y(n_4252)
);

BUFx3_ASAP7_75t_L g4253 ( 
.A(n_4004),
.Y(n_4253)
);

BUFx3_ASAP7_75t_L g4254 ( 
.A(n_4096),
.Y(n_4254)
);

INVx2_ASAP7_75t_L g4255 ( 
.A(n_3996),
.Y(n_4255)
);

BUFx3_ASAP7_75t_L g4256 ( 
.A(n_4096),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_4189),
.B(n_3963),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_4005),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_3999),
.Y(n_4259)
);

AND2x2_ASAP7_75t_L g4260 ( 
.A(n_4105),
.B(n_3963),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4007),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4008),
.Y(n_4262)
);

HB1xp67_ASAP7_75t_L g4263 ( 
.A(n_4060),
.Y(n_4263)
);

INVx2_ASAP7_75t_L g4264 ( 
.A(n_4001),
.Y(n_4264)
);

OR2x2_ASAP7_75t_L g4265 ( 
.A(n_4056),
.B(n_3963),
.Y(n_4265)
);

AND2x2_ASAP7_75t_L g4266 ( 
.A(n_4095),
.B(n_3648),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4015),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4148),
.B(n_3946),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4098),
.B(n_3803),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4009),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_4044),
.B(n_4112),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4010),
.Y(n_4272)
);

HB1xp67_ASAP7_75t_L g4273 ( 
.A(n_4068),
.Y(n_4273)
);

HB1xp67_ASAP7_75t_L g4274 ( 
.A(n_4071),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_4141),
.B(n_4075),
.Y(n_4275)
);

BUFx2_ASAP7_75t_L g4276 ( 
.A(n_4160),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4024),
.Y(n_4277)
);

INVx2_ASAP7_75t_L g4278 ( 
.A(n_4020),
.Y(n_4278)
);

INVx2_ASAP7_75t_L g4279 ( 
.A(n_4023),
.Y(n_4279)
);

INVx2_ASAP7_75t_L g4280 ( 
.A(n_4025),
.Y(n_4280)
);

OR2x2_ASAP7_75t_L g4281 ( 
.A(n_4061),
.B(n_3927),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4026),
.Y(n_4282)
);

OR2x2_ASAP7_75t_L g4283 ( 
.A(n_4064),
.B(n_3759),
.Y(n_4283)
);

AND2x4_ASAP7_75t_SL g4284 ( 
.A(n_4110),
.B(n_3901),
.Y(n_4284)
);

BUFx2_ASAP7_75t_L g4285 ( 
.A(n_4160),
.Y(n_4285)
);

INVx2_ASAP7_75t_L g4286 ( 
.A(n_4030),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_4118),
.B(n_3986),
.Y(n_4287)
);

OR2x2_ASAP7_75t_L g4288 ( 
.A(n_4090),
.B(n_3679),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4028),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4121),
.B(n_3987),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4029),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4014),
.Y(n_4292)
);

HB1xp67_ASAP7_75t_L g4293 ( 
.A(n_4132),
.Y(n_4293)
);

BUFx6f_ASAP7_75t_L g4294 ( 
.A(n_4134),
.Y(n_4294)
);

BUFx2_ASAP7_75t_L g4295 ( 
.A(n_4033),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4032),
.Y(n_4296)
);

INVx2_ASAP7_75t_SL g4297 ( 
.A(n_4134),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_4017),
.Y(n_4298)
);

HB1xp67_ASAP7_75t_L g4299 ( 
.A(n_4067),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4017),
.Y(n_4300)
);

BUFx2_ASAP7_75t_L g4301 ( 
.A(n_4041),
.Y(n_4301)
);

INVx2_ASAP7_75t_L g4302 ( 
.A(n_4034),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_4019),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4038),
.Y(n_4304)
);

HB1xp67_ASAP7_75t_L g4305 ( 
.A(n_4067),
.Y(n_4305)
);

AND2x2_ASAP7_75t_L g4306 ( 
.A(n_4123),
.B(n_3892),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_4128),
.B(n_3906),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_4156),
.B(n_3834),
.Y(n_4308)
);

AND2x2_ASAP7_75t_L g4309 ( 
.A(n_4119),
.B(n_3761),
.Y(n_4309)
);

OR2x2_ASAP7_75t_L g4310 ( 
.A(n_4100),
.B(n_4016),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4037),
.Y(n_4311)
);

AOI221xp5_ASAP7_75t_L g4312 ( 
.A1(n_4108),
.A2(n_3846),
.B1(n_3622),
.B2(n_3875),
.C(n_3842),
.Y(n_4312)
);

INVx2_ASAP7_75t_L g4313 ( 
.A(n_4049),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4169),
.B(n_3746),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_4050),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4207),
.B(n_3981),
.Y(n_4316)
);

NOR2x1_ASAP7_75t_L g4317 ( 
.A(n_4069),
.B(n_3911),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_4170),
.B(n_3674),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_4171),
.B(n_3674),
.Y(n_4319)
);

HB1xp67_ASAP7_75t_L g4320 ( 
.A(n_4089),
.Y(n_4320)
);

HB1xp67_ASAP7_75t_L g4321 ( 
.A(n_4089),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_4110),
.Y(n_4322)
);

AND2x2_ASAP7_75t_L g4323 ( 
.A(n_4081),
.B(n_3981),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_4039),
.Y(n_4324)
);

INVx2_ASAP7_75t_L g4325 ( 
.A(n_4076),
.Y(n_4325)
);

AND2x2_ASAP7_75t_L g4326 ( 
.A(n_4070),
.B(n_3898),
.Y(n_4326)
);

AND2x4_ASAP7_75t_L g4327 ( 
.A(n_4018),
.B(n_3702),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4174),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_4078),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4085),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_4019),
.Y(n_4331)
);

BUFx6f_ASAP7_75t_L g4332 ( 
.A(n_4134),
.Y(n_4332)
);

INVx2_ASAP7_75t_SL g4333 ( 
.A(n_4143),
.Y(n_4333)
);

NOR2x1_ASAP7_75t_SL g4334 ( 
.A(n_4069),
.B(n_3733),
.Y(n_4334)
);

AND2x2_ASAP7_75t_L g4335 ( 
.A(n_4087),
.B(n_3898),
.Y(n_4335)
);

OR2x2_ASAP7_75t_L g4336 ( 
.A(n_4157),
.B(n_3681),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4178),
.Y(n_4337)
);

HB1xp67_ASAP7_75t_L g4338 ( 
.A(n_4159),
.Y(n_4338)
);

NOR2x1_ASAP7_75t_SL g4339 ( 
.A(n_4054),
.B(n_3801),
.Y(n_4339)
);

INVx1_ASAP7_75t_SL g4340 ( 
.A(n_4103),
.Y(n_4340)
);

INVx2_ASAP7_75t_SL g4341 ( 
.A(n_4002),
.Y(n_4341)
);

BUFx2_ASAP7_75t_L g4342 ( 
.A(n_4203),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_4031),
.B(n_3681),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4101),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4036),
.B(n_3836),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4040),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_4021),
.B(n_3836),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4129),
.B(n_3830),
.Y(n_4348)
);

BUFx2_ASAP7_75t_L g4349 ( 
.A(n_4146),
.Y(n_4349)
);

AND2x2_ASAP7_75t_L g4350 ( 
.A(n_4130),
.B(n_3833),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4046),
.Y(n_4351)
);

INVx4_ASAP7_75t_SL g4352 ( 
.A(n_4204),
.Y(n_4352)
);

HB1xp67_ASAP7_75t_L g4353 ( 
.A(n_4188),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4048),
.Y(n_4354)
);

OR2x2_ASAP7_75t_L g4355 ( 
.A(n_4133),
.B(n_3971),
.Y(n_4355)
);

OR2x2_ASAP7_75t_L g4356 ( 
.A(n_4072),
.B(n_4161),
.Y(n_4356)
);

AND2x2_ASAP7_75t_L g4357 ( 
.A(n_4045),
.B(n_3840),
.Y(n_4357)
);

OR2x2_ASAP7_75t_L g4358 ( 
.A(n_4163),
.B(n_3977),
.Y(n_4358)
);

NOR2xp33_ASAP7_75t_L g4359 ( 
.A(n_4212),
.B(n_3675),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4022),
.Y(n_4360)
);

HB1xp67_ASAP7_75t_L g4361 ( 
.A(n_4150),
.Y(n_4361)
);

NAND2x1p5_ASAP7_75t_L g4362 ( 
.A(n_4053),
.B(n_3839),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4153),
.B(n_3845),
.Y(n_4363)
);

HB1xp67_ASAP7_75t_L g4364 ( 
.A(n_4162),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4120),
.Y(n_4365)
);

NAND2xp5_ASAP7_75t_L g4366 ( 
.A(n_4099),
.B(n_4102),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4125),
.Y(n_4367)
);

AND2x4_ASAP7_75t_L g4368 ( 
.A(n_4327),
.B(n_4018),
.Y(n_4368)
);

NAND3xp33_ASAP7_75t_L g4369 ( 
.A(n_4312),
.B(n_4115),
.C(n_4080),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_4273),
.B(n_4136),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_L g4371 ( 
.A(n_4274),
.B(n_4104),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4266),
.B(n_4175),
.Y(n_4372)
);

OAI22xp5_ASAP7_75t_L g4373 ( 
.A1(n_4276),
.A2(n_4097),
.B1(n_4198),
.B2(n_4073),
.Y(n_4373)
);

OAI22xp5_ASAP7_75t_L g4374 ( 
.A1(n_4285),
.A2(n_4097),
.B1(n_4198),
.B2(n_4073),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_4293),
.B(n_4182),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4260),
.B(n_4155),
.Y(n_4376)
);

AND2x2_ASAP7_75t_L g4377 ( 
.A(n_4244),
.B(n_4077),
.Y(n_4377)
);

NOR2xp33_ASAP7_75t_L g4378 ( 
.A(n_4359),
.B(n_4079),
.Y(n_4378)
);

NAND3xp33_ASAP7_75t_L g4379 ( 
.A(n_4299),
.B(n_4227),
.C(n_4047),
.Y(n_4379)
);

NAND3xp33_ASAP7_75t_L g4380 ( 
.A(n_4305),
.B(n_4214),
.C(n_4199),
.Y(n_4380)
);

AOI22xp33_ASAP7_75t_SL g4381 ( 
.A1(n_4339),
.A2(n_3874),
.B1(n_4219),
.B2(n_4217),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4338),
.B(n_4196),
.Y(n_4382)
);

OAI221xp5_ASAP7_75t_SL g4383 ( 
.A1(n_4246),
.A2(n_4202),
.B1(n_4184),
.B2(n_4027),
.C(n_4206),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4287),
.B(n_4183),
.Y(n_4384)
);

OAI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_4322),
.A2(n_4256),
.B1(n_4254),
.B2(n_4317),
.Y(n_4385)
);

OAI221xp5_ASAP7_75t_L g4386 ( 
.A1(n_4269),
.A2(n_4091),
.B1(n_3814),
.B2(n_3656),
.C(n_4083),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_4361),
.B(n_4186),
.Y(n_4387)
);

NAND3xp33_ASAP7_75t_L g4388 ( 
.A(n_4320),
.B(n_4201),
.C(n_4216),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_4271),
.B(n_4107),
.Y(n_4389)
);

INVx1_ASAP7_75t_L g4390 ( 
.A(n_4234),
.Y(n_4390)
);

AND2x2_ASAP7_75t_L g4391 ( 
.A(n_4248),
.B(n_4185),
.Y(n_4391)
);

AND2x2_ASAP7_75t_L g4392 ( 
.A(n_4275),
.B(n_4185),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4250),
.B(n_4208),
.Y(n_4393)
);

NAND2xp5_ASAP7_75t_SL g4394 ( 
.A(n_4294),
.B(n_4172),
.Y(n_4394)
);

OAI21xp5_ASAP7_75t_SL g4395 ( 
.A1(n_4284),
.A2(n_4035),
.B(n_4131),
.Y(n_4395)
);

AND2x2_ASAP7_75t_L g4396 ( 
.A(n_4251),
.B(n_4208),
.Y(n_4396)
);

OAI21xp33_ASAP7_75t_L g4397 ( 
.A1(n_4263),
.A2(n_3957),
.B(n_3751),
.Y(n_4397)
);

OAI22xp5_ASAP7_75t_L g4398 ( 
.A1(n_4340),
.A2(n_4202),
.B1(n_4184),
.B2(n_4054),
.Y(n_4398)
);

NAND3xp33_ASAP7_75t_L g4399 ( 
.A(n_4321),
.B(n_4223),
.C(n_4149),
.Y(n_4399)
);

OAI21xp5_ASAP7_75t_SL g4400 ( 
.A1(n_4362),
.A2(n_3664),
.B(n_3701),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_4353),
.B(n_4308),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4257),
.B(n_4220),
.Y(n_4402)
);

NAND4xp25_ASAP7_75t_L g4403 ( 
.A(n_4343),
.B(n_3699),
.C(n_3789),
.D(n_3912),
.Y(n_4403)
);

OAI221xp5_ASAP7_75t_SL g4404 ( 
.A1(n_4336),
.A2(n_3960),
.B1(n_4114),
.B2(n_4113),
.C(n_4197),
.Y(n_4404)
);

NAND3xp33_ASAP7_75t_L g4405 ( 
.A(n_4364),
.B(n_4221),
.C(n_4138),
.Y(n_4405)
);

NOR3xp33_ASAP7_75t_L g4406 ( 
.A(n_4314),
.B(n_4145),
.C(n_4164),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_4342),
.B(n_4109),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_4356),
.B(n_4051),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4278),
.B(n_4052),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4279),
.B(n_4205),
.Y(n_4410)
);

NAND3xp33_ASAP7_75t_L g4411 ( 
.A(n_4288),
.B(n_4181),
.C(n_4165),
.Y(n_4411)
);

AOI22xp33_ASAP7_75t_L g4412 ( 
.A1(n_4316),
.A2(n_4093),
.B1(n_4113),
.B2(n_4111),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4323),
.B(n_4220),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4268),
.B(n_4154),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4280),
.B(n_4211),
.Y(n_4415)
);

NOR2xp33_ASAP7_75t_L g4416 ( 
.A(n_4252),
.B(n_4086),
.Y(n_4416)
);

OAI21xp5_ASAP7_75t_SL g4417 ( 
.A1(n_4294),
.A2(n_4063),
.B(n_3659),
.Y(n_4417)
);

NAND3xp33_ASAP7_75t_L g4418 ( 
.A(n_4295),
.B(n_3874),
.C(n_4116),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4286),
.B(n_4302),
.Y(n_4419)
);

NOR2xp33_ASAP7_75t_SL g4420 ( 
.A(n_4294),
.B(n_3685),
.Y(n_4420)
);

AOI221xp5_ASAP7_75t_L g4421 ( 
.A1(n_4235),
.A2(n_4088),
.B1(n_3772),
.B2(n_4058),
.C(n_3903),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4304),
.B(n_4213),
.Y(n_4422)
);

NAND3xp33_ASAP7_75t_L g4423 ( 
.A(n_4318),
.B(n_4319),
.C(n_4301),
.Y(n_4423)
);

INVx1_ASAP7_75t_L g4424 ( 
.A(n_4258),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4313),
.B(n_4315),
.Y(n_4425)
);

OAI21xp33_ASAP7_75t_L g4426 ( 
.A1(n_4310),
.A2(n_3700),
.B(n_4222),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_4290),
.B(n_4177),
.Y(n_4427)
);

AOI22xp33_ASAP7_75t_L g4428 ( 
.A1(n_4326),
.A2(n_4093),
.B1(n_4111),
.B2(n_3984),
.Y(n_4428)
);

OAI22xp5_ASAP7_75t_L g4429 ( 
.A1(n_4349),
.A2(n_3691),
.B1(n_4000),
.B2(n_4006),
.Y(n_4429)
);

AOI21xp33_ASAP7_75t_L g4430 ( 
.A1(n_4283),
.A2(n_4215),
.B(n_4210),
.Y(n_4430)
);

NAND2xp5_ASAP7_75t_L g4431 ( 
.A(n_4328),
.B(n_4092),
.Y(n_4431)
);

NAND2xp5_ASAP7_75t_SL g4432 ( 
.A(n_4332),
.B(n_4042),
.Y(n_4432)
);

NAND2xp5_ASAP7_75t_SL g4433 ( 
.A(n_4332),
.B(n_4042),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4337),
.B(n_4094),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4357),
.B(n_4139),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4346),
.B(n_4022),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4363),
.B(n_4147),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4238),
.B(n_4225),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4238),
.B(n_4239),
.Y(n_4439)
);

AND2x2_ASAP7_75t_L g4440 ( 
.A(n_4335),
.B(n_4084),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4239),
.B(n_4228),
.Y(n_4441)
);

AND2x2_ASAP7_75t_L g4442 ( 
.A(n_4247),
.B(n_4084),
.Y(n_4442)
);

NAND3xp33_ASAP7_75t_L g4443 ( 
.A(n_4281),
.B(n_3824),
.C(n_4215),
.Y(n_4443)
);

NAND3xp33_ASAP7_75t_L g4444 ( 
.A(n_4236),
.B(n_4166),
.C(n_4224),
.Y(n_4444)
);

OAI221xp5_ASAP7_75t_L g4445 ( 
.A1(n_4333),
.A2(n_3721),
.B1(n_3890),
.B2(n_3967),
.C(n_4137),
.Y(n_4445)
);

AND2x2_ASAP7_75t_L g4446 ( 
.A(n_4237),
.B(n_4065),
.Y(n_4446)
);

NAND4xp25_ASAP7_75t_L g4447 ( 
.A(n_4306),
.B(n_3791),
.C(n_3633),
.D(n_3748),
.Y(n_4447)
);

NOR3xp33_ASAP7_75t_L g4448 ( 
.A(n_4297),
.B(n_3895),
.C(n_3959),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4240),
.B(n_4066),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4237),
.B(n_4151),
.Y(n_4450)
);

NAND2xp5_ASAP7_75t_SL g4451 ( 
.A(n_4332),
.B(n_4012),
.Y(n_4451)
);

NAND3xp33_ASAP7_75t_L g4452 ( 
.A(n_4243),
.B(n_4168),
.C(n_4124),
.Y(n_4452)
);

NOR2xp33_ASAP7_75t_L g4453 ( 
.A(n_4253),
.B(n_4057),
.Y(n_4453)
);

AND2x2_ASAP7_75t_L g4454 ( 
.A(n_4243),
.B(n_4179),
.Y(n_4454)
);

NOR3xp33_ASAP7_75t_L g4455 ( 
.A(n_4341),
.B(n_3914),
.C(n_3858),
.Y(n_4455)
);

OAI221xp5_ASAP7_75t_L g4456 ( 
.A1(n_4366),
.A2(n_3832),
.B1(n_4122),
.B2(n_3703),
.C(n_3878),
.Y(n_4456)
);

AND2x2_ASAP7_75t_L g4457 ( 
.A(n_4249),
.B(n_4167),
.Y(n_4457)
);

NAND2xp5_ASAP7_75t_SL g4458 ( 
.A(n_4352),
.B(n_4193),
.Y(n_4458)
);

NAND4xp25_ASAP7_75t_L g4459 ( 
.A(n_4307),
.B(n_3624),
.C(n_3767),
.D(n_3760),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4249),
.B(n_4127),
.Y(n_4460)
);

OAI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4345),
.A2(n_4000),
.B1(n_4144),
.B2(n_3825),
.Y(n_4461)
);

NOR2xp33_ASAP7_75t_L g4462 ( 
.A(n_4352),
.B(n_4187),
.Y(n_4462)
);

OAI22xp5_ASAP7_75t_L g4463 ( 
.A1(n_4347),
.A2(n_4144),
.B1(n_3776),
.B2(n_3983),
.Y(n_4463)
);

AND2x2_ASAP7_75t_SL g4464 ( 
.A(n_4327),
.B(n_3642),
.Y(n_4464)
);

AOI221xp5_ASAP7_75t_L g4465 ( 
.A1(n_4261),
.A2(n_3629),
.B1(n_3976),
.B2(n_3972),
.C(n_4117),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4240),
.B(n_4140),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_4242),
.B(n_4142),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4390),
.Y(n_4468)
);

INVx1_ASAP7_75t_SL g4469 ( 
.A(n_4372),
.Y(n_4469)
);

INVxp67_ASAP7_75t_L g4470 ( 
.A(n_4391),
.Y(n_4470)
);

OR2x2_ASAP7_75t_L g4471 ( 
.A(n_4401),
.B(n_4330),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4439),
.Y(n_4472)
);

AND2x4_ASAP7_75t_L g4473 ( 
.A(n_4368),
.B(n_4339),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4419),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4425),
.Y(n_4475)
);

INVx2_ASAP7_75t_L g4476 ( 
.A(n_4424),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4446),
.Y(n_4477)
);

INVx2_ASAP7_75t_L g4478 ( 
.A(n_4460),
.Y(n_4478)
);

AND2x2_ASAP7_75t_L g4479 ( 
.A(n_4450),
.B(n_4309),
.Y(n_4479)
);

INVx3_ASAP7_75t_L g4480 ( 
.A(n_4464),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4436),
.Y(n_4481)
);

AND2x2_ASAP7_75t_L g4482 ( 
.A(n_4392),
.B(n_4348),
.Y(n_4482)
);

INVx2_ASAP7_75t_L g4483 ( 
.A(n_4382),
.Y(n_4483)
);

OR2x2_ASAP7_75t_L g4484 ( 
.A(n_4408),
.B(n_4344),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4454),
.B(n_4350),
.Y(n_4485)
);

NOR2xp67_ASAP7_75t_L g4486 ( 
.A(n_4395),
.B(n_4233),
.Y(n_4486)
);

AND2x2_ASAP7_75t_L g4487 ( 
.A(n_4457),
.B(n_4265),
.Y(n_4487)
);

AND2x2_ASAP7_75t_L g4488 ( 
.A(n_4402),
.B(n_4262),
.Y(n_4488)
);

HB1xp67_ASAP7_75t_L g4489 ( 
.A(n_4385),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4393),
.B(n_4270),
.Y(n_4490)
);

OR2x2_ASAP7_75t_L g4491 ( 
.A(n_4384),
.B(n_4355),
.Y(n_4491)
);

HB1xp67_ASAP7_75t_L g4492 ( 
.A(n_4387),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4409),
.Y(n_4493)
);

INVx3_ASAP7_75t_L g4494 ( 
.A(n_4368),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4431),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_4406),
.B(n_4272),
.Y(n_4496)
);

INVx2_ASAP7_75t_L g4497 ( 
.A(n_4466),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4396),
.B(n_4277),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_4410),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_4415),
.Y(n_4500)
);

NAND2xp5_ASAP7_75t_L g4501 ( 
.A(n_4379),
.B(n_4282),
.Y(n_4501)
);

AND2x2_ASAP7_75t_SL g4502 ( 
.A(n_4420),
.B(n_3642),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4467),
.Y(n_4503)
);

OR2x2_ASAP7_75t_L g4504 ( 
.A(n_4371),
.B(n_4365),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4438),
.Y(n_4505)
);

OA21x2_ASAP7_75t_L g4506 ( 
.A1(n_4426),
.A2(n_4074),
.B(n_4190),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4440),
.B(n_4289),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_4441),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4377),
.B(n_4291),
.Y(n_4509)
);

HB1xp67_ASAP7_75t_L g4510 ( 
.A(n_4407),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4442),
.B(n_4296),
.Y(n_4511)
);

OR2x2_ASAP7_75t_L g4512 ( 
.A(n_4389),
.B(n_4367),
.Y(n_4512)
);

INVx2_ASAP7_75t_SL g4513 ( 
.A(n_4458),
.Y(n_4513)
);

OR2x2_ASAP7_75t_L g4514 ( 
.A(n_4423),
.B(n_4241),
.Y(n_4514)
);

AND2x4_ASAP7_75t_L g4515 ( 
.A(n_4405),
.B(n_4399),
.Y(n_4515)
);

INVx2_ASAP7_75t_L g4516 ( 
.A(n_4449),
.Y(n_4516)
);

AND2x4_ASAP7_75t_L g4517 ( 
.A(n_4411),
.B(n_4334),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4437),
.B(n_4311),
.Y(n_4518)
);

INVx2_ASAP7_75t_SL g4519 ( 
.A(n_4413),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4375),
.B(n_4324),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4370),
.B(n_4351),
.Y(n_4521)
);

NOR2x1_ASAP7_75t_L g4522 ( 
.A(n_4417),
.B(n_4176),
.Y(n_4522)
);

INVx1_ASAP7_75t_L g4523 ( 
.A(n_4422),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4434),
.Y(n_4524)
);

NAND2x1p5_ASAP7_75t_L g4525 ( 
.A(n_4451),
.B(n_3854),
.Y(n_4525)
);

INVxp67_ASAP7_75t_SL g4526 ( 
.A(n_4388),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4435),
.Y(n_4527)
);

INVx2_ASAP7_75t_L g4528 ( 
.A(n_4376),
.Y(n_4528)
);

INVxp67_ASAP7_75t_L g4529 ( 
.A(n_4462),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4414),
.B(n_4354),
.Y(n_4530)
);

AND2x2_ASAP7_75t_L g4531 ( 
.A(n_4427),
.B(n_4255),
.Y(n_4531)
);

AND2x2_ASAP7_75t_SL g4532 ( 
.A(n_4412),
.B(n_4428),
.Y(n_4532)
);

OR2x2_ASAP7_75t_L g4533 ( 
.A(n_4444),
.B(n_4259),
.Y(n_4533)
);

AND2x4_ASAP7_75t_L g4534 ( 
.A(n_4432),
.B(n_4334),
.Y(n_4534)
);

NAND2xp5_ASAP7_75t_L g4535 ( 
.A(n_4380),
.B(n_4360),
.Y(n_4535)
);

NOR2x1_ASAP7_75t_SL g4536 ( 
.A(n_4433),
.B(n_3688),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4426),
.B(n_4360),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4373),
.Y(n_4538)
);

HB1xp67_ASAP7_75t_L g4539 ( 
.A(n_4416),
.Y(n_4539)
);

INVx1_ASAP7_75t_L g4540 ( 
.A(n_4374),
.Y(n_4540)
);

INVx1_ASAP7_75t_SL g4541 ( 
.A(n_4453),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_4461),
.B(n_4398),
.Y(n_4542)
);

AND2x2_ASAP7_75t_L g4543 ( 
.A(n_4463),
.B(n_4264),
.Y(n_4543)
);

NOR2xp33_ASAP7_75t_L g4544 ( 
.A(n_4378),
.B(n_4369),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4430),
.B(n_4267),
.Y(n_4545)
);

INVx2_ASAP7_75t_L g4546 ( 
.A(n_4452),
.Y(n_4546)
);

AND2x2_ASAP7_75t_L g4547 ( 
.A(n_4394),
.B(n_4325),
.Y(n_4547)
);

NAND2xp5_ASAP7_75t_L g4548 ( 
.A(n_4465),
.B(n_4242),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4474),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4494),
.B(n_4429),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4474),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4475),
.Y(n_4552)
);

OR2x2_ASAP7_75t_L g4553 ( 
.A(n_4491),
.B(n_4329),
.Y(n_4553)
);

INVx2_ASAP7_75t_L g4554 ( 
.A(n_4533),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4494),
.B(n_4381),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4475),
.Y(n_4556)
);

AND2x2_ASAP7_75t_L g4557 ( 
.A(n_4538),
.B(n_4418),
.Y(n_4557)
);

INVx1_ASAP7_75t_L g4558 ( 
.A(n_4472),
.Y(n_4558)
);

AND2x2_ASAP7_75t_L g4559 ( 
.A(n_4538),
.B(n_4540),
.Y(n_4559)
);

AND2x4_ASAP7_75t_L g4560 ( 
.A(n_4473),
.B(n_4418),
.Y(n_4560)
);

INVxp67_ASAP7_75t_L g4561 ( 
.A(n_4544),
.Y(n_4561)
);

OR2x2_ASAP7_75t_L g4562 ( 
.A(n_4512),
.B(n_4358),
.Y(n_4562)
);

INVx1_ASAP7_75t_SL g4563 ( 
.A(n_4522),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4540),
.B(n_4448),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4472),
.Y(n_4565)
);

NOR2xp33_ASAP7_75t_L g4566 ( 
.A(n_4529),
.B(n_4386),
.Y(n_4566)
);

OR2x2_ASAP7_75t_L g4567 ( 
.A(n_4471),
.B(n_4404),
.Y(n_4567)
);

OR2x2_ASAP7_75t_L g4568 ( 
.A(n_4484),
.B(n_4245),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4548),
.B(n_4245),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4499),
.Y(n_4570)
);

BUFx2_ASAP7_75t_SL g4571 ( 
.A(n_4534),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4499),
.Y(n_4572)
);

OAI21xp33_ASAP7_75t_SL g4573 ( 
.A1(n_4489),
.A2(n_3994),
.B(n_4200),
.Y(n_4573)
);

INVx2_ASAP7_75t_L g4574 ( 
.A(n_4534),
.Y(n_4574)
);

AND2x2_ASAP7_75t_L g4575 ( 
.A(n_4542),
.B(n_4397),
.Y(n_4575)
);

AND2x2_ASAP7_75t_L g4576 ( 
.A(n_4543),
.B(n_4397),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4504),
.B(n_4292),
.Y(n_4577)
);

NOR3xp33_ASAP7_75t_L g4578 ( 
.A(n_4526),
.B(n_4383),
.C(n_4445),
.Y(n_4578)
);

HB1xp67_ASAP7_75t_L g4579 ( 
.A(n_4514),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_4546),
.B(n_4292),
.Y(n_4580)
);

OR2x2_ASAP7_75t_L g4581 ( 
.A(n_4497),
.B(n_4298),
.Y(n_4581)
);

AND2x2_ASAP7_75t_L g4582 ( 
.A(n_4545),
.B(n_4298),
.Y(n_4582)
);

INVx2_ASAP7_75t_L g4583 ( 
.A(n_4468),
.Y(n_4583)
);

INVx1_ASAP7_75t_L g4584 ( 
.A(n_4500),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4500),
.Y(n_4585)
);

AND2x2_ASAP7_75t_L g4586 ( 
.A(n_4513),
.B(n_4300),
.Y(n_4586)
);

OAI21xp33_ASAP7_75t_L g4587 ( 
.A1(n_4532),
.A2(n_4400),
.B(n_4447),
.Y(n_4587)
);

AND2x4_ASAP7_75t_L g4588 ( 
.A(n_4473),
.B(n_4300),
.Y(n_4588)
);

OR2x2_ASAP7_75t_L g4589 ( 
.A(n_4503),
.B(n_4303),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_L g4590 ( 
.A(n_4496),
.B(n_4303),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4523),
.Y(n_4591)
);

INVx2_ASAP7_75t_L g4592 ( 
.A(n_4476),
.Y(n_4592)
);

OR2x2_ASAP7_75t_L g4593 ( 
.A(n_4505),
.B(n_4331),
.Y(n_4593)
);

OR2x2_ASAP7_75t_L g4594 ( 
.A(n_4508),
.B(n_4331),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4523),
.Y(n_4595)
);

INVxp33_ASAP7_75t_L g4596 ( 
.A(n_4486),
.Y(n_4596)
);

OR2x2_ASAP7_75t_L g4597 ( 
.A(n_4516),
.B(n_4230),
.Y(n_4597)
);

NOR2x1p5_ASAP7_75t_L g4598 ( 
.A(n_4480),
.B(n_4403),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_4524),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_4539),
.B(n_4455),
.Y(n_4600)
);

INVxp67_ASAP7_75t_L g4601 ( 
.A(n_4541),
.Y(n_4601)
);

INVx1_ASAP7_75t_L g4602 ( 
.A(n_4524),
.Y(n_4602)
);

NOR2x1_ASAP7_75t_L g4603 ( 
.A(n_4517),
.B(n_4443),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4492),
.B(n_4231),
.Y(n_4604)
);

INVx1_ASAP7_75t_L g4605 ( 
.A(n_4493),
.Y(n_4605)
);

INVx1_ASAP7_75t_L g4606 ( 
.A(n_4481),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4515),
.B(n_4421),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4495),
.Y(n_4608)
);

OR2x2_ASAP7_75t_L g4609 ( 
.A(n_4580),
.B(n_4535),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4581),
.Y(n_4610)
);

AND2x2_ASAP7_75t_L g4611 ( 
.A(n_4571),
.B(n_4517),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4571),
.B(n_4560),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4559),
.B(n_4515),
.Y(n_4613)
);

AND2x4_ASAP7_75t_L g4614 ( 
.A(n_4560),
.B(n_4480),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_L g4615 ( 
.A(n_4564),
.B(n_4557),
.Y(n_4615)
);

OAI22xp33_ASAP7_75t_L g4616 ( 
.A1(n_4563),
.A2(n_4469),
.B1(n_4519),
.B2(n_4525),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4555),
.B(n_4547),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_L g4618 ( 
.A(n_4607),
.B(n_4501),
.Y(n_4618)
);

HB1xp67_ASAP7_75t_L g4619 ( 
.A(n_4579),
.Y(n_4619)
);

AND2x2_ASAP7_75t_L g4620 ( 
.A(n_4550),
.B(n_4574),
.Y(n_4620)
);

AND2x2_ASAP7_75t_L g4621 ( 
.A(n_4588),
.B(n_4510),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4589),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4588),
.B(n_4482),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4575),
.B(n_4527),
.Y(n_4624)
);

INVx1_ASAP7_75t_SL g4625 ( 
.A(n_4600),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4562),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_4569),
.B(n_4520),
.Y(n_4627)
);

OAI21xp5_ASAP7_75t_L g4628 ( 
.A1(n_4587),
.A2(n_4502),
.B(n_4537),
.Y(n_4628)
);

OR2x2_ASAP7_75t_L g4629 ( 
.A(n_4568),
.B(n_4521),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4582),
.B(n_4470),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4554),
.B(n_4487),
.Y(n_4631)
);

INVx1_ASAP7_75t_SL g4632 ( 
.A(n_4596),
.Y(n_4632)
);

NAND2x1_ASAP7_75t_L g4633 ( 
.A(n_4603),
.B(n_4528),
.Y(n_4633)
);

NAND2xp5_ASAP7_75t_L g4634 ( 
.A(n_4608),
.B(n_4527),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_4597),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4577),
.Y(n_4636)
);

AND2x2_ASAP7_75t_L g4637 ( 
.A(n_4576),
.B(n_4483),
.Y(n_4637)
);

INVx1_ASAP7_75t_L g4638 ( 
.A(n_4608),
.Y(n_4638)
);

INVxp67_ASAP7_75t_L g4639 ( 
.A(n_4566),
.Y(n_4639)
);

OR2x6_ASAP7_75t_L g4640 ( 
.A(n_4601),
.B(n_3854),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4593),
.Y(n_4641)
);

BUFx2_ASAP7_75t_L g4642 ( 
.A(n_4573),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4605),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4606),
.Y(n_4644)
);

OR2x2_ASAP7_75t_L g4645 ( 
.A(n_4604),
.B(n_4477),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4599),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4602),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4594),
.Y(n_4648)
);

OR2x2_ASAP7_75t_SL g4649 ( 
.A(n_4567),
.B(n_4536),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4561),
.B(n_4509),
.Y(n_4650)
);

OAI21xp5_ASAP7_75t_L g4651 ( 
.A1(n_4578),
.A2(n_4456),
.B(n_4459),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_L g4652 ( 
.A(n_4570),
.B(n_4572),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4586),
.B(n_4485),
.Y(n_4653)
);

NOR2xp33_ASAP7_75t_L g4654 ( 
.A(n_4590),
.B(n_3627),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4553),
.Y(n_4655)
);

INVxp67_ASAP7_75t_SL g4656 ( 
.A(n_4598),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4584),
.Y(n_4657)
);

NAND2xp5_ASAP7_75t_L g4658 ( 
.A(n_4585),
.B(n_4518),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_L g4659 ( 
.A(n_4591),
.B(n_4488),
.Y(n_4659)
);

OR2x2_ASAP7_75t_L g4660 ( 
.A(n_4549),
.B(n_4478),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4551),
.B(n_4490),
.Y(n_4661)
);

OR2x6_ASAP7_75t_L g4662 ( 
.A(n_4595),
.B(n_3765),
.Y(n_4662)
);

NOR2xp33_ASAP7_75t_L g4663 ( 
.A(n_4552),
.B(n_3671),
.Y(n_4663)
);

INVx1_ASAP7_75t_L g4664 ( 
.A(n_4556),
.Y(n_4664)
);

INVx3_ASAP7_75t_L g4665 ( 
.A(n_4583),
.Y(n_4665)
);

AND2x2_ASAP7_75t_L g4666 ( 
.A(n_4558),
.B(n_4498),
.Y(n_4666)
);

BUFx2_ASAP7_75t_L g4667 ( 
.A(n_4565),
.Y(n_4667)
);

AOI211xp5_ASAP7_75t_L g4668 ( 
.A1(n_4592),
.A2(n_3920),
.B(n_3916),
.C(n_3697),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4562),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4619),
.Y(n_4670)
);

AOI22xp5_ASAP7_75t_L g4671 ( 
.A1(n_4656),
.A2(n_3947),
.B1(n_3975),
.B2(n_4158),
.Y(n_4671)
);

INVx2_ASAP7_75t_L g4672 ( 
.A(n_4665),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4612),
.B(n_4611),
.Y(n_4673)
);

INVx1_ASAP7_75t_SL g4674 ( 
.A(n_4640),
.Y(n_4674)
);

NOR2x1_ASAP7_75t_L g4675 ( 
.A(n_4640),
.B(n_3939),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4639),
.B(n_4530),
.Y(n_4676)
);

NOR2xp33_ASAP7_75t_L g4677 ( 
.A(n_4632),
.B(n_4195),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4634),
.Y(n_4678)
);

INVx1_ASAP7_75t_L g4679 ( 
.A(n_4652),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4626),
.Y(n_4680)
);

HB1xp67_ASAP7_75t_L g4681 ( 
.A(n_4625),
.Y(n_4681)
);

HB1xp67_ASAP7_75t_L g4682 ( 
.A(n_4667),
.Y(n_4682)
);

INVx1_ASAP7_75t_L g4683 ( 
.A(n_4669),
.Y(n_4683)
);

HB1xp67_ASAP7_75t_L g4684 ( 
.A(n_4643),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4658),
.Y(n_4685)
);

INVx4_ASAP7_75t_L g4686 ( 
.A(n_4662),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_R g4687 ( 
.A(n_4614),
.B(n_3968),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4665),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4624),
.B(n_4531),
.Y(n_4689)
);

AOI22xp33_ASAP7_75t_L g4690 ( 
.A1(n_4614),
.A2(n_4506),
.B1(n_4192),
.B2(n_4479),
.Y(n_4690)
);

INVx1_ASAP7_75t_SL g4691 ( 
.A(n_4649),
.Y(n_4691)
);

HB1xp67_ASAP7_75t_L g4692 ( 
.A(n_4644),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4617),
.B(n_4511),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4650),
.Y(n_4694)
);

AOI22xp33_ASAP7_75t_L g4695 ( 
.A1(n_4651),
.A2(n_4506),
.B1(n_4192),
.B2(n_3923),
.Y(n_4695)
);

AOI22xp5_ASAP7_75t_L g4696 ( 
.A1(n_4615),
.A2(n_3965),
.B1(n_3939),
.B2(n_4195),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4620),
.Y(n_4697)
);

INVx2_ASAP7_75t_L g4698 ( 
.A(n_4645),
.Y(n_4698)
);

XNOR2x2_ASAP7_75t_L g4699 ( 
.A(n_4628),
.B(n_4126),
.Y(n_4699)
);

AOI22xp33_ASAP7_75t_L g4700 ( 
.A1(n_4642),
.A2(n_4507),
.B1(n_3922),
.B2(n_3882),
.Y(n_4700)
);

AND2x2_ASAP7_75t_L g4701 ( 
.A(n_4621),
.B(n_4536),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4637),
.B(n_4218),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4638),
.Y(n_4703)
);

AOI22xp5_ASAP7_75t_L g4704 ( 
.A1(n_4618),
.A2(n_4135),
.B1(n_3739),
.B2(n_3938),
.Y(n_4704)
);

INVx1_ASAP7_75t_L g4705 ( 
.A(n_4629),
.Y(n_4705)
);

INVx1_ASAP7_75t_SL g4706 ( 
.A(n_4662),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4646),
.Y(n_4707)
);

INVx1_ASAP7_75t_L g4708 ( 
.A(n_4681),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4670),
.Y(n_4709)
);

NAND2xp33_ASAP7_75t_L g4710 ( 
.A(n_4675),
.B(n_4613),
.Y(n_4710)
);

INVxp67_ASAP7_75t_L g4711 ( 
.A(n_4677),
.Y(n_4711)
);

INVx1_ASAP7_75t_L g4712 ( 
.A(n_4680),
.Y(n_4712)
);

INVxp67_ASAP7_75t_L g4713 ( 
.A(n_4671),
.Y(n_4713)
);

AOI22xp5_ASAP7_75t_L g4714 ( 
.A1(n_4674),
.A2(n_4616),
.B1(n_4663),
.B2(n_4654),
.Y(n_4714)
);

OR2x2_ASAP7_75t_L g4715 ( 
.A(n_4683),
.B(n_4705),
.Y(n_4715)
);

OAI211xp5_ASAP7_75t_L g4716 ( 
.A1(n_4691),
.A2(n_4668),
.B(n_4633),
.C(n_4636),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4682),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4694),
.B(n_4627),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4673),
.B(n_4610),
.Y(n_4719)
);

A2O1A1Ixp33_ASAP7_75t_L g4720 ( 
.A1(n_4706),
.A2(n_4609),
.B(n_4622),
.C(n_4610),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4701),
.B(n_4623),
.Y(n_4721)
);

NAND3xp33_ASAP7_75t_L g4722 ( 
.A(n_4686),
.B(n_4657),
.C(n_4647),
.Y(n_4722)
);

OAI22xp33_ASAP7_75t_SL g4723 ( 
.A1(n_4686),
.A2(n_4664),
.B1(n_4622),
.B2(n_4641),
.Y(n_4723)
);

INVxp67_ASAP7_75t_L g4724 ( 
.A(n_4671),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4698),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4684),
.Y(n_4726)
);

AOI21xp33_ASAP7_75t_L g4727 ( 
.A1(n_4692),
.A2(n_4641),
.B(n_3944),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4672),
.Y(n_4728)
);

AOI22xp33_ASAP7_75t_L g4729 ( 
.A1(n_4699),
.A2(n_4655),
.B1(n_4648),
.B2(n_4635),
.Y(n_4729)
);

INVxp67_ASAP7_75t_L g4730 ( 
.A(n_4696),
.Y(n_4730)
);

OR2x2_ASAP7_75t_L g4731 ( 
.A(n_4678),
.B(n_4660),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4688),
.Y(n_4732)
);

OAI21xp5_ASAP7_75t_L g4733 ( 
.A1(n_4696),
.A2(n_4630),
.B(n_4659),
.Y(n_4733)
);

NOR2xp33_ASAP7_75t_L g4734 ( 
.A(n_4697),
.B(n_4631),
.Y(n_4734)
);

OAI221xp5_ASAP7_75t_L g4735 ( 
.A1(n_4695),
.A2(n_3881),
.B1(n_3737),
.B2(n_3794),
.C(n_3894),
.Y(n_4735)
);

OR2x2_ASAP7_75t_L g4736 ( 
.A(n_4679),
.B(n_4661),
.Y(n_4736)
);

OAI221xp5_ASAP7_75t_L g4737 ( 
.A1(n_4700),
.A2(n_3951),
.B1(n_3921),
.B2(n_3790),
.C(n_3649),
.Y(n_4737)
);

BUFx2_ASAP7_75t_L g4738 ( 
.A(n_4711),
.Y(n_4738)
);

OAI21xp5_ASAP7_75t_SL g4739 ( 
.A1(n_4730),
.A2(n_4704),
.B(n_4690),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_4708),
.B(n_4685),
.Y(n_4740)
);

AND2x2_ASAP7_75t_L g4741 ( 
.A(n_4721),
.B(n_4693),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4726),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4713),
.B(n_4676),
.Y(n_4743)
);

AND2x2_ASAP7_75t_L g4744 ( 
.A(n_4714),
.B(n_4653),
.Y(n_4744)
);

AND2x2_ASAP7_75t_L g4745 ( 
.A(n_4714),
.B(n_4702),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4715),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4725),
.Y(n_4747)
);

INVx2_ASAP7_75t_SL g4748 ( 
.A(n_4728),
.Y(n_4748)
);

INVx1_ASAP7_75t_SL g4749 ( 
.A(n_4717),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_4724),
.B(n_4707),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4733),
.B(n_4689),
.Y(n_4751)
);

INVxp67_ASAP7_75t_L g4752 ( 
.A(n_4709),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4732),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4720),
.B(n_4703),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4712),
.B(n_4704),
.Y(n_4755)
);

AND2x2_ASAP7_75t_L g4756 ( 
.A(n_4729),
.B(n_4666),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4734),
.B(n_4687),
.Y(n_4757)
);

NAND2xp33_ASAP7_75t_L g4758 ( 
.A(n_4719),
.B(n_3922),
.Y(n_4758)
);

NAND2xp5_ASAP7_75t_L g4759 ( 
.A(n_4723),
.B(n_3762),
.Y(n_4759)
);

AND2x2_ASAP7_75t_L g4760 ( 
.A(n_4710),
.B(n_3956),
.Y(n_4760)
);

NOR2xp33_ASAP7_75t_L g4761 ( 
.A(n_4716),
.B(n_3961),
.Y(n_4761)
);

HB1xp67_ASAP7_75t_L g4762 ( 
.A(n_4718),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4736),
.B(n_4727),
.Y(n_4763)
);

OR2x2_ASAP7_75t_L g4764 ( 
.A(n_4747),
.B(n_4731),
.Y(n_4764)
);

OAI21xp33_ASAP7_75t_L g4765 ( 
.A1(n_4739),
.A2(n_4722),
.B(n_4735),
.Y(n_4765)
);

OAI211xp5_ASAP7_75t_L g4766 ( 
.A1(n_4738),
.A2(n_4739),
.B(n_4761),
.C(n_4742),
.Y(n_4766)
);

OAI21xp5_ASAP7_75t_L g4767 ( 
.A1(n_4748),
.A2(n_4737),
.B(n_3973),
.Y(n_4767)
);

AOI22xp5_ASAP7_75t_L g4768 ( 
.A1(n_4745),
.A2(n_3882),
.B1(n_3770),
.B2(n_3889),
.Y(n_4768)
);

OAI21xp5_ASAP7_75t_SL g4769 ( 
.A1(n_4760),
.A2(n_3847),
.B(n_3815),
.Y(n_4769)
);

OAI221xp5_ASAP7_75t_L g4770 ( 
.A1(n_4749),
.A2(n_3693),
.B1(n_3808),
.B2(n_3774),
.C(n_3899),
.Y(n_4770)
);

OAI211xp5_ASAP7_75t_L g4771 ( 
.A1(n_4749),
.A2(n_3850),
.B(n_3940),
.C(n_3991),
.Y(n_4771)
);

OAI211xp5_ASAP7_75t_L g4772 ( 
.A1(n_4762),
.A2(n_3934),
.B(n_3928),
.C(n_3900),
.Y(n_4772)
);

AOI221xp5_ASAP7_75t_L g4773 ( 
.A1(n_4746),
.A2(n_3755),
.B1(n_3800),
.B2(n_3872),
.C(n_3780),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4753),
.Y(n_4774)
);

AOI21xp5_ASAP7_75t_L g4775 ( 
.A1(n_4754),
.A2(n_3778),
.B(n_3569),
.Y(n_4775)
);

OAI32xp33_ASAP7_75t_L g4776 ( 
.A1(n_4743),
.A2(n_3688),
.A3(n_3966),
.B1(n_3964),
.B2(n_3564),
.Y(n_4776)
);

INVx1_ASAP7_75t_L g4777 ( 
.A(n_4740),
.Y(n_4777)
);

A2O1A1Ixp33_ASAP7_75t_L g4778 ( 
.A1(n_4744),
.A2(n_3880),
.B(n_3831),
.C(n_3539),
.Y(n_4778)
);

NAND3xp33_ASAP7_75t_SL g4779 ( 
.A(n_4740),
.B(n_3919),
.C(n_3907),
.Y(n_4779)
);

AOI321xp33_ASAP7_75t_L g4780 ( 
.A1(n_4755),
.A2(n_4194),
.A3(n_4173),
.B1(n_4191),
.B2(n_4180),
.C(n_3625),
.Y(n_4780)
);

OAI211xp5_ASAP7_75t_SL g4781 ( 
.A1(n_4752),
.A2(n_3565),
.B(n_3988),
.C(n_3575),
.Y(n_4781)
);

NOR2x1_ASAP7_75t_L g4782 ( 
.A(n_4766),
.B(n_4750),
.Y(n_4782)
);

INVxp67_ASAP7_75t_L g4783 ( 
.A(n_4774),
.Y(n_4783)
);

AO22x2_ASAP7_75t_L g4784 ( 
.A1(n_4777),
.A2(n_4755),
.B1(n_4759),
.B2(n_4751),
.Y(n_4784)
);

NOR3xp33_ASAP7_75t_L g4785 ( 
.A(n_4765),
.B(n_4763),
.C(n_4756),
.Y(n_4785)
);

OAI21xp33_ASAP7_75t_SL g4786 ( 
.A1(n_4764),
.A2(n_4741),
.B(n_4757),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4767),
.B(n_4758),
.Y(n_4787)
);

NAND4xp25_ASAP7_75t_L g4788 ( 
.A(n_4778),
.B(n_3949),
.C(n_3548),
.D(n_4152),
.Y(n_4788)
);

NOR3xp33_ASAP7_75t_L g4789 ( 
.A(n_4776),
.B(n_3793),
.C(n_3753),
.Y(n_4789)
);

NAND3xp33_ASAP7_75t_L g4790 ( 
.A(n_4775),
.B(n_3797),
.C(n_3783),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4772),
.Y(n_4791)
);

AO22x2_ASAP7_75t_L g4792 ( 
.A1(n_4779),
.A2(n_3915),
.B1(n_3936),
.B2(n_3909),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4780),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4768),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4792),
.Y(n_4795)
);

NAND3xp33_ASAP7_75t_L g4796 ( 
.A(n_4783),
.B(n_4769),
.C(n_4771),
.Y(n_4796)
);

NOR2xp33_ASAP7_75t_L g4797 ( 
.A(n_4786),
.B(n_4781),
.Y(n_4797)
);

NOR2xp33_ASAP7_75t_L g4798 ( 
.A(n_4791),
.B(n_4770),
.Y(n_4798)
);

NOR5xp2_ASAP7_75t_L g4799 ( 
.A(n_4793),
.B(n_4773),
.C(n_3694),
.D(n_3242),
.E(n_887),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4792),
.Y(n_4800)
);

OAI21xp33_ASAP7_75t_SL g4801 ( 
.A1(n_4782),
.A2(n_3891),
.B(n_3817),
.Y(n_4801)
);

AOI21xp5_ASAP7_75t_L g4802 ( 
.A1(n_4785),
.A2(n_3512),
.B(n_3891),
.Y(n_4802)
);

INVx1_ASAP7_75t_L g4803 ( 
.A(n_4795),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_SL g4804 ( 
.A(n_4798),
.B(n_4794),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4797),
.B(n_4784),
.Y(n_4805)
);

NAND3x1_ASAP7_75t_L g4806 ( 
.A(n_4805),
.B(n_4800),
.C(n_4787),
.Y(n_4806)
);

AOI221xp5_ASAP7_75t_L g4807 ( 
.A1(n_4804),
.A2(n_4796),
.B1(n_4803),
.B2(n_4788),
.C(n_4801),
.Y(n_4807)
);

NOR2x1_ASAP7_75t_L g4808 ( 
.A(n_4804),
.B(n_4790),
.Y(n_4808)
);

INVx1_ASAP7_75t_L g4809 ( 
.A(n_4808),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4809),
.Y(n_4810)
);

NOR3xp33_ASAP7_75t_L g4811 ( 
.A(n_4810),
.B(n_4807),
.C(n_4806),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4811),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_4812),
.Y(n_4813)
);

AOI22xp5_ASAP7_75t_L g4814 ( 
.A1(n_4813),
.A2(n_4789),
.B1(n_4802),
.B2(n_4799),
.Y(n_4814)
);

OR2x6_ASAP7_75t_L g4815 ( 
.A(n_4814),
.B(n_3783),
.Y(n_4815)
);

AOI322xp5_ASAP7_75t_L g4816 ( 
.A1(n_4815),
.A2(n_3705),
.A3(n_3813),
.B1(n_3826),
.B2(n_3902),
.C1(n_3924),
.C2(n_4229),
.Y(n_4816)
);

AOI221xp5_ASAP7_75t_L g4817 ( 
.A1(n_4816),
.A2(n_3783),
.B1(n_3798),
.B2(n_3797),
.C(n_3716),
.Y(n_4817)
);

AOI211xp5_ASAP7_75t_L g4818 ( 
.A1(n_4817),
.A2(n_3798),
.B(n_3797),
.C(n_4082),
.Y(n_4818)
);


endmodule