module fake_netlist_5_551_n_111 (n_16, n_0, n_12, n_9, n_18, n_1, n_8, n_10, n_4, n_11, n_17, n_19, n_7, n_15, n_5, n_14, n_2, n_13, n_3, n_6, n_111);

input n_16;
input n_0;
input n_12;
input n_9;
input n_18;
input n_1;
input n_8;
input n_10;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_5;
input n_14;
input n_2;
input n_13;
input n_3;
input n_6;

output n_111;

wire n_91;
wire n_82;
wire n_24;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_96;
wire n_37;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_42;
wire n_22;
wire n_45;
wire n_46;
wire n_21;
wire n_94;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_30;
wire n_33;
wire n_84;
wire n_23;
wire n_29;
wire n_79;
wire n_47;
wire n_25;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_85;
wire n_95;
wire n_59;
wire n_26;
wire n_55;
wire n_99;
wire n_49;
wire n_20;
wire n_39;
wire n_54;
wire n_67;
wire n_36;
wire n_76;
wire n_87;
wire n_27;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_28;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVxp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_26),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_20),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2x1p5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_31),
.Y(n_57)
);

NAND2x1p5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_23),
.Y(n_58)
);

AND2x4_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_53),
.A2(n_48),
.B1(n_46),
.B2(n_41),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_41),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_43),
.B(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_47),
.B1(n_42),
.B2(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

OAI21x1_ASAP7_75t_L g65 ( 
.A1(n_62),
.A2(n_57),
.B(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_57),
.B(n_42),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_37),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_SL g69 ( 
.A(n_63),
.B(n_30),
.C(n_21),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_69),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g71 ( 
.A(n_69),
.B(n_60),
.C(n_32),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_R g73 ( 
.A(n_64),
.B(n_16),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_60),
.Y(n_74)
);

OAI221xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_66),
.B1(n_64),
.B2(n_67),
.C(n_28),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_68),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_68),
.B1(n_67),
.B2(n_65),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_77),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_70),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_74),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AO21x2_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_73),
.B(n_65),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_72),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_85),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_27),
.B1(n_25),
.B2(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_88),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_83),
.B(n_92),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_90),
.B(n_87),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_87),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_95),
.B(n_96),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_91),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_6),
.C2(n_7),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_68),
.B1(n_56),
.B2(n_55),
.Y(n_100)
);

OAI211xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_47),
.B(n_4),
.C(n_6),
.Y(n_101)
);

AOI311xp33_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_0),
.A3(n_7),
.B(n_56),
.C(n_55),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_0),
.Y(n_103)
);

NAND4xp75_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_37),
.C(n_15),
.D(n_14),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_103),
.Y(n_105)
);

OAI22x1_ASAP7_75t_SL g106 ( 
.A1(n_102),
.A2(n_101),
.B1(n_57),
.B2(n_65),
.Y(n_106)
);

AOI21x1_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_104),
.B(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_107),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_109),
.A2(n_106),
.B1(n_52),
.B2(n_49),
.Y(n_110)
);

O2A1O1Ixp33_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_49),
.B(n_108),
.C(n_109),
.Y(n_111)
);


endmodule