module fake_netlist_6_3620_n_1803 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1803);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1803;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g163 ( 
.A(n_27),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_80),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_12),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_16),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_10),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_23),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_72),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_49),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_128),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_90),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_32),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_112),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_0),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_98),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_73),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_105),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_15),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_34),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_17),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_115),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_117),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_48),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_129),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_42),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_82),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_103),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_30),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_62),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_28),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_48),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_47),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_135),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_89),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_100),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_107),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_38),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_7),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_19),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_119),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_70),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_88),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_87),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_124),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_33),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_65),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_150),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_141),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_32),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_93),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_54),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_154),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_137),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_153),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_76),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_113),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_56),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_51),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_24),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_125),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_39),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_61),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_54),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_39),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_38),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_147),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_30),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_50),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_121),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_37),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_8),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_151),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_96),
.Y(n_263)
);

BUFx10_ASAP7_75t_L g264 ( 
.A(n_51),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_116),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_22),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_43),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_114),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_15),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_69),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_41),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_42),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_11),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_155),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_0),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_49),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_66),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_11),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_59),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_52),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_19),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_74),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_12),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_13),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_81),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_71),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_132),
.Y(n_292)
);

BUFx8_ASAP7_75t_SL g293 ( 
.A(n_143),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_111),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_92),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_14),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_63),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_25),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_45),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_79),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_83),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_29),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_148),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_58),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_123),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_44),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_16),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_35),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_46),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_14),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_94),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_146),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_6),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_106),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_24),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_43),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_1),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_134),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_4),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_126),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_157),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_244),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_178),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_286),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_320),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_194),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_194),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_194),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_194),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_293),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_194),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_230),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_237),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_165),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_203),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_230),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_165),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_208),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_170),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_230),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_209),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_170),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_212),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_219),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_220),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_277),
.Y(n_350)
);

INVxp33_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_230),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_256),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_226),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_277),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_282),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_241),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_229),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_179),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_179),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_282),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_197),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_234),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_232),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_163),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_232),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_184),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_198),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_163),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_210),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_213),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_235),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_215),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_240),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_238),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_176),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_257),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_176),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_284),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_242),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_245),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_246),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_307),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_308),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_247),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_250),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_262),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_266),
.Y(n_394)
);

INVxp33_ASAP7_75t_SL g395 ( 
.A(n_168),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_292),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_172),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_172),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_295),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_297),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_302),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_328),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_329),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_337),
.B(n_173),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_325),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_173),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_324),
.A2(n_254),
.B1(n_190),
.B2(n_189),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_330),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_379),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_357),
.B(n_360),
.C(n_359),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_265),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_327),
.Y(n_420)
);

INVx2_ASAP7_75t_SL g421 ( 
.A(n_361),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_363),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g423 ( 
.A1(n_338),
.A2(n_188),
.B(n_186),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_333),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_343),
.B(n_186),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_333),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_368),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_345),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_347),
.B(n_188),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_377),
.B(n_253),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_342),
.B(n_222),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_348),
.B(n_222),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_369),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_373),
.B(n_195),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_375),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_352),
.B(n_175),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_366),
.B(n_169),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_370),
.A2(n_276),
.B1(n_291),
.B2(n_288),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_363),
.B(n_183),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_326),
.A2(n_171),
.B1(n_315),
.B2(n_312),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_336),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_336),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_381),
.B(n_382),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_351),
.A2(n_190),
.B1(n_189),
.B2(n_174),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_395),
.A2(n_268),
.B1(n_315),
.B2(n_312),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_354),
.A2(n_168),
.B1(n_311),
.B2(n_309),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_339),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_392),
.B(n_227),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_394),
.B(n_205),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_365),
.B(n_206),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_399),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_371),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_372),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_339),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_367),
.B(n_253),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_400),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_401),
.B(n_358),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_341),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_372),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_367),
.B(n_171),
.Y(n_469)
);

INVx5_ASAP7_75t_L g470 ( 
.A(n_341),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_344),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_397),
.B(n_207),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_344),
.B(n_191),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_332),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_439),
.B(n_364),
.Y(n_479)
);

AO21x2_ASAP7_75t_L g480 ( 
.A1(n_458),
.A2(n_217),
.B(n_216),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_457),
.B(n_384),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_456),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_411),
.B(n_388),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_450),
.B(n_396),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_405),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_450),
.B(n_169),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_174),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_420),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_431),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_431),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_450),
.B(n_429),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_438),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_438),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_397),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_378),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_435),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_407),
.B(n_398),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_435),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_442),
.A2(n_275),
.B1(n_182),
.B2(n_322),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_409),
.B(n_263),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_435),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_406),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_427),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_402),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_417),
.Y(n_515)
);

OAI21xp33_ASAP7_75t_SL g516 ( 
.A1(n_433),
.A2(n_423),
.B(n_425),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_427),
.Y(n_517)
);

INVxp67_ASAP7_75t_R g518 ( 
.A(n_443),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_402),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_454),
.B(n_453),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_432),
.B(n_398),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_433),
.B(n_346),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_436),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_450),
.B(n_169),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_447),
.Y(n_526)
);

INVxp33_ASAP7_75t_L g527 ( 
.A(n_451),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_422),
.B(n_230),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_447),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_440),
.B(n_374),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_447),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_410),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_460),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_417),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_403),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_447),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_441),
.B(n_285),
.Y(n_540)
);

CKINVDCx6p67_ASAP7_75t_R g541 ( 
.A(n_410),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_403),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_419),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_230),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_441),
.B(n_323),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_412),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_469),
.B(n_214),
.C(n_211),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_412),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_441),
.B(n_218),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_444),
.B(n_349),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_465),
.A2(n_466),
.B1(n_443),
.B2(n_451),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_414),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_441),
.B(n_224),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_444),
.B(n_228),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_444),
.B(n_231),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g556 ( 
.A(n_426),
.Y(n_556)
);

BUFx6f_ASAP7_75t_SL g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_414),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_426),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_447),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_L g561 ( 
.A(n_464),
.B(n_230),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_447),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_459),
.B(n_374),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_459),
.B(n_259),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_455),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_455),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_455),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_464),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

BUFx10_ASAP7_75t_L g571 ( 
.A(n_475),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_424),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_455),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_424),
.Y(n_574)
);

BUFx10_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_459),
.B(n_271),
.Y(n_576)
);

BUFx6f_ASAP7_75t_SL g577 ( 
.A(n_456),
.Y(n_577)
);

CKINVDCx14_ASAP7_75t_R g578 ( 
.A(n_445),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_419),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_428),
.Y(n_580)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_445),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_428),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_421),
.B(n_204),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_434),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_416),
.B(n_187),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_455),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_427),
.B(n_289),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_427),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_437),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_437),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_449),
.A2(n_393),
.B1(n_391),
.B2(n_390),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_L g593 ( 
.A(n_421),
.B(n_230),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_449),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_413),
.B(n_290),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_463),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_452),
.B(n_349),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_452),
.Y(n_599)
);

AOI21x1_ASAP7_75t_L g600 ( 
.A1(n_473),
.A2(n_462),
.B(n_461),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_413),
.B(n_294),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_413),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_463),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_461),
.B(n_164),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_473),
.B(n_187),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_462),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_463),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_468),
.A2(n_393),
.B1(n_391),
.B2(n_390),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_468),
.B(n_376),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_474),
.B(n_187),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_463),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_413),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_463),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_413),
.B(n_301),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_471),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_446),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_R g618 ( 
.A(n_471),
.B(n_164),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_471),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_446),
.B(n_196),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_413),
.B(n_304),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_471),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_467),
.B(n_196),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_470),
.B(n_305),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_471),
.B(n_166),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_470),
.B(n_306),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_501),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_523),
.B(n_471),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_523),
.B(n_166),
.Y(n_629)
);

AO221x1_ASAP7_75t_L g630 ( 
.A1(n_594),
.A2(n_313),
.B1(n_314),
.B2(n_387),
.C(n_386),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_501),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_569),
.B(n_252),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_509),
.B(n_167),
.Y(n_633)
);

AOI21x1_ASAP7_75t_L g634 ( 
.A1(n_600),
.A2(n_467),
.B(n_356),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_504),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_504),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_507),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_569),
.B(n_474),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_516),
.B(n_252),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_595),
.B(n_252),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_595),
.B(n_252),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_479),
.B(n_167),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_595),
.B(n_252),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_483),
.B(n_536),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_515),
.B(n_474),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_507),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_510),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_563),
.B(n_376),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_617),
.B(n_580),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_617),
.B(n_474),
.Y(n_650)
);

OR2x6_ASAP7_75t_L g651 ( 
.A(n_500),
.B(n_380),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_510),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_580),
.B(n_582),
.Y(n_653)
);

NAND2x1_ASAP7_75t_L g654 ( 
.A(n_495),
.B(n_524),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_582),
.B(n_474),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_584),
.B(n_474),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_499),
.B(n_255),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_538),
.B(n_252),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_481),
.B(n_177),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_513),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_478),
.B(n_177),
.Y(n_661)
);

NOR2x1p5_ASAP7_75t_L g662 ( 
.A(n_541),
.B(n_201),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_480),
.A2(n_561),
.B1(n_563),
.B2(n_550),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_478),
.B(n_180),
.Y(n_664)
);

AND2x4_ASAP7_75t_SL g665 ( 
.A(n_571),
.B(n_163),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_482),
.B(n_180),
.Y(n_666)
);

AND2x2_ASAP7_75t_SL g667 ( 
.A(n_561),
.B(n_380),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_584),
.B(n_587),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_480),
.A2(n_563),
.B1(n_550),
.B2(n_587),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_513),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_520),
.A2(n_298),
.B1(n_387),
.B2(n_386),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_R g672 ( 
.A(n_533),
.B(n_181),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_519),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_590),
.B(n_591),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_519),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_590),
.B(n_470),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_499),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_591),
.B(n_470),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_SL g679 ( 
.A(n_520),
.B(n_201),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_538),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_484),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_599),
.A2(n_185),
.B1(n_182),
.B2(n_192),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_482),
.B(n_181),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_538),
.B(n_252),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_583),
.B(n_264),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_607),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_599),
.B(n_185),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_607),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_505),
.B(n_470),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_521),
.B(n_470),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_598),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_538),
.B(n_252),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_522),
.B(n_192),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_535),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_522),
.B(n_193),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_538),
.B(n_193),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_575),
.B(n_199),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_583),
.B(n_264),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_575),
.B(n_199),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_535),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_542),
.Y(n_701)
);

OR2x6_ASAP7_75t_L g702 ( 
.A(n_500),
.B(n_383),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_575),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_614),
.B(n_200),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_610),
.B(n_383),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_598),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_614),
.B(n_200),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_542),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_546),
.B(n_202),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_600),
.B(n_202),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_546),
.B(n_243),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_541),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_548),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_548),
.B(n_243),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_500),
.B(n_269),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_552),
.Y(n_716)
);

AOI22x1_ASAP7_75t_L g717 ( 
.A1(n_552),
.A2(n_279),
.B1(n_269),
.B2(n_275),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_558),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_533),
.B(n_278),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_530),
.B(n_264),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_503),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_530),
.B(n_385),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_558),
.Y(n_723)
);

HB1xp67_ASAP7_75t_L g724 ( 
.A(n_484),
.Y(n_724)
);

AND2x6_ASAP7_75t_SL g725 ( 
.A(n_530),
.B(n_385),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_572),
.B(n_278),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_571),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_572),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_500),
.B(n_279),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_574),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_574),
.Y(n_731)
);

BUFx8_ASAP7_75t_L g732 ( 
.A(n_559),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_578),
.B(n_221),
.C(n_223),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_495),
.B(n_281),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_619),
.A2(n_322),
.B(n_316),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_619),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_540),
.A2(n_281),
.B1(n_316),
.B2(n_236),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_610),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_610),
.Y(n_739)
);

AOI221xp5_ASAP7_75t_L g740 ( 
.A1(n_581),
.A2(n_276),
.B1(n_270),
.B2(n_273),
.C(n_274),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_604),
.B(n_225),
.C(n_233),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_545),
.B(n_239),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_557),
.A2(n_248),
.B1(n_249),
.B2(n_251),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_495),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_480),
.B(n_258),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_524),
.B(n_534),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_524),
.B(n_260),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_557),
.A2(n_261),
.B1(n_267),
.B2(n_287),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_SL g749 ( 
.A(n_496),
.B(n_270),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_549),
.A2(n_273),
.B1(n_274),
.B2(n_280),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_553),
.A2(n_280),
.B1(n_283),
.B2(n_288),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_534),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_476),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_476),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_534),
.B(n_299),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_492),
.B(n_303),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_477),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_488),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_503),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_537),
.B(n_300),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_488),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_554),
.A2(n_311),
.B1(n_291),
.B2(n_309),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_537),
.B(n_362),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_571),
.Y(n_764)
);

BUFx6f_ASAP7_75t_SL g765 ( 
.A(n_530),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_490),
.Y(n_766)
);

O2A1O1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_528),
.A2(n_362),
.B(n_356),
.C(n_355),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_537),
.B(n_355),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_543),
.B(n_350),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_543),
.B(n_350),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_508),
.B(n_283),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_543),
.B(n_162),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_490),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_567),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_477),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_623),
.B(n_159),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_SL g777 ( 
.A(n_551),
.B(n_527),
.C(n_532),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_567),
.B(n_152),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_567),
.B(n_149),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_555),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_620),
.B(n_3),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_487),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_487),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_564),
.B(n_145),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_492),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_613),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_576),
.B(n_142),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_502),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_506),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_620),
.B(n_5),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_502),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_559),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_493),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_526),
.B(n_140),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_547),
.B(n_139),
.Y(n_795)
);

OAI22xp33_ASAP7_75t_L g796 ( 
.A1(n_489),
.A2(n_8),
.B1(n_9),
.B2(n_17),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_525),
.B(n_9),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_486),
.B(n_18),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_667),
.A2(n_557),
.B1(n_577),
.B2(n_593),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_721),
.B(n_556),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_738),
.B(n_585),
.Y(n_801)
);

AND3x1_ASAP7_75t_SL g802 ( 
.A(n_740),
.B(n_491),
.C(n_518),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_667),
.B(n_526),
.Y(n_803)
);

NAND2x1p5_ASAP7_75t_L g804 ( 
.A(n_736),
.B(n_589),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_636),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_652),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_679),
.A2(n_528),
.B1(n_544),
.B2(n_491),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_652),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_633),
.B(n_579),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_627),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_792),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_721),
.B(n_759),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_649),
.B(n_579),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_669),
.B(n_529),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_686),
.B(n_493),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_785),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_759),
.B(n_577),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_629),
.B(n_577),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_792),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_660),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_685),
.B(n_518),
.Y(n_821)
);

INVx5_ASAP7_75t_L g822 ( 
.A(n_680),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_688),
.B(n_494),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_663),
.B(n_529),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_785),
.B(n_544),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_631),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_736),
.B(n_744),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_660),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_670),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_786),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_713),
.B(n_494),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_716),
.B(n_497),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_786),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_677),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_698),
.B(n_485),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_670),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_727),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_635),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_718),
.B(n_497),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_730),
.B(n_498),
.Y(n_840)
);

OR2x2_ASAP7_75t_L g841 ( 
.A(n_657),
.B(n_681),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_736),
.B(n_531),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_637),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_673),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_724),
.B(n_693),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_744),
.B(n_531),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_687),
.B(n_777),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_722),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_646),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_731),
.B(n_498),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_647),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_673),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_675),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_653),
.B(n_589),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_668),
.B(n_602),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_675),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_SL g857 ( 
.A(n_771),
.B(n_485),
.C(n_606),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_744),
.B(n_539),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_679),
.A2(n_593),
.B1(n_514),
.B2(n_511),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_752),
.B(n_539),
.Y(n_860)
);

INVx5_ASAP7_75t_L g861 ( 
.A(n_680),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_674),
.B(n_602),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_SL g863 ( 
.A1(n_781),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_694),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_694),
.B(n_602),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_700),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_672),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_739),
.B(n_611),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_700),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_701),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_701),
.Y(n_871)
);

INVx1_ASAP7_75t_SL g872 ( 
.A(n_756),
.Y(n_872)
);

AND3x2_ASAP7_75t_SL g873 ( 
.A(n_796),
.B(n_20),
.C(n_21),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_720),
.Y(n_874)
);

AOI21xp33_ASAP7_75t_L g875 ( 
.A1(n_642),
.A2(n_625),
.B(n_588),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_708),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_786),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_705),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_708),
.B(n_613),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_723),
.B(n_728),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_723),
.B(n_612),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_728),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_789),
.A2(n_506),
.B(n_512),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_756),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_789),
.A2(n_506),
.B(n_512),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_741),
.B(n_596),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_758),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_786),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_628),
.B(n_622),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_659),
.B(n_622),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_752),
.B(n_608),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_761),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_651),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_671),
.A2(n_511),
.B1(n_514),
.B2(n_605),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_766),
.Y(n_895)
);

BUFx4f_ASAP7_75t_L g896 ( 
.A(n_776),
.Y(n_896)
);

BUFx4f_ASAP7_75t_L g897 ( 
.A(n_776),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_773),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_691),
.B(n_612),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_706),
.B(n_592),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_793),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_703),
.Y(n_902)
);

OR2x6_ASAP7_75t_L g903 ( 
.A(n_727),
.B(n_601),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_661),
.B(n_597),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_705),
.Y(n_905)
);

NOR2x1p5_ASAP7_75t_L g906 ( 
.A(n_764),
.B(n_621),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_752),
.B(n_586),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_671),
.A2(n_798),
.B1(n_797),
.B2(n_790),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_774),
.B(n_586),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_753),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_671),
.A2(n_597),
.B1(n_560),
.B2(n_562),
.Y(n_911)
);

AND2x6_ASAP7_75t_SL g912 ( 
.A(n_715),
.B(n_615),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_754),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_651),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_634),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_664),
.B(n_573),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_666),
.B(n_573),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_754),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_774),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_696),
.A2(n_570),
.B1(n_560),
.B2(n_562),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_705),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_SL g922 ( 
.A1(n_665),
.A2(n_618),
.B1(n_565),
.B2(n_603),
.Y(n_922)
);

AOI211xp5_ASAP7_75t_L g923 ( 
.A1(n_729),
.A2(n_626),
.B(n_624),
.C(n_616),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_680),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_695),
.B(n_609),
.Y(n_925)
);

BUFx2_ASAP7_75t_SL g926 ( 
.A(n_764),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_SL g927 ( 
.A(n_682),
.B(n_22),
.C(n_23),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_648),
.B(n_703),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_654),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_683),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_732),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_757),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_775),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_774),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_712),
.B(n_78),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_SL g936 ( 
.A1(n_712),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_789),
.A2(n_512),
.B(n_517),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_648),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_742),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_648),
.B(n_616),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_696),
.A2(n_608),
.B(n_605),
.C(n_603),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_704),
.B(n_517),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_760),
.A2(n_570),
.B1(n_568),
.B2(n_566),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_780),
.A2(n_568),
.B(n_566),
.C(n_565),
.Y(n_944)
);

AND2x6_ASAP7_75t_L g945 ( 
.A(n_776),
.B(n_57),
.Y(n_945)
);

OR2x2_ASAP7_75t_SL g946 ( 
.A(n_745),
.B(n_26),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_784),
.B(n_517),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_719),
.B(n_29),
.Y(n_948)
);

AND2x6_ASAP7_75t_L g949 ( 
.A(n_772),
.B(n_60),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_782),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_782),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_780),
.A2(n_31),
.B(n_34),
.C(n_35),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_707),
.B(n_31),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_783),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_672),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_665),
.B(n_40),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_732),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_783),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_788),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_651),
.B(n_40),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_732),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_630),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_962)
);

INVx5_ASAP7_75t_L g963 ( 
.A(n_651),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_702),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_638),
.B(n_47),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_644),
.B(n_50),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_709),
.B(n_53),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_791),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_702),
.B(n_53),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_788),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_778),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_791),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_791),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_763),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_768),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_746),
.Y(n_976)
);

INVx4_ASAP7_75t_L g977 ( 
.A(n_702),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_769),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_770),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_SL g980 ( 
.A(n_733),
.B(n_55),
.C(n_64),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_702),
.B(n_762),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_765),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_779),
.A2(n_68),
.B1(n_84),
.B2(n_86),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_655),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_711),
.B(n_91),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_725),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_656),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_939),
.B(n_726),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_847),
.A2(n_697),
.B1(n_699),
.B2(n_749),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_847),
.B(n_714),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_807),
.A2(n_699),
.B1(n_697),
.B2(n_710),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_908),
.A2(n_750),
.B(n_751),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_925),
.B(n_755),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_947),
.A2(n_645),
.B(n_692),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_805),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_806),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_947),
.A2(n_692),
.B(n_658),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_930),
.B(n_743),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_830),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_807),
.A2(n_897),
.B1(n_896),
.B2(n_890),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_900),
.B(n_747),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_808),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_SL g1003 ( 
.A1(n_985),
.A2(n_787),
.B(n_767),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_824),
.A2(n_942),
.B(n_814),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_818),
.B(n_748),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_890),
.B(n_760),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_818),
.B(n_737),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_974),
.B(n_734),
.Y(n_1008)
);

AOI22xp33_ASAP7_75t_SL g1009 ( 
.A1(n_821),
.A2(n_765),
.B1(n_717),
.B2(n_662),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_800),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_841),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_908),
.A2(n_779),
.B1(n_632),
.B2(n_795),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_978),
.B(n_734),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_R g1014 ( 
.A(n_816),
.B(n_765),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_824),
.A2(n_684),
.B(n_658),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_967),
.A2(n_632),
.B(n_641),
.C(n_640),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_828),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_942),
.A2(n_684),
.B(n_710),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_810),
.B(n_641),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_828),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_814),
.A2(n_650),
.B(n_639),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_848),
.B(n_640),
.Y(n_1022)
);

O2A1O1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_953),
.A2(n_643),
.B(n_639),
.C(n_735),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_829),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_829),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_830),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_811),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_830),
.Y(n_1028)
);

AOI33xp33_ASAP7_75t_L g1029 ( 
.A1(n_962),
.A2(n_643),
.A3(n_794),
.B1(n_690),
.B2(n_689),
.B3(n_676),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_811),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_854),
.A2(n_794),
.B(n_678),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_928),
.B(n_825),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_848),
.B(n_99),
.Y(n_1033)
);

AO21x2_ASAP7_75t_L g1034 ( 
.A1(n_944),
.A2(n_875),
.B(n_965),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_837),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_967),
.A2(n_109),
.B(n_118),
.C(n_120),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_845),
.B(n_133),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_857),
.A2(n_138),
.B(n_952),
.C(n_966),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_896),
.A2(n_897),
.B1(n_799),
.B2(n_809),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_836),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_819),
.Y(n_1041)
);

AND2x6_ASAP7_75t_L g1042 ( 
.A(n_971),
.B(n_915),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_836),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_826),
.B(n_838),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_928),
.B(n_825),
.Y(n_1045)
);

BUFx4_ASAP7_75t_SL g1046 ( 
.A(n_957),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_844),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_843),
.B(n_849),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_867),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_938),
.B(n_878),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_962),
.A2(n_945),
.B1(n_983),
.B2(n_980),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_955),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_834),
.B(n_812),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_883),
.A2(n_937),
.B(n_885),
.Y(n_1054)
);

OAI21xp33_ASAP7_75t_SL g1055 ( 
.A1(n_851),
.A2(n_859),
.B(n_887),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_987),
.B(n_984),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_952),
.A2(n_874),
.B(n_927),
.C(n_944),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_987),
.B(n_975),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_868),
.A2(n_801),
.B(n_817),
.C(n_895),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_876),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_819),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_880),
.A2(n_859),
.B1(n_963),
.B2(n_934),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_975),
.B(n_979),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_855),
.A2(n_862),
.B(n_904),
.Y(n_1064)
);

OAI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_835),
.A2(n_817),
.B(n_884),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_977),
.B(n_905),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_876),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_882),
.Y(n_1068)
);

CKINVDCx14_ASAP7_75t_R g1069 ( 
.A(n_935),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_882),
.Y(n_1070)
);

OAI22x1_ASAP7_75t_L g1071 ( 
.A1(n_981),
.A2(n_964),
.B1(n_893),
.B2(n_914),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_916),
.A2(n_917),
.B(n_889),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_872),
.B(n_892),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_898),
.B(n_901),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_921),
.B(n_912),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_927),
.A2(n_948),
.B(n_899),
.C(n_960),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_827),
.A2(n_803),
.B(n_879),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_893),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_827),
.A2(n_803),
.B(n_979),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_933),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_977),
.B(n_914),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_976),
.B(n_852),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_933),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_954),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_801),
.A2(n_956),
.B(n_894),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_868),
.A2(n_886),
.B(n_976),
.C(n_871),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_853),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_963),
.A2(n_934),
.B1(n_919),
.B2(n_870),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_982),
.Y(n_1089)
);

BUFx12f_ASAP7_75t_L g1090 ( 
.A(n_931),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_R g1091 ( 
.A(n_837),
.B(n_902),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_SL g1092 ( 
.A(n_936),
.B(n_873),
.C(n_940),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_964),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_963),
.B(n_902),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_856),
.B(n_864),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_815),
.A2(n_850),
.B(n_839),
.C(n_832),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_866),
.B(n_820),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_813),
.B(n_869),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_941),
.A2(n_923),
.B(n_911),
.C(n_831),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_894),
.B(n_840),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_954),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_913),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_911),
.A2(n_823),
.B(n_983),
.C(n_943),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_919),
.A2(n_920),
.B(n_950),
.C(n_918),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_963),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_830),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_961),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_945),
.A2(n_969),
.B1(n_949),
.B2(n_959),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_958),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_910),
.B(n_970),
.Y(n_1110)
);

OAI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_969),
.A2(n_873),
.B1(n_902),
.B2(n_903),
.Y(n_1111)
);

NOR2x1_ASAP7_75t_L g1112 ( 
.A(n_926),
.B(n_877),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_932),
.B(n_951),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_945),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_822),
.A2(n_924),
.B1(n_861),
.B2(n_804),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_906),
.B(n_902),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_986),
.B(n_946),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_SL g1118 ( 
.A(n_945),
.B(n_877),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_945),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_915),
.A2(n_842),
.B(n_881),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_922),
.B(n_804),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_842),
.A2(n_909),
.B(n_891),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_972),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_846),
.A2(n_907),
.B(n_891),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_968),
.A2(n_971),
.B1(n_833),
.B2(n_888),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_863),
.B(n_903),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_SL g1127 ( 
.A(n_935),
.B(n_971),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_846),
.A2(n_909),
.B(n_858),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_949),
.A2(n_973),
.B1(n_972),
.B2(n_860),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_865),
.A2(n_907),
.B(n_858),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_860),
.A2(n_971),
.B(n_929),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_903),
.B(n_929),
.Y(n_1132)
);

AO32x1_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_948),
.A3(n_523),
.B1(n_670),
.B2(n_673),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_929),
.A2(n_949),
.B(n_802),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1001),
.B(n_929),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_SL g1136 ( 
.A1(n_991),
.A2(n_802),
.B(n_949),
.C(n_1007),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1044),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_989),
.A2(n_992),
.B(n_1006),
.C(n_1038),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1048),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1102),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_1091),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_988),
.B(n_1073),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_L g1144 ( 
.A1(n_1111),
.A2(n_1051),
.B1(n_1092),
.B2(n_1000),
.C(n_1057),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_1021),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1072),
.A2(n_1064),
.B(n_1096),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1051),
.A2(n_1012),
.B(n_1008),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_SL g1148 ( 
.A(n_1089),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_990),
.A2(n_1005),
.B(n_998),
.C(n_1059),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1030),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1063),
.B(n_1056),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_994),
.A2(n_997),
.B(n_1016),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1058),
.B(n_993),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1076),
.A2(n_1037),
.B(n_1103),
.C(n_1012),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1124),
.A2(n_1122),
.B(n_1015),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1081),
.B(n_1116),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1079),
.A2(n_1077),
.B(n_1120),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1100),
.B(n_1022),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_1126),
.A2(n_1073),
.B1(n_1117),
.B2(n_1093),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_1041),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1130),
.A2(n_1031),
.B(n_1062),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1022),
.B(n_1074),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1003),
.A2(n_1099),
.B(n_1023),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_R g1165 ( 
.A(n_1090),
.B(n_1107),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1011),
.B(n_1010),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1032),
.B(n_1045),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1010),
.B(n_1011),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1134),
.A2(n_1115),
.B(n_1125),
.Y(n_1169)
);

BUFx4f_ASAP7_75t_SL g1170 ( 
.A(n_1035),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1039),
.A2(n_1086),
.B(n_1118),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1065),
.A2(n_1111),
.B(n_1092),
.C(n_1121),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1055),
.A2(n_1104),
.B(n_1129),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1074),
.B(n_1085),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1061),
.B(n_1041),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1034),
.A2(n_1019),
.B(n_1129),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_995),
.Y(n_1177)
);

AOI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1037),
.A2(n_1117),
.B1(n_1075),
.B2(n_1127),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1088),
.A2(n_1113),
.B(n_1082),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1029),
.A2(n_1097),
.B(n_1095),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_1114),
.B(n_1119),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_1112),
.B(n_1094),
.Y(n_1182)
);

BUFx10_ASAP7_75t_L g1183 ( 
.A(n_1049),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1036),
.A2(n_1093),
.B(n_1078),
.C(n_1075),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1053),
.B(n_1078),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1053),
.B(n_1052),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_SL g1187 ( 
.A1(n_1110),
.A2(n_1060),
.B(n_1105),
.C(n_1132),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_996),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1097),
.A2(n_1095),
.B(n_1033),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1034),
.A2(n_1133),
.B(n_1108),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1002),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1069),
.B(n_1033),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1026),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1020),
.B(n_1070),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1009),
.A2(n_1132),
.B1(n_1071),
.B2(n_1050),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1024),
.B(n_1043),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1025),
.B(n_1047),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1040),
.B(n_1068),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1123),
.A2(n_1083),
.B(n_1109),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1026),
.A2(n_1028),
.B(n_1066),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1081),
.B(n_1027),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1133),
.A2(n_1108),
.B(n_1066),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1087),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1067),
.A2(n_1084),
.B(n_1101),
.C(n_1080),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1091),
.B(n_1014),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_999),
.A2(n_1105),
.B(n_1106),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_999),
.A2(n_1106),
.B(n_1042),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1026),
.Y(n_1208)
);

O2A1O1Ixp5_ASAP7_75t_L g1209 ( 
.A1(n_1042),
.A2(n_1026),
.B(n_1028),
.C(n_1014),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1042),
.B(n_1028),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1089),
.B(n_1028),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1042),
.A2(n_1054),
.B(n_1131),
.Y(n_1212)
);

NAND3xp33_ASAP7_75t_SL g1213 ( 
.A(n_1046),
.B(n_908),
.C(n_533),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1046),
.B(n_821),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1010),
.B(n_821),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1061),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_1049),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1030),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1044),
.Y(n_1222)
);

CKINVDCx8_ASAP7_75t_R g1223 ( 
.A(n_1049),
.Y(n_1223)
);

BUFx5_ASAP7_75t_L g1224 ( 
.A(n_1042),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1072),
.A2(n_1018),
.B(n_1004),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_989),
.A2(n_847),
.B(n_798),
.C(n_992),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1010),
.B(n_821),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1065),
.A2(n_857),
.B1(n_327),
.B2(n_324),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1017),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1044),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1030),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1091),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1091),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1112),
.B(n_963),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1061),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1044),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1099),
.A2(n_944),
.A3(n_991),
.B(n_1004),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1044),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1051),
.A2(n_807),
.B1(n_908),
.B2(n_1111),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1244)
);

AND3x4_ASAP7_75t_L g1245 ( 
.A(n_1092),
.B(n_733),
.C(n_727),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_SL g1246 ( 
.A1(n_1051),
.A2(n_857),
.B(n_485),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1011),
.B(n_841),
.Y(n_1247)
);

NAND3xp33_ASAP7_75t_L g1248 ( 
.A(n_989),
.B(n_847),
.C(n_659),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1044),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1072),
.A2(n_1064),
.B(n_1018),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1054),
.A2(n_1131),
.B(n_1128),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1072),
.A2(n_1064),
.B(n_1018),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1032),
.B(n_926),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_1021),
.Y(n_1255)
);

NOR3xp33_ASAP7_75t_L g1256 ( 
.A(n_1005),
.B(n_857),
.C(n_481),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1073),
.B(n_930),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_988),
.B(n_324),
.Y(n_1258)
);

HB1xp67_ASAP7_75t_L g1259 ( 
.A(n_1041),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1049),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1099),
.A2(n_944),
.A3(n_991),
.B(n_1004),
.Y(n_1262)
);

AOI211x1_ASAP7_75t_L g1263 ( 
.A1(n_992),
.A2(n_1111),
.B(n_796),
.C(n_1085),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1010),
.B(n_821),
.Y(n_1264)
);

AOI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1018),
.A2(n_1004),
.B(n_1021),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1017),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_1099),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_992),
.A2(n_857),
.B1(n_847),
.B2(n_798),
.Y(n_1270)
);

NOR4xp25_ASAP7_75t_L g1271 ( 
.A(n_992),
.B(n_908),
.C(n_1111),
.D(n_1038),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1272)
);

OAI22x1_ASAP7_75t_L g1273 ( 
.A1(n_989),
.A2(n_491),
.B1(n_847),
.B2(n_551),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_1021),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1026),
.Y(n_1275)
);

A2O1A1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_989),
.A2(n_847),
.B(n_798),
.C(n_992),
.Y(n_1276)
);

BUFx3_ASAP7_75t_L g1277 ( 
.A(n_1030),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1017),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1004),
.A2(n_1018),
.B(n_1021),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1001),
.B(n_1063),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1072),
.A2(n_1064),
.B(n_1018),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1051),
.A2(n_857),
.B(n_485),
.Y(n_1283)
);

INVx3_ASAP7_75t_SL g1284 ( 
.A(n_1217),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1199),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1248),
.A2(n_1276),
.B(n_1226),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1164),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1221),
.A2(n_1235),
.B(n_1234),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1142),
.B(n_1232),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1138),
.A2(n_1149),
.B(n_1154),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1238),
.A2(n_1251),
.B(n_1244),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1215),
.B(n_1227),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1143),
.B(n_1246),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1193),
.Y(n_1294)
);

AOI222xp33_ASAP7_75t_L g1295 ( 
.A1(n_1273),
.A2(n_1283),
.B1(n_1243),
.B2(n_1144),
.C1(n_1213),
.C2(n_1270),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1243),
.A2(n_1144),
.B1(n_1256),
.B2(n_1147),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1167),
.B(n_1156),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1158),
.A2(n_1155),
.B(n_1265),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1146),
.A2(n_1253),
.B(n_1282),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1178),
.A2(n_1163),
.B1(n_1228),
.B2(n_1258),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1250),
.A2(n_1225),
.B(n_1152),
.Y(n_1301)
);

BUFx2_ASAP7_75t_SL g1302 ( 
.A(n_1223),
.Y(n_1302)
);

OAI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1189),
.A2(n_1136),
.B(n_1271),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1192),
.A2(n_1189),
.B1(n_1163),
.B2(n_1186),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1162),
.A2(n_1255),
.B(n_1145),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1145),
.A2(n_1255),
.B(n_1280),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1159),
.A2(n_1174),
.B(n_1172),
.C(n_1173),
.Y(n_1307)
);

BUFx3_ASAP7_75t_L g1308 ( 
.A(n_1233),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1247),
.B(n_1175),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1174),
.A2(n_1245),
.B1(n_1159),
.B2(n_1137),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1211),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1167),
.B(n_1156),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1274),
.A2(n_1280),
.B(n_1169),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1264),
.B(n_1185),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1261),
.Y(n_1315)
);

INVx2_ASAP7_75t_SL g1316 ( 
.A(n_1201),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1229),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1216),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1173),
.A2(n_1202),
.B(n_1180),
.Y(n_1319)
);

AO21x2_ASAP7_75t_L g1320 ( 
.A1(n_1180),
.A2(n_1187),
.B(n_1179),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1168),
.Y(n_1321)
);

BUFx4f_ASAP7_75t_SL g1322 ( 
.A(n_1183),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_SL g1323 ( 
.A(n_1170),
.B(n_1205),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1239),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1167),
.B(n_1181),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1268),
.A2(n_1157),
.B(n_1151),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1177),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1207),
.A2(n_1206),
.B(n_1209),
.Y(n_1328)
);

INVx3_ASAP7_75t_SL g1329 ( 
.A(n_1183),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1266),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1150),
.Y(n_1331)
);

NOR2x1_ASAP7_75t_R g1332 ( 
.A(n_1231),
.B(n_1277),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1257),
.A2(n_1184),
.B(n_1166),
.C(n_1249),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1140),
.A2(n_1222),
.B1(n_1230),
.B2(n_1240),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1278),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1242),
.B(n_1272),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1218),
.B(n_1279),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1148),
.Y(n_1338)
);

CKINVDCx11_ASAP7_75t_R g1339 ( 
.A(n_1254),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1210),
.A2(n_1135),
.B(n_1182),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1188),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1157),
.A2(n_1151),
.B(n_1281),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1135),
.A2(n_1204),
.B(n_1279),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1160),
.A2(n_1153),
.A3(n_1218),
.B(n_1281),
.Y(n_1344)
);

INVx4_ASAP7_75t_SL g1345 ( 
.A(n_1254),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1236),
.B(n_1252),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1259),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1148),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1236),
.A2(n_1272),
.B(n_1269),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1219),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1252),
.B(n_1269),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1210),
.A2(n_1182),
.B(n_1237),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1254),
.B(n_1181),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1191),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1260),
.A2(n_1267),
.B(n_1153),
.C(n_1195),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1214),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1237),
.A2(n_1197),
.B(n_1198),
.Y(n_1357)
);

INVx3_ASAP7_75t_SL g1358 ( 
.A(n_1193),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1208),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1260),
.A2(n_1267),
.B(n_1203),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1181),
.Y(n_1361)
);

AO21x2_ASAP7_75t_L g1362 ( 
.A1(n_1194),
.A2(n_1196),
.B(n_1197),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1200),
.A2(n_1196),
.B(n_1198),
.Y(n_1363)
);

A2O1A1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1263),
.A2(n_1161),
.B(n_1241),
.C(n_1262),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1275),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1241),
.B(n_1262),
.Y(n_1366)
);

NAND2x1p5_ASAP7_75t_L g1367 ( 
.A(n_1224),
.B(n_1165),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1241),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1262),
.A2(n_1243),
.B1(n_1283),
.B2(n_1246),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1224),
.A2(n_1212),
.B(n_1139),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1224),
.B(n_1143),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1224),
.B(n_1215),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1224),
.A2(n_1212),
.B(n_1139),
.Y(n_1373)
);

BUFx4f_ASAP7_75t_SL g1374 ( 
.A(n_1183),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1243),
.A2(n_1283),
.B1(n_1246),
.B2(n_1273),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1243),
.A2(n_847),
.B1(n_781),
.B2(n_790),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1143),
.B(n_1163),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1141),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1167),
.B(n_1254),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1212),
.A2(n_1220),
.B(n_1139),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1199),
.Y(n_1381)
);

OAI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1248),
.A2(n_1276),
.B(n_1226),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1190),
.A2(n_1146),
.A3(n_1164),
.B(n_1176),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1141),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1212),
.A2(n_1220),
.B(n_1139),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1199),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1167),
.B(n_1156),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1248),
.B(n_1270),
.C(n_1256),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1199),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1215),
.B(n_1227),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1215),
.B(n_1227),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1167),
.B(n_1156),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1193),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1175),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1141),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1141),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1142),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1224),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1141),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1141),
.Y(n_1400)
);

INVx1_ASAP7_75t_SL g1401 ( 
.A(n_1216),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1141),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1170),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1215),
.B(n_1227),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1212),
.A2(n_1220),
.B(n_1139),
.Y(n_1405)
);

AO31x2_ASAP7_75t_L g1406 ( 
.A1(n_1190),
.A2(n_1146),
.A3(n_1164),
.B(n_1176),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1167),
.B(n_1156),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1143),
.B(n_1163),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1199),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1243),
.A2(n_1273),
.B1(n_992),
.B2(n_1144),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1193),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1141),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1247),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1314),
.B(n_1292),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1377),
.B(n_1408),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1299),
.A2(n_1301),
.B(n_1349),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1331),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1309),
.B(n_1394),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1337),
.B(n_1346),
.Y(n_1419)
);

OAI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1376),
.A2(n_1293),
.B1(n_1410),
.B2(n_1304),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1368),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1360),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1290),
.A2(n_1355),
.B(n_1342),
.Y(n_1423)
);

CKINVDCx6p67_ASAP7_75t_R g1424 ( 
.A(n_1284),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1345),
.B(n_1297),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1300),
.A2(n_1375),
.B(n_1382),
.C(n_1293),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1315),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1375),
.A2(n_1295),
.B(n_1355),
.C(n_1388),
.Y(n_1429)
);

NOR2xp67_ASAP7_75t_R g1430 ( 
.A(n_1315),
.B(n_1331),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1410),
.A2(n_1310),
.B1(n_1296),
.B2(n_1334),
.Y(n_1431)
);

O2A1O1Ixp5_ASAP7_75t_L g1432 ( 
.A1(n_1303),
.A2(n_1287),
.B(n_1369),
.C(n_1326),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1344),
.B(n_1413),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1351),
.B(n_1336),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1331),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1310),
.A2(n_1296),
.B1(n_1334),
.B2(n_1289),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1322),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1321),
.B(n_1404),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1333),
.A2(n_1367),
.B(n_1379),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1371),
.B(n_1324),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1313),
.A2(n_1298),
.B(n_1305),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_L g1442 ( 
.A1(n_1307),
.A2(n_1369),
.B(n_1364),
.C(n_1347),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1367),
.A2(n_1379),
.B(n_1332),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1307),
.B(n_1318),
.Y(n_1444)
);

OAI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1356),
.A2(n_1323),
.B1(n_1397),
.B2(n_1289),
.C(n_1401),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1364),
.A2(n_1316),
.B(n_1379),
.C(n_1402),
.Y(n_1446)
);

OAI22xp5_ASAP7_75t_L g1447 ( 
.A1(n_1308),
.A2(n_1353),
.B1(n_1316),
.B2(n_1392),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1308),
.A2(n_1353),
.B1(n_1407),
.B2(n_1387),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1360),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1327),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1341),
.Y(n_1451)
);

O2A1O1Ixp33_ASAP7_75t_L g1452 ( 
.A1(n_1412),
.A2(n_1378),
.B(n_1384),
.C(n_1354),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1395),
.A2(n_1399),
.B(n_1400),
.C(n_1396),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1322),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1298),
.A2(n_1305),
.B(n_1306),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1353),
.A2(n_1312),
.B1(n_1407),
.B2(n_1392),
.Y(n_1456)
);

OAI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1329),
.A2(n_1363),
.B1(n_1311),
.B2(n_1284),
.C(n_1302),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1325),
.A2(n_1387),
.B(n_1407),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1344),
.B(n_1366),
.Y(n_1459)
);

BUFx4f_ASAP7_75t_L g1460 ( 
.A(n_1329),
.Y(n_1460)
);

O2A1O1Ixp5_ASAP7_75t_L g1461 ( 
.A1(n_1285),
.A2(n_1389),
.B(n_1409),
.C(n_1386),
.Y(n_1461)
);

OA21x2_ASAP7_75t_L g1462 ( 
.A1(n_1306),
.A2(n_1291),
.B(n_1288),
.Y(n_1462)
);

OA22x2_ASAP7_75t_L g1463 ( 
.A1(n_1325),
.A2(n_1312),
.B1(n_1392),
.B2(n_1372),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1317),
.B(n_1335),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1374),
.A2(n_1350),
.B1(n_1338),
.B2(n_1361),
.Y(n_1465)
);

CKINVDCx16_ASAP7_75t_R g1466 ( 
.A(n_1403),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1350),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1361),
.B(n_1330),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1319),
.A2(n_1359),
.B(n_1365),
.C(n_1381),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1319),
.B(n_1362),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1359),
.B(n_1358),
.Y(n_1471)
);

O2A1O1Ixp5_ASAP7_75t_L g1472 ( 
.A1(n_1386),
.A2(n_1398),
.B(n_1411),
.C(n_1406),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1320),
.A2(n_1343),
.B(n_1358),
.C(n_1398),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1383),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1339),
.B(n_1340),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1339),
.B(n_1393),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1294),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1374),
.Y(n_1478)
);

CKINVDCx14_ASAP7_75t_R g1479 ( 
.A(n_1338),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1294),
.B(n_1393),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1383),
.B(n_1357),
.Y(n_1481)
);

CKINVDCx12_ASAP7_75t_R g1482 ( 
.A(n_1348),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1411),
.B(n_1352),
.Y(n_1483)
);

AOI221x1_ASAP7_75t_SL g1484 ( 
.A1(n_1348),
.A2(n_1328),
.B1(n_1373),
.B2(n_1370),
.C(n_1398),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1370),
.B(n_1373),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1380),
.B(n_1385),
.Y(n_1486)
);

CKINVDCx12_ASAP7_75t_R g1487 ( 
.A(n_1405),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1377),
.B(n_1408),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1314),
.B(n_1292),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1377),
.B(n_1408),
.Y(n_1490)
);

O2A1O1Ixp5_ASAP7_75t_L g1491 ( 
.A1(n_1290),
.A2(n_1286),
.B(n_1382),
.C(n_1243),
.Y(n_1491)
);

AND2x6_ASAP7_75t_L g1492 ( 
.A(n_1325),
.B(n_1398),
.Y(n_1492)
);

NOR2xp67_ASAP7_75t_L g1493 ( 
.A(n_1315),
.B(n_1186),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1421),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1483),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1461),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1485),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1459),
.B(n_1470),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1421),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_1457),
.B(n_1433),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1462),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1455),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1422),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1437),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1426),
.B(n_1420),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_1492),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1455),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1481),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1449),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1449),
.Y(n_1510)
);

OR2x6_ASAP7_75t_L g1511 ( 
.A(n_1423),
.B(n_1416),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1441),
.Y(n_1512)
);

OAI211xp5_ASAP7_75t_L g1513 ( 
.A1(n_1429),
.A2(n_1426),
.B(n_1442),
.C(n_1431),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1472),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1468),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1474),
.B(n_1463),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1441),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1486),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1450),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1451),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1463),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1472),
.B(n_1432),
.Y(n_1522)
);

OR2x6_ASAP7_75t_L g1523 ( 
.A(n_1446),
.B(n_1473),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1469),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1432),
.A2(n_1491),
.B(n_1475),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1440),
.B(n_1418),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1487),
.Y(n_1527)
);

NOR3xp33_ASAP7_75t_L g1528 ( 
.A(n_1429),
.B(n_1491),
.C(n_1436),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1452),
.Y(n_1529)
);

AO21x2_ASAP7_75t_L g1530 ( 
.A1(n_1446),
.A2(n_1442),
.B(n_1453),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1464),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1452),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1419),
.B(n_1434),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1444),
.A2(n_1490),
.B1(n_1415),
.B2(n_1488),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1447),
.B(n_1438),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1492),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1509),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1509),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1509),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1530),
.B(n_1439),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1526),
.B(n_1534),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1531),
.B(n_1484),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1510),
.Y(n_1543)
);

INVx5_ASAP7_75t_L g1544 ( 
.A(n_1511),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1516),
.B(n_1428),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1498),
.B(n_1414),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_1504),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1531),
.B(n_1453),
.Y(n_1548)
);

AOI31xp33_ASAP7_75t_L g1549 ( 
.A1(n_1505),
.A2(n_1448),
.A3(n_1456),
.B(n_1465),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1489),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1510),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1497),
.B(n_1492),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1494),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1517),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1498),
.B(n_1445),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1499),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1498),
.B(n_1476),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1508),
.B(n_1477),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1505),
.A2(n_1513),
.B1(n_1528),
.B2(n_1511),
.C(n_1534),
.Y(n_1559)
);

AND2x4_ASAP7_75t_L g1560 ( 
.A(n_1497),
.B(n_1425),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1527),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1497),
.B(n_1480),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1503),
.Y(n_1563)
);

BUFx2_ASAP7_75t_SL g1564 ( 
.A(n_1500),
.Y(n_1564)
);

BUFx2_ASAP7_75t_SL g1565 ( 
.A(n_1500),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1518),
.B(n_1471),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1537),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1559),
.A2(n_1528),
.B1(n_1513),
.B2(n_1533),
.C(n_1529),
.Y(n_1569)
);

OAI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1559),
.A2(n_1511),
.B1(n_1533),
.B2(n_1535),
.C(n_1523),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1540),
.A2(n_1502),
.B(n_1512),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1546),
.B(n_1518),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1540),
.A2(n_1521),
.B1(n_1511),
.B2(n_1523),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1549),
.A2(n_1521),
.B1(n_1511),
.B2(n_1523),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1541),
.A2(n_1530),
.B1(n_1511),
.B2(n_1555),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1542),
.A2(n_1514),
.B(n_1496),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1542),
.A2(n_1514),
.B(n_1496),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1537),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1555),
.B(n_1525),
.C(n_1529),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1552),
.B(n_1521),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1515),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1538),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1564),
.A2(n_1511),
.B1(n_1530),
.B2(n_1532),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1561),
.Y(n_1584)
);

INVx1_ASAP7_75t_SL g1585 ( 
.A(n_1557),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1556),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1538),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1539),
.Y(n_1588)
);

INVx1_ASAP7_75t_SL g1589 ( 
.A(n_1566),
.Y(n_1589)
);

OAI321xp33_ASAP7_75t_L g1590 ( 
.A1(n_1548),
.A2(n_1523),
.A3(n_1522),
.B1(n_1532),
.B2(n_1524),
.C(n_1535),
.Y(n_1590)
);

AND2x6_ASAP7_75t_SL g1591 ( 
.A(n_1545),
.B(n_1479),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1545),
.B(n_1526),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1558),
.B(n_1563),
.Y(n_1593)
);

NOR3xp33_ASAP7_75t_L g1594 ( 
.A(n_1549),
.B(n_1561),
.C(n_1548),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1550),
.B(n_1495),
.Y(n_1595)
);

INVx4_ASAP7_75t_R g1596 ( 
.A(n_1553),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1554),
.A2(n_1507),
.B(n_1501),
.Y(n_1597)
);

OAI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1544),
.A2(n_1532),
.B(n_1443),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1518),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1564),
.A2(n_1523),
.B1(n_1535),
.B2(n_1458),
.Y(n_1600)
);

OAI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1565),
.A2(n_1523),
.B1(n_1493),
.B2(n_1526),
.C(n_1527),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1565),
.A2(n_1522),
.B1(n_1524),
.B2(n_1520),
.C(n_1519),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1543),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1552),
.B(n_1523),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1567),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1576),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1597),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1576),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1594),
.B(n_1544),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1578),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1582),
.Y(n_1611)
);

INVx4_ASAP7_75t_SL g1612 ( 
.A(n_1604),
.Y(n_1612)
);

CKINVDCx14_ASAP7_75t_R g1613 ( 
.A(n_1568),
.Y(n_1613)
);

BUFx3_ASAP7_75t_L g1614 ( 
.A(n_1577),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1587),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1571),
.A2(n_1579),
.B(n_1583),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1588),
.Y(n_1617)
);

AND2x6_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1506),
.Y(n_1618)
);

NOR2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1568),
.B(n_1424),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1577),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1596),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1584),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1604),
.B(n_1552),
.Y(n_1623)
);

INVx4_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1603),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1572),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1592),
.B(n_1551),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1563),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1530),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1572),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1604),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1628),
.B(n_1593),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1612),
.B(n_1604),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1624),
.B(n_1466),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1606),
.Y(n_1635)
);

NAND4xp25_ASAP7_75t_SL g1636 ( 
.A(n_1629),
.B(n_1569),
.C(n_1575),
.D(n_1570),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1612),
.B(n_1595),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1612),
.B(n_1595),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1605),
.B(n_1585),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1605),
.B(n_1586),
.Y(n_1640)
);

AOI211x1_ASAP7_75t_SL g1641 ( 
.A1(n_1609),
.A2(n_1574),
.B(n_1573),
.C(n_1598),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1628),
.B(n_1626),
.Y(n_1642)
);

OR2x6_ASAP7_75t_L g1643 ( 
.A(n_1624),
.B(n_1536),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1610),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1621),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1610),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1612),
.B(n_1552),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1612),
.B(n_1580),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1631),
.B(n_1580),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1611),
.B(n_1602),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1612),
.B(n_1589),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1612),
.B(n_1566),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1628),
.B(n_1626),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1631),
.B(n_1562),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1562),
.Y(n_1655)
);

NOR3xp33_ASAP7_75t_SL g1656 ( 
.A(n_1609),
.B(n_1427),
.C(n_1601),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1607),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1611),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1622),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1615),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1630),
.B(n_1581),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1606),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1623),
.B(n_1599),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1623),
.B(n_1560),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1560),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1624),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1644),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1624),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1644),
.Y(n_1670)
);

INVxp33_ASAP7_75t_L g1671 ( 
.A(n_1634),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1646),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1657),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1657),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1647),
.Y(n_1676)
);

INVxp33_ASAP7_75t_L g1677 ( 
.A(n_1656),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1646),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1660),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1657),
.Y(n_1680)
);

CKINVDCx14_ASAP7_75t_R g1681 ( 
.A(n_1643),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1641),
.B(n_1624),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1645),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1641),
.B(n_1613),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1645),
.B(n_1613),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1645),
.B(n_1622),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1648),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1633),
.B(n_1621),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1636),
.A2(n_1600),
.B1(n_1618),
.B2(n_1619),
.Y(n_1689)
);

NAND2xp33_ASAP7_75t_L g1690 ( 
.A(n_1656),
.B(n_1619),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1650),
.B(n_1660),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1666),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1662),
.B(n_1627),
.Y(n_1693)
);

INVxp33_ASAP7_75t_L g1694 ( 
.A(n_1633),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1658),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1658),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1659),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1649),
.B(n_1622),
.Y(n_1698)
);

OR2x2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.B(n_1617),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1632),
.B(n_1625),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1659),
.Y(n_1701)
);

O2A1O1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1643),
.A2(n_1608),
.B(n_1620),
.C(n_1614),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1676),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1673),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1676),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1682),
.B(n_1649),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1679),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1669),
.B(n_1649),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1669),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1670),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1672),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1671),
.B(n_1664),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1691),
.B(n_1632),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1678),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1671),
.B(n_1664),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1685),
.Y(n_1718)
);

AND3x1_ASAP7_75t_L g1719 ( 
.A(n_1684),
.B(n_1629),
.C(n_1636),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1695),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1688),
.B(n_1637),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1673),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1687),
.B(n_1647),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1690),
.A2(n_1643),
.B(n_1616),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1677),
.A2(n_1643),
.B1(n_1647),
.B2(n_1638),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1688),
.B(n_1637),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1676),
.B(n_1638),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1700),
.B(n_1642),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1719),
.A2(n_1677),
.B(n_1690),
.Y(n_1729)
);

OAI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1707),
.A2(n_1689),
.B1(n_1694),
.B2(n_1590),
.Y(n_1730)
);

AND4x1_ASAP7_75t_L g1731 ( 
.A(n_1725),
.B(n_1667),
.C(n_1702),
.D(n_1686),
.Y(n_1731)
);

AOI22x1_ASAP7_75t_L g1732 ( 
.A1(n_1724),
.A2(n_1687),
.B1(n_1683),
.B2(n_1674),
.Y(n_1732)
);

A2O1A1Ixp33_ASAP7_75t_L g1733 ( 
.A1(n_1719),
.A2(n_1694),
.B(n_1681),
.C(n_1674),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_L g1734 ( 
.A(n_1705),
.B(n_1698),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1718),
.A2(n_1681),
.B(n_1692),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1721),
.B(n_1666),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1710),
.B(n_1696),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_SL g1738 ( 
.A1(n_1706),
.A2(n_1614),
.B1(n_1616),
.B2(n_1608),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1721),
.B(n_1697),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1717),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1726),
.A2(n_1643),
.B1(n_1647),
.B2(n_1651),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1726),
.B(n_1701),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1727),
.B(n_1654),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1705),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1717),
.Y(n_1745)
);

OAI322xp33_ASAP7_75t_L g1746 ( 
.A1(n_1714),
.A2(n_1620),
.A3(n_1699),
.B1(n_1663),
.B2(n_1635),
.C1(n_1653),
.C2(n_1693),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1654),
.Y(n_1747)
);

O2A1O1Ixp5_ASAP7_75t_L g1748 ( 
.A1(n_1703),
.A2(n_1723),
.B(n_1716),
.C(n_1713),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1743),
.B(n_1727),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1744),
.B(n_1714),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1736),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1735),
.B(n_1728),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1740),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1745),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1734),
.B(n_1723),
.Y(n_1755)
);

NOR2x1_ASAP7_75t_L g1756 ( 
.A(n_1729),
.B(n_1703),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1731),
.B(n_1708),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1739),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1746),
.B(n_1728),
.Y(n_1759)
);

AOI211x1_ASAP7_75t_L g1760 ( 
.A1(n_1757),
.A2(n_1730),
.B(n_1737),
.C(n_1742),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1759),
.A2(n_1733),
.B(n_1730),
.Y(n_1761)
);

OAI211xp5_ASAP7_75t_L g1762 ( 
.A1(n_1759),
.A2(n_1732),
.B(n_1738),
.C(n_1741),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_L g1763 ( 
.A(n_1756),
.B(n_1748),
.C(n_1738),
.Y(n_1763)
);

AOI211xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1752),
.A2(n_1747),
.B(n_1708),
.C(n_1711),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1752),
.A2(n_1751),
.B1(n_1749),
.B2(n_1758),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1753),
.A2(n_1748),
.B1(n_1711),
.B2(n_1712),
.C(n_1715),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1750),
.A2(n_1715),
.B1(n_1712),
.B2(n_1720),
.C(n_1614),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1755),
.A2(n_1720),
.B(n_1723),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1751),
.Y(n_1769)
);

AOI321xp33_ASAP7_75t_L g1770 ( 
.A1(n_1761),
.A2(n_1754),
.A3(n_1723),
.B1(n_1722),
.B2(n_1704),
.C(n_1675),
.Y(n_1770)
);

OAI211xp5_ASAP7_75t_L g1771 ( 
.A1(n_1763),
.A2(n_1722),
.B(n_1704),
.C(n_1635),
.Y(n_1771)
);

OAI211xp5_ASAP7_75t_L g1772 ( 
.A1(n_1760),
.A2(n_1722),
.B(n_1704),
.C(n_1663),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1769),
.Y(n_1773)
);

XNOR2xp5_ASAP7_75t_SL g1774 ( 
.A(n_1765),
.B(n_1482),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1773),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1770),
.B(n_1454),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1772),
.B(n_1764),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1771),
.Y(n_1778)
);

INVx2_ASAP7_75t_SL g1779 ( 
.A(n_1774),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1773),
.B(n_1768),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1780),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1775),
.Y(n_1782)
);

AOI321xp33_ASAP7_75t_L g1783 ( 
.A1(n_1777),
.A2(n_1762),
.A3(n_1767),
.B1(n_1766),
.B2(n_1675),
.C(n_1680),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1776),
.A2(n_1616),
.B1(n_1651),
.B2(n_1680),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1775),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1781),
.B(n_1779),
.Y(n_1786)
);

NOR3xp33_ASAP7_75t_L g1787 ( 
.A(n_1782),
.B(n_1778),
.C(n_1776),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1785),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1788),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1787),
.B1(n_1786),
.B2(n_1784),
.Y(n_1790)
);

OR5x1_ASAP7_75t_L g1791 ( 
.A(n_1790),
.B(n_1783),
.C(n_1788),
.D(n_1614),
.E(n_1478),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1790),
.B(n_1504),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1791),
.A2(n_1661),
.B(n_1655),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1793),
.Y(n_1795)
);

NOR2x1p5_ASAP7_75t_L g1796 ( 
.A(n_1794),
.B(n_1467),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_SL g1797 ( 
.A1(n_1795),
.A2(n_1435),
.B1(n_1417),
.B2(n_1460),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1796),
.A2(n_1460),
.B1(n_1653),
.B2(n_1661),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1640),
.B(n_1639),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1797),
.B(n_1430),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1800),
.B(n_1640),
.Y(n_1801)
);

AOI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_1655),
.B1(n_1652),
.B2(n_1665),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1417),
.B(n_1639),
.C(n_1652),
.Y(n_1803)
);


endmodule