module fake_jpeg_6705_n_283 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_283);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_45;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_36),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_16),
.B1(n_15),
.B2(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_17),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_28),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_34),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_33),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_41),
.B1(n_30),
.B2(n_38),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_29),
.B1(n_21),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_56),
.B1(n_41),
.B2(n_17),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_62),
.B1(n_16),
.B2(n_15),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_21),
.B1(n_34),
.B2(n_35),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_46),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_41),
.B(n_40),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_49),
.Y(n_90)
);

NOR2x1_ASAP7_75t_R g68 ( 
.A(n_49),
.B(n_41),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_74),
.B(n_61),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_38),
.B1(n_48),
.B2(n_47),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_72),
.Y(n_95)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_78),
.B1(n_81),
.B2(n_62),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_22),
.B(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_42),
.B1(n_37),
.B2(n_47),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_27),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_27),
.Y(n_82)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_24),
.B(n_16),
.Y(n_119)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_86),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_52),
.B1(n_56),
.B2(n_51),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_92),
.B1(n_94),
.B2(n_24),
.Y(n_117)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_51),
.C(n_64),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_98),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_100),
.B1(n_80),
.B2(n_66),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_71),
.B(n_24),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_49),
.B1(n_63),
.B2(n_59),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_50),
.B1(n_57),
.B2(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_96),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_57),
.B1(n_47),
.B2(n_48),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_101),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_13),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_115),
.B1(n_122),
.B2(n_92),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_66),
.B1(n_67),
.B2(n_38),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_119),
.B(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_86),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_76),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_90),
.B(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_120),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_47),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_88),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_72),
.B1(n_71),
.B2(n_31),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_19),
.B1(n_13),
.B2(n_25),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_124),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_130),
.B1(n_117),
.B2(n_110),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_127),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_135),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_96),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_98),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_101),
.B(n_17),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_17),
.Y(n_162)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_102),
.B1(n_105),
.B2(n_106),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_139),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_114),
.B1(n_121),
.B2(n_118),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_103),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_123),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_162),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_112),
.C(n_119),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_158),
.C(n_160),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_99),
.C(n_58),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_128),
.C(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_25),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_99),
.C(n_58),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_124),
.C(n_58),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_70),
.B1(n_26),
.B2(n_25),
.Y(n_166)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_171),
.C(n_181),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_143),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_180),
.B(n_26),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_130),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_141),
.C(n_125),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_178),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_179),
.B(n_183),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_133),
.B(n_140),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_140),
.C(n_58),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_146),
.C(n_162),
.Y(n_196)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

A2O1A1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_18),
.B(n_36),
.C(n_32),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_43),
.B1(n_45),
.B2(n_36),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_188),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_26),
.B1(n_19),
.B2(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_187),
.Y(n_189)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_174),
.A2(n_152),
.A3(n_151),
.B1(n_150),
.B2(n_157),
.C1(n_146),
.C2(n_165),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_23),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_198),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_192),
.C(n_175),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_205),
.B1(n_207),
.B2(n_23),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_23),
.C(n_20),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_58),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_0),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_204),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_185),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_175),
.B(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_0),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_214),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_213),
.B(n_218),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_185),
.C(n_18),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_185),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_215),
.A2(n_225),
.B(n_194),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_198),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_208),
.B(n_199),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_200),
.C(n_201),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_195),
.B(n_0),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_219),
.A2(n_222),
.B(n_223),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_18),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_203),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_1),
.C(n_3),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_1),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_233),
.B(n_234),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_191),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_20),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_1),
.C(n_3),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_229),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_200),
.B(n_206),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_198),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_235),
.A2(n_238),
.B(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_193),
.B1(n_189),
.B2(n_207),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_221),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_189),
.B1(n_14),
.B2(n_23),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_220),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_214),
.B(n_22),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_32),
.B1(n_31),
.B2(n_20),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_210),
.A2(n_20),
.B1(n_14),
.B2(n_45),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_245),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_227),
.B(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_244),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_251),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_18),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_247),
.A2(n_248),
.B(n_22),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_18),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_250),
.C(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_45),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_239),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_228),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_255),
.B(n_259),
.Y(n_268)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_250),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_43),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_252),
.A2(n_43),
.B(n_45),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_262),
.C(n_4),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_43),
.B(n_45),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_270),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_8),
.Y(n_273)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_9),
.B(n_10),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_266),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_6),
.C(n_7),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_267),
.A2(n_269),
.B(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_6),
.C(n_7),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_7),
.B(n_8),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_271),
.Y(n_279)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_274),
.B(n_276),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_9),
.C(n_10),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_278),
.A2(n_272),
.B(n_11),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_281),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_279),
.A2(n_11),
.B(n_12),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_282),
.A2(n_277),
.B(n_11),
.Y(n_283)
);


endmodule