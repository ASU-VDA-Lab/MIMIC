module real_jpeg_5603_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_0),
.B(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_0),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_0),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_0),
.B(n_235),
.Y(n_234)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_2),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_2),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_2),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_2),
.B(n_58),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_2),
.B(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_2),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_2),
.B(n_393),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_3),
.Y(n_139)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_4),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_4),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_4),
.B(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_4),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_4),
.B(n_41),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_4),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_4),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_5),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_5),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_5),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_5),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_5),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_5),
.B(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_7),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_7),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_7),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_7),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_7),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_7),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_7),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_7),
.B(n_329),
.Y(n_328)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_8),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_8),
.Y(n_427)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_9),
.Y(n_170)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_11),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_11),
.B(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_11),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_11),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_11),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_11),
.B(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_11),
.B(n_418),
.Y(n_417)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g229 ( 
.A(n_12),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_12),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_13),
.B(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_13),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_13),
.B(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_13),
.B(n_178),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_13),
.B(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_14),
.Y(n_184)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_14),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_14),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_15),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_26),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_15),
.B(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_15),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_15),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_15),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_104),
.B(n_320),
.C(n_502),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_24),
.C(n_28),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_20),
.A2(n_28),
.B1(n_74),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_20),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_20),
.A2(n_85),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_20),
.B(n_225),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g502 ( 
.A(n_20),
.B(n_44),
.C(n_100),
.Y(n_502)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_22),
.Y(n_117)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_23),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g262 ( 
.A(n_23),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_23),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_24),
.A2(n_25),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_24),
.A2(n_25),
.B1(n_327),
.B2(n_333),
.Y(n_326)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_25),
.B(n_328),
.C(n_332),
.Y(n_483)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_27),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_28),
.A2(n_39),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_28),
.A2(n_74),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_28),
.B(n_147),
.C(n_152),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_32),
.Y(n_133)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_32),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_32),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_40),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_33),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_94),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_80),
.C(n_81),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_36),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_61),
.C(n_71),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_37),
.B(n_490),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_52),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_57),
.C(n_59),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_44),
.C(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_74),
.C(n_79),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_39),
.A2(n_75),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_39),
.B(n_115),
.C(n_119),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_39),
.A2(n_75),
.B1(n_478),
.B2(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_42),
.B(n_167),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_43),
.Y(n_370)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_43),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_44),
.A2(n_97),
.B1(n_98),
.B2(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_44),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_102),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_45),
.Y(n_175)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_47),
.A2(n_48),
.B1(n_129),
.B2(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_47),
.A2(n_48),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_48),
.B(n_126),
.C(n_129),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_48),
.B(n_191),
.C(n_320),
.Y(n_482)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_51),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_56),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_57),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_61),
.B(n_71),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_64),
.C(n_67),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_62),
.A2(n_64),
.B1(n_65),
.B2(n_473),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_62),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_64),
.A2(n_65),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_65),
.B(n_136),
.C(n_234),
.Y(n_308)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_66),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_67),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_76),
.B2(n_79),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_76),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_76),
.A2(n_79),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_79),
.B(n_191),
.C(n_287),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_80),
.B(n_81),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_86),
.B1(n_87),
.B2(n_93),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_85),
.B(n_226),
.C(n_228),
.Y(n_282)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_90),
.C(n_93),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_99),
.A2(n_100),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_99),
.A2(n_100),
.B1(n_345),
.B2(n_348),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_99),
.B(n_341),
.C(n_348),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_100),
.B(n_304),
.C(n_308),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_497),
.B(n_501),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_465),
.B(n_494),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_349),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_276),
.B(n_310),
.C(n_311),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_247),
.B(n_275),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_109),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_218),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_110),
.B(n_218),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_171),
.C(n_202),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_111),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_143),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_112),
.B(n_144),
.C(n_154),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_125),
.C(n_134),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_113),
.B(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g361 ( 
.A(n_124),
.Y(n_361)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_124),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_125),
.A2(n_134),
.B1(n_135),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_125),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_126),
.B(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_128),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_129),
.Y(n_256)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_133),
.Y(n_268)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_140),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_136),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_136),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_236),
.Y(n_269)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_139),
.Y(n_415)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_148),
.B(n_191),
.Y(n_365)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_150),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_150),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_156),
.B(n_157),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_155),
.B(n_162),
.C(n_166),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_171),
.B(n_202),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_186),
.C(n_188),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_172),
.A2(n_186),
.B1(n_187),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_172),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_177),
.C(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_174),
.B(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_174),
.B(n_430),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_180),
.B1(n_181),
.B2(n_185),
.Y(n_176)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_180),
.A2(n_181),
.B1(n_292),
.B2(n_295),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_181),
.B(n_234),
.C(n_293),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_183),
.Y(n_227)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_183),
.Y(n_364)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_184),
.Y(n_407)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_188),
.B(n_251),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.C(n_198),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_189),
.A2(n_190),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_191),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_191),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_191),
.A2(n_284),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_194),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_453)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_217),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_205),
.C(n_217),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_212),
.C(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_212),
.A2(n_328),
.B1(n_331),
.B2(n_332),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_212),
.Y(n_332)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_219),
.B(n_221),
.C(n_237),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_237),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_223),
.B(n_224),
.C(n_230),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_233),
.A2(n_234),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_233),
.A2(n_234),
.B1(n_357),
.B2(n_358),
.Y(n_394)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_234),
.B(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_238),
.B(n_240),
.C(n_241),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_243),
.B(n_245),
.C(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_273),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_248),
.B(n_273),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_253),
.C(n_270),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_249),
.A2(n_250),
.B1(n_457),
.B2(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_253),
.B(n_270),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_269),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_254),
.B(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_257),
.B(n_269),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_263),
.C(n_264),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_258),
.A2(n_259),
.B1(n_264),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_263),
.B(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_264),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_265),
.B(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_265),
.B(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_277),
.B(n_312),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_313),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_279),
.B(n_313),
.Y(n_464)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_296),
.CI(n_309),
.CON(n_279),
.SN(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_291),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_283),
.C(n_291),
.Y(n_336)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_293),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_299),
.C(n_301),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_308),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_314),
.B(n_316),
.C(n_334),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_334),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_317),
.B(n_325),
.C(n_326),
.Y(n_474)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

INVx8_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_328),
.Y(n_331)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_337),
.B2(n_338),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_335),
.B(n_339),
.C(n_340),
.Y(n_484)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

AO22x1_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_345),
.Y(n_348)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OAI31xp33_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_461),
.A3(n_462),
.B(n_464),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_455),
.B(n_460),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_442),
.B(n_454),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_395),
.B(n_441),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_381),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_354),
.B(n_381),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_366),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_355),
.B(n_367),
.C(n_378),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_362),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_356),
.B(n_363),
.C(n_365),
.Y(n_450)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_365),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_378),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.C(n_373),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_368),
.B(n_383),
.Y(n_382)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_371),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_383)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx8_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.C(n_394),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_382),
.B(n_438),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_384),
.A2(n_385),
.B1(n_394),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_391),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_386),
.A2(n_387),
.B1(n_391),
.B2(n_392),
.Y(n_408)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx5_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_394),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_435),
.B(n_440),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_420),
.B(n_434),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_409),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_409),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_408),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_406),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_406),
.C(n_408),
.Y(n_436)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx5_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_416),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_411),
.B1(n_416),
.B2(n_417),
.Y(n_432)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_428),
.B(n_433),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_429),
.B(n_432),
.Y(n_433)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_437),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_444),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_448),
.B2(n_449),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_450),
.C(n_451),
.Y(n_459)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_459),
.Y(n_460)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_491),
.Y(n_465)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_485),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_485),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_475),
.C(n_484),
.Y(n_467)
);

FAx1_ASAP7_75t_SL g493 ( 
.A(n_468),
.B(n_475),
.CI(n_484),
.CON(n_493),
.SN(n_493)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_474),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_471),
.C(n_474),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_481),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_482),
.C(n_483),
.Y(n_488)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_488),
.C(n_489),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_493),
.Y(n_495)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_493),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_500),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_500),
.Y(n_501)
);


endmodule