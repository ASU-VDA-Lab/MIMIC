module fake_netlist_1_2300_n_1489 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1489);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1489;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_1474;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g328 ( .A(n_50), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_212), .Y(n_329) );
BUFx5_ASAP7_75t_L g330 ( .A(n_270), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_258), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_11), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g333 ( .A(n_292), .B(n_163), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_221), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_5), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_57), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_184), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_190), .Y(n_338) );
CKINVDCx14_ASAP7_75t_R g339 ( .A(n_318), .Y(n_339) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_229), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_25), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_131), .Y(n_342) );
CKINVDCx5p33_ASAP7_75t_R g343 ( .A(n_60), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_322), .B(n_159), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_78), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_20), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_157), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_105), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_79), .B(n_21), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_43), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_57), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_74), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_260), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_294), .Y(n_354) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_320), .Y(n_355) );
INVx1_ASAP7_75t_SL g356 ( .A(n_312), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_96), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_205), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_75), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_3), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_68), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_11), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_150), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_13), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_324), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_154), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_145), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_123), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_172), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_280), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_0), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_87), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_199), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_166), .Y(n_374) );
CKINVDCx20_ASAP7_75t_R g375 ( .A(n_117), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_10), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_91), .Y(n_377) );
CKINVDCx16_ASAP7_75t_R g378 ( .A(n_326), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_152), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_92), .Y(n_380) );
BUFx2_ASAP7_75t_L g381 ( .A(n_251), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_6), .Y(n_382) );
BUFx3_ASAP7_75t_L g383 ( .A(n_256), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_197), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_101), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_325), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g387 ( .A(n_238), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_64), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_149), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_283), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_70), .Y(n_391) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_118), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_189), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_5), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_285), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_85), .B(n_211), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_119), .Y(n_397) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_6), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_135), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_179), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_126), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_217), .Y(n_402) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_90), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_64), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_206), .Y(n_405) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_307), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_176), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_253), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_98), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_96), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_44), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_83), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_46), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_246), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_45), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_213), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_245), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_49), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_121), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_43), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_261), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_209), .B(n_94), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_182), .Y(n_423) );
BUFx5_ASAP7_75t_L g424 ( .A(n_88), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_216), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_68), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_81), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_177), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_142), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_83), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_32), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_7), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_288), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_18), .Y(n_434) );
INVx1_ASAP7_75t_SL g435 ( .A(n_317), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_299), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_284), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_32), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_129), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_49), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_295), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_210), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_122), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_105), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_72), .Y(n_445) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_146), .Y(n_446) );
INVxp67_ASAP7_75t_L g447 ( .A(n_267), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_309), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_168), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_196), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_54), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_94), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_186), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_302), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_173), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_125), .Y(n_456) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_97), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_269), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_116), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_100), .Y(n_460) );
CKINVDCx14_ASAP7_75t_R g461 ( .A(n_114), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_55), .Y(n_462) );
CKINVDCx5p33_ASAP7_75t_R g463 ( .A(n_120), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_127), .B(n_88), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_160), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_227), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_239), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_52), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_45), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_38), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_228), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g472 ( .A(n_8), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_178), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_241), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_115), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_9), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_4), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_8), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_54), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_70), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_315), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_243), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_139), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_98), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_214), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_316), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_91), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_175), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_124), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_100), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_215), .Y(n_491) );
INVxp67_ASAP7_75t_L g492 ( .A(n_226), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_286), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_208), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_155), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_192), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_151), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_225), .Y(n_498) );
INVx3_ASAP7_75t_L g499 ( .A(n_374), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_424), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_330), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_424), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_461), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_424), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_424), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_381), .B(n_0), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_424), .Y(n_507) );
XNOR2xp5_ASAP7_75t_L g508 ( .A(n_351), .B(n_1), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_419), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_374), .B(n_1), .Y(n_510) );
CKINVDCx11_ASAP7_75t_R g511 ( .A(n_351), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_330), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_337), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_461), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_514) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_342), .Y(n_515) );
INVx4_ASAP7_75t_L g516 ( .A(n_424), .Y(n_516) );
BUFx3_ASAP7_75t_L g517 ( .A(n_337), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_330), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_330), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_424), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_380), .B(n_2), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_342), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_330), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_330), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_418), .B(n_432), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_404), .B(n_7), .Y(n_526) );
AND2x4_ASAP7_75t_L g527 ( .A(n_418), .B(n_9), .Y(n_527) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_329), .A2(n_10), .B(n_12), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_432), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_335), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_410), .B(n_12), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_445), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_342), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_342), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_335), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_411), .B(n_13), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_445), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_451), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_451), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_503), .B(n_398), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_503), .Y(n_541) );
INVx4_ASAP7_75t_L g542 ( .A(n_510), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_509), .B(n_370), .Y(n_543) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_515), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_520), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_503), .B(n_378), .Y(n_546) );
INVx2_ASAP7_75t_SL g547 ( .A(n_535), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_520), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_509), .B(n_387), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_535), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_510), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_527), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_527), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_535), .B(n_430), .Y(n_556) );
INVx3_ASAP7_75t_L g557 ( .A(n_510), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_527), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_538), .B(n_447), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_531), .A2(n_403), .B1(n_444), .B2(n_430), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_520), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_527), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_527), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_516), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_538), .B(n_466), .Y(n_565) );
BUFx10_ASAP7_75t_L g566 ( .A(n_510), .Y(n_566) );
AND2x6_ASAP7_75t_L g567 ( .A(n_510), .B(n_383), .Y(n_567) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_515), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_516), .Y(n_569) );
BUFx3_ASAP7_75t_L g570 ( .A(n_513), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_527), .A2(n_332), .B1(n_336), .B2(n_328), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_510), .B(n_358), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_538), .B(n_358), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_539), .B(n_444), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_516), .Y(n_575) );
OR2x6_ASAP7_75t_L g576 ( .A(n_514), .B(n_427), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_539), .B(n_490), .Y(n_577) );
INVx5_ASAP7_75t_L g578 ( .A(n_516), .Y(n_578) );
AND2x4_ASAP7_75t_L g579 ( .A(n_539), .B(n_470), .Y(n_579) );
AND2x6_ASAP7_75t_L g580 ( .A(n_499), .B(n_383), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_499), .B(n_491), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_525), .B(n_363), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_516), .Y(n_583) );
AND2x6_ASAP7_75t_L g584 ( .A(n_499), .B(n_498), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_499), .B(n_492), .Y(n_585) );
BUFx10_ASAP7_75t_L g586 ( .A(n_506), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_525), .B(n_363), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_499), .B(n_490), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_547), .B(n_531), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_557), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_547), .B(n_531), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_559), .B(n_521), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_551), .A2(n_549), .B1(n_541), .B2(n_543), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_551), .A2(n_536), .B1(n_506), .B2(n_526), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_553), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g596 ( .A(n_560), .B(n_530), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_557), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_542), .B(n_516), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_565), .B(n_536), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_566), .Y(n_601) );
NAND2xp33_ASAP7_75t_L g602 ( .A(n_567), .B(n_330), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_588), .B(n_536), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_556), .B(n_513), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_573), .B(n_521), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_574), .A2(n_526), .B1(n_514), .B2(n_375), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_557), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_542), .B(n_501), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_558), .A2(n_528), .B1(n_502), .B2(n_505), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_577), .B(n_513), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_572), .A2(n_507), .B(n_504), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_571), .A2(n_375), .B1(n_392), .B2(n_355), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_540), .A2(n_392), .B1(n_493), .B2(n_355), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_542), .B(n_501), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_579), .B(n_513), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_570), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_579), .B(n_517), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_562), .A2(n_537), .B(n_501), .C(n_518), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_563), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_579), .B(n_517), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_576), .A2(n_493), .B1(n_371), .B2(n_460), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_552), .Y(n_622) );
AND2x2_ASAP7_75t_SL g623 ( .A(n_552), .B(n_528), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_540), .A2(n_346), .B1(n_372), .B2(n_343), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_582), .B(n_525), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_546), .B(n_517), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_581), .B(n_517), .Y(n_627) );
OR2x2_ASAP7_75t_SL g628 ( .A(n_576), .B(n_511), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_566), .Y(n_629) );
INVx3_ASAP7_75t_L g630 ( .A(n_566), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_567), .A2(n_528), .B1(n_502), .B2(n_505), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_586), .B(n_457), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_587), .Y(n_633) );
BUFx3_ASAP7_75t_L g634 ( .A(n_570), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_585), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_576), .A2(n_385), .B1(n_413), .B2(n_376), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_576), .B(n_525), .Y(n_637) );
BUFx2_ASAP7_75t_L g638 ( .A(n_567), .Y(n_638) );
AOI22xp33_ASAP7_75t_SL g639 ( .A1(n_586), .A2(n_352), .B1(n_460), .B2(n_371), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_567), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_567), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_567), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_580), .B(n_525), .Y(n_643) );
BUFx3_ASAP7_75t_L g644 ( .A(n_580), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_545), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_545), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_554), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_580), .B(n_525), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_554), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_578), .B(n_528), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_586), .B(n_529), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_584), .A2(n_420), .B1(n_472), .B2(n_415), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_580), .B(n_530), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_580), .Y(n_654) );
BUFx3_ASAP7_75t_L g655 ( .A(n_580), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_561), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_584), .B(n_530), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_564), .B(n_529), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_564), .A2(n_504), .B(n_502), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_584), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_584), .B(n_548), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_584), .Y(n_662) );
NAND2xp33_ASAP7_75t_L g663 ( .A(n_578), .B(n_344), .Y(n_663) );
INVx5_ASAP7_75t_L g664 ( .A(n_578), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_578), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_578), .B(n_501), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_561), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_548), .B(n_368), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_550), .B(n_368), .Y(n_669) );
AND3x1_ASAP7_75t_L g670 ( .A(n_550), .B(n_508), .C(n_511), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_569), .B(n_512), .Y(n_671) );
BUFx2_ASAP7_75t_L g672 ( .A(n_575), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_575), .Y(n_673) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_569), .A2(n_352), .B1(n_470), .B2(n_345), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_583), .B(n_433), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_583), .B(n_433), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_544), .B(n_532), .Y(n_677) );
INVx3_ASAP7_75t_L g678 ( .A(n_544), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_544), .Y(n_679) );
AND2x4_ASAP7_75t_L g680 ( .A(n_544), .B(n_532), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_544), .B(n_436), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_568), .A2(n_478), .B1(n_359), .B2(n_452), .Y(n_682) );
AND2x6_ASAP7_75t_SL g683 ( .A(n_568), .B(n_508), .Y(n_683) );
NAND2x1_ASAP7_75t_L g684 ( .A(n_568), .B(n_528), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_568), .B(n_508), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_651), .B(n_388), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_637), .A2(n_339), .B1(n_422), .B2(n_436), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_637), .B(n_469), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_598), .A2(n_505), .B(n_500), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_624), .B(n_341), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_608), .A2(n_500), .B(n_512), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_589), .B(n_528), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_637), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_592), .A2(n_339), .B1(n_350), .B2(n_348), .Y(n_694) );
OAI21xp33_ASAP7_75t_SL g695 ( .A1(n_631), .A2(n_349), .B(n_537), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_685), .Y(n_696) );
O2A1O1Ixp33_ASAP7_75t_L g697 ( .A1(n_674), .A2(n_357), .B(n_361), .C(n_360), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_594), .A2(n_446), .B1(n_448), .B2(n_441), .Y(n_698) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_601), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_608), .A2(n_518), .B(n_512), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_601), .B(n_441), .Y(n_701) );
O2A1O1Ixp33_ASAP7_75t_L g702 ( .A1(n_674), .A2(n_362), .B(n_377), .C(n_364), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_591), .B(n_446), .Y(n_703) );
O2A1O1Ixp33_ASAP7_75t_L g704 ( .A1(n_599), .A2(n_382), .B(n_394), .C(n_391), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_601), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_614), .A2(n_519), .B(n_518), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_614), .A2(n_519), .B(n_518), .Y(n_707) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_644), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_622), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_612), .A2(n_489), .B1(n_412), .B2(n_426), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_632), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_613), .A2(n_489), .B1(n_434), .B2(n_438), .Y(n_712) );
AO21x1_ASAP7_75t_L g713 ( .A1(n_650), .A2(n_523), .B(n_519), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_593), .A2(n_440), .B1(n_462), .B2(n_409), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_603), .A2(n_475), .B1(n_476), .B2(n_468), .Y(n_715) );
AND2x4_ASAP7_75t_SL g716 ( .A(n_636), .B(n_477), .Y(n_716) );
NOR3xp33_ASAP7_75t_SL g717 ( .A(n_621), .B(n_605), .C(n_628), .Y(n_717) );
OR2x6_ASAP7_75t_L g718 ( .A(n_638), .B(n_479), .Y(n_718) );
BUFx2_ASAP7_75t_L g719 ( .A(n_683), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_590), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_592), .B(n_605), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g722 ( .A1(n_618), .A2(n_480), .B(n_487), .C(n_523), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_630), .B(n_373), .Y(n_723) );
NAND2xp5_ASAP7_75t_SL g724 ( .A(n_630), .B(n_393), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_671), .A2(n_524), .B(n_523), .Y(n_725) );
OAI22x1_ASAP7_75t_L g726 ( .A1(n_606), .A2(n_349), .B1(n_396), .B2(n_340), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_595), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_633), .B(n_356), .Y(n_728) );
INVx3_ASAP7_75t_L g729 ( .A(n_664), .Y(n_729) );
INVx4_ASAP7_75t_L g730 ( .A(n_664), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g731 ( .A1(n_671), .A2(n_524), .B(n_496), .Y(n_731) );
AND2x4_ASAP7_75t_L g732 ( .A(n_596), .B(n_537), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_600), .A2(n_524), .B1(n_484), .B2(n_431), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_619), .Y(n_734) );
O2A1O1Ixp5_ASAP7_75t_L g735 ( .A1(n_684), .A2(n_396), .B(n_365), .C(n_369), .Y(n_735) );
NAND2xp5_ASAP7_75t_SL g736 ( .A(n_664), .B(n_405), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_627), .A2(n_334), .B(n_331), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_604), .A2(n_610), .B(n_626), .Y(n_738) );
BUFx2_ASAP7_75t_L g739 ( .A(n_621), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_625), .B(n_668), .Y(n_740) );
OAI21xp33_ASAP7_75t_SL g741 ( .A1(n_631), .A2(n_464), .B(n_347), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_590), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_658), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_664), .B(n_414), .Y(n_744) );
OR2x6_ASAP7_75t_SL g745 ( .A(n_639), .B(n_421), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_623), .A2(n_353), .B(n_338), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_625), .B(n_463), .Y(n_747) );
AOI21x1_ASAP7_75t_L g748 ( .A1(n_653), .A2(n_333), .B(n_354), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_672), .B(n_465), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_623), .A2(n_367), .B(n_366), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_663), .A2(n_384), .B1(n_386), .B2(n_379), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_643), .A2(n_484), .B1(n_431), .B2(n_390), .Y(n_752) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_644), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_658), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_615), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_669), .B(n_435), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_597), .A2(n_484), .B1(n_431), .B2(n_395), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_652), .B(n_494), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_659), .A2(n_399), .B(n_389), .Y(n_759) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_655), .Y(n_760) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_655), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_648), .A2(n_402), .B1(n_407), .B2(n_401), .Y(n_762) );
INVx6_ASAP7_75t_L g763 ( .A(n_680), .Y(n_763) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_665), .Y(n_764) );
NOR2xp67_ASAP7_75t_L g765 ( .A(n_597), .B(n_128), .Y(n_765) );
AO21x1_ASAP7_75t_L g766 ( .A1(n_650), .A2(n_417), .B(n_416), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_L g767 ( .A1(n_618), .A2(n_428), .B(n_429), .C(n_423), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_617), .Y(n_768) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_675), .B(n_439), .C(n_437), .Y(n_769) );
NOR3xp33_ASAP7_75t_SL g770 ( .A(n_670), .B(n_443), .C(n_442), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g771 ( .A1(n_611), .A2(n_450), .B(n_453), .C(n_449), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g772 ( .A(n_629), .B(n_454), .Y(n_772) );
BUFx3_ASAP7_75t_L g773 ( .A(n_680), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g774 ( .A1(n_607), .A2(n_456), .B(n_455), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_620), .B(n_484), .Y(n_775) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_634), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_660), .B(n_458), .Y(n_777) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_640), .B(n_459), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_607), .A2(n_473), .B(n_471), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_676), .B(n_481), .Y(n_780) );
BUFx12f_ASAP7_75t_L g781 ( .A(n_634), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_682), .B(n_482), .Y(n_782) );
INVx6_ASAP7_75t_L g783 ( .A(n_677), .Y(n_783) );
OA21x2_ASAP7_75t_L g784 ( .A1(n_609), .A2(n_365), .B(n_329), .Y(n_784) );
O2A1O1Ixp5_ASAP7_75t_L g785 ( .A1(n_657), .A2(n_397), .B(n_400), .C(n_369), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g786 ( .A(n_660), .B(n_483), .Y(n_786) );
NOR2xp33_ASAP7_75t_SL g787 ( .A(n_641), .B(n_485), .Y(n_787) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_642), .Y(n_788) );
O2A1O1Ixp33_ASAP7_75t_L g789 ( .A1(n_602), .A2(n_488), .B(n_495), .C(n_486), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_649), .B(n_497), .Y(n_790) );
BUFx3_ASAP7_75t_L g791 ( .A(n_677), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_609), .A2(n_400), .B1(n_425), .B2(n_397), .Y(n_792) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_661), .A2(n_467), .B(n_425), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_654), .B(n_14), .Y(n_794) );
OR2x6_ASAP7_75t_L g795 ( .A(n_662), .B(n_467), .Y(n_795) );
NOR2x1_ASAP7_75t_L g796 ( .A(n_681), .B(n_406), .Y(n_796) );
OR2x2_ASAP7_75t_L g797 ( .A(n_649), .B(n_14), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_666), .Y(n_798) );
BUFx12f_ASAP7_75t_L g799 ( .A(n_679), .Y(n_799) );
NAND2xp5_ASAP7_75t_SL g800 ( .A(n_656), .B(n_406), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_667), .B(n_406), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_673), .A2(n_408), .B1(n_474), .B2(n_406), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_616), .B(n_15), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_667), .B(n_16), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_666), .A2(n_568), .B(n_474), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_645), .Y(n_806) );
NOR2x1_ASAP7_75t_R g807 ( .A(n_646), .B(n_408), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g808 ( .A1(n_647), .A2(n_474), .B(n_408), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_678), .A2(n_474), .B1(n_408), .B2(n_515), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_678), .A2(n_522), .B(n_515), .Y(n_810) );
OAI21x1_ASAP7_75t_L g811 ( .A1(n_684), .A2(n_132), .B(n_130), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_624), .B(n_16), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_651), .B(n_17), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_637), .A2(n_522), .B1(n_533), .B2(n_515), .Y(n_814) );
AOI21xp33_ASAP7_75t_L g815 ( .A1(n_651), .A2(n_18), .B(n_19), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_624), .B(n_19), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_622), .Y(n_817) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_637), .B(n_515), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_651), .B(n_20), .Y(n_819) );
BUFx3_ASAP7_75t_L g820 ( .A(n_665), .Y(n_820) );
AND2x2_ASAP7_75t_SL g821 ( .A(n_670), .B(n_21), .Y(n_821) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_601), .Y(n_822) );
AO32x1_ASAP7_75t_L g823 ( .A1(n_635), .A2(n_534), .A3(n_533), .B1(n_522), .B2(n_515), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_637), .B(n_22), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_L g825 ( .A1(n_674), .A2(n_24), .B(n_22), .C(n_23), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g826 ( .A1(n_637), .A2(n_533), .B1(n_522), .B2(n_534), .Y(n_826) );
OR2x6_ASAP7_75t_SL g827 ( .A(n_612), .B(n_23), .Y(n_827) );
BUFx6f_ASAP7_75t_L g828 ( .A(n_601), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_651), .B(n_24), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g830 ( .A1(n_739), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_711), .B(n_26), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_721), .A2(n_533), .B1(n_534), .B2(n_522), .Y(n_832) );
OAI21xp5_ASAP7_75t_L g833 ( .A1(n_735), .A2(n_738), .B(n_785), .Y(n_833) );
BUFx2_ASAP7_75t_L g834 ( .A(n_718), .Y(n_834) );
A2O1A1Ixp33_ASAP7_75t_L g835 ( .A1(n_740), .A2(n_534), .B(n_533), .C(n_522), .Y(n_835) );
OAI22x1_ASAP7_75t_L g836 ( .A1(n_827), .A2(n_29), .B1(n_27), .B2(n_28), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_710), .B(n_28), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_727), .Y(n_838) );
AO32x2_ASAP7_75t_L g839 ( .A1(n_792), .A2(n_534), .A3(n_533), .B1(n_522), .B2(n_33), .Y(n_839) );
OAI21xp5_ASAP7_75t_SL g840 ( .A1(n_716), .A2(n_29), .B(n_30), .Y(n_840) );
BUFx3_ASAP7_75t_L g841 ( .A(n_781), .Y(n_841) );
AND2x4_ASAP7_75t_L g842 ( .A(n_693), .B(n_30), .Y(n_842) );
BUFx3_ASAP7_75t_L g843 ( .A(n_799), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_696), .A2(n_534), .B1(n_533), .B2(n_34), .Y(n_844) );
A2O1A1Ixp33_ASAP7_75t_L g845 ( .A1(n_695), .A2(n_534), .B(n_533), .C(n_34), .Y(n_845) );
OA21x2_ASAP7_75t_L g846 ( .A1(n_811), .A2(n_534), .B(n_133), .Y(n_846) );
INVxp67_ASAP7_75t_L g847 ( .A(n_745), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_712), .A2(n_534), .B1(n_35), .B2(n_31), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_734), .Y(n_849) );
AO32x2_ASAP7_75t_L g850 ( .A1(n_752), .A2(n_31), .A3(n_33), .B1(n_35), .B2(n_36), .Y(n_850) );
AOI222xp33_ASAP7_75t_L g851 ( .A1(n_821), .A2(n_36), .B1(n_37), .B2(n_38), .C1(n_39), .C2(n_40), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_692), .A2(n_136), .B(n_134), .Y(n_852) );
O2A1O1Ixp33_ASAP7_75t_L g853 ( .A1(n_704), .A2(n_37), .B(n_39), .C(n_40), .Y(n_853) );
A2O1A1Ixp33_ASAP7_75t_L g854 ( .A1(n_722), .A2(n_41), .B(n_42), .C(n_44), .Y(n_854) );
OR2x2_ASAP7_75t_L g855 ( .A(n_698), .B(n_41), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_688), .B(n_42), .Y(n_856) );
AO31x2_ASAP7_75t_L g857 ( .A1(n_713), .A2(n_46), .A3(n_47), .B(n_48), .Y(n_857) );
OR2x2_ASAP7_75t_L g858 ( .A(n_719), .B(n_47), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_743), .B(n_48), .Y(n_859) );
INVx4_ASAP7_75t_L g860 ( .A(n_699), .Y(n_860) );
INVx2_ASAP7_75t_L g861 ( .A(n_720), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_746), .A2(n_138), .B(n_137), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_750), .A2(n_141), .B(n_140), .Y(n_863) );
AO31x2_ASAP7_75t_L g864 ( .A1(n_766), .A2(n_767), .A3(n_771), .B(n_726), .Y(n_864) );
BUFx3_ASAP7_75t_L g865 ( .A(n_820), .Y(n_865) );
OAI21xp5_ASAP7_75t_L g866 ( .A1(n_689), .A2(n_144), .B(n_143), .Y(n_866) );
A2O1A1Ixp33_ASAP7_75t_L g867 ( .A1(n_754), .A2(n_50), .B(n_51), .C(n_52), .Y(n_867) );
INVx2_ASAP7_75t_SL g868 ( .A(n_764), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_690), .B(n_51), .Y(n_869) );
O2A1O1Ixp33_ASAP7_75t_L g870 ( .A1(n_825), .A2(n_53), .B(n_55), .C(n_56), .Y(n_870) );
OAI22xp33_ASAP7_75t_L g871 ( .A1(n_718), .A2(n_53), .B1(n_56), .B2(n_58), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_717), .B(n_58), .Y(n_872) );
OAI21xp5_ASAP7_75t_L g873 ( .A1(n_691), .A2(n_148), .B(n_147), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_812), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_874) );
BUFx10_ASAP7_75t_L g875 ( .A(n_764), .Y(n_875) );
INVx3_ASAP7_75t_L g876 ( .A(n_730), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_700), .A2(n_156), .B(n_153), .Y(n_877) );
BUFx6f_ASAP7_75t_L g878 ( .A(n_699), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g879 ( .A1(n_816), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_709), .Y(n_880) );
OR2x2_ASAP7_75t_L g881 ( .A(n_686), .B(n_62), .Y(n_881) );
OAI21xp5_ASAP7_75t_L g882 ( .A1(n_706), .A2(n_161), .B(n_158), .Y(n_882) );
INVx5_ASAP7_75t_L g883 ( .A(n_699), .Y(n_883) );
AO32x2_ASAP7_75t_L g884 ( .A1(n_714), .A2(n_65), .A3(n_66), .B1(n_67), .B2(n_69), .Y(n_884) );
AO31x2_ASAP7_75t_L g885 ( .A1(n_778), .A2(n_65), .A3(n_66), .B(n_67), .Y(n_885) );
AO31x2_ASAP7_75t_L g886 ( .A1(n_826), .A2(n_69), .A3(n_71), .B(n_72), .Y(n_886) );
OAI21xp33_ASAP7_75t_L g887 ( .A1(n_694), .A2(n_71), .B(n_73), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_817), .Y(n_888) );
AO221x1_ASAP7_75t_L g889 ( .A1(n_687), .A2(n_73), .B1(n_74), .B2(n_75), .C(n_76), .Y(n_889) );
OAI21x1_ASAP7_75t_L g890 ( .A1(n_796), .A2(n_164), .B(n_162), .Y(n_890) );
AO32x2_ASAP7_75t_L g891 ( .A1(n_741), .A2(n_76), .A3(n_77), .B1(n_78), .B2(n_79), .Y(n_891) );
O2A1O1Ixp5_ASAP7_75t_L g892 ( .A1(n_748), .A2(n_829), .B(n_819), .C(n_813), .Y(n_892) );
NAND2x1p5_ASAP7_75t_L g893 ( .A(n_822), .B(n_77), .Y(n_893) );
AO31x2_ASAP7_75t_L g894 ( .A1(n_794), .A2(n_80), .A3(n_81), .B(n_82), .Y(n_894) );
INVx5_ASAP7_75t_L g895 ( .A(n_822), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_755), .B(n_80), .Y(n_896) );
OR2x2_ASAP7_75t_L g897 ( .A(n_715), .B(n_82), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_768), .B(n_84), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_764), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_707), .A2(n_236), .B(n_323), .Y(n_900) );
O2A1O1Ixp33_ASAP7_75t_L g901 ( .A1(n_697), .A2(n_84), .B(n_85), .C(n_86), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_824), .A2(n_87), .B1(n_89), .B2(n_90), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_769), .B(n_89), .Y(n_903) );
A2O1A1Ixp33_ASAP7_75t_L g904 ( .A1(n_737), .A2(n_92), .B(n_93), .C(n_95), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_797), .Y(n_905) );
HB1xp67_ASAP7_75t_L g906 ( .A(n_718), .Y(n_906) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_756), .B(n_93), .C(n_95), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_790), .Y(n_908) );
INVx2_ASAP7_75t_SL g909 ( .A(n_732), .Y(n_909) );
BUFx6f_ASAP7_75t_L g910 ( .A(n_822), .Y(n_910) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_773), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_725), .A2(n_242), .B(n_321), .Y(n_912) );
OAI21xp5_ASAP7_75t_L g913 ( .A1(n_731), .A2(n_240), .B(n_319), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_732), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_742), .Y(n_915) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_751), .B(n_97), .C(n_99), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_770), .B(n_99), .Y(n_917) );
OAI21x1_ASAP7_75t_L g918 ( .A1(n_805), .A2(n_237), .B(n_314), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_758), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g920 ( .A1(n_783), .A2(n_103), .B1(n_104), .B2(n_106), .Y(n_920) );
BUFx8_ASAP7_75t_SL g921 ( .A(n_798), .Y(n_921) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_703), .B(n_104), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_789), .A2(n_106), .B(n_107), .C(n_108), .Y(n_923) );
AO31x2_ASAP7_75t_L g924 ( .A1(n_793), .A2(n_107), .A3(n_108), .B(n_109), .Y(n_924) );
INVx2_ASAP7_75t_SL g925 ( .A(n_730), .Y(n_925) );
AND2x4_ASAP7_75t_L g926 ( .A(n_729), .B(n_109), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_806), .Y(n_927) );
INVx3_ASAP7_75t_L g928 ( .A(n_828), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_702), .B(n_110), .Y(n_929) );
AO31x2_ASAP7_75t_L g930 ( .A1(n_803), .A2(n_110), .A3(n_111), .B(n_112), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_804), .Y(n_931) );
OAI21x1_ASAP7_75t_L g932 ( .A1(n_818), .A2(n_247), .B(n_313), .Y(n_932) );
NOR2xp67_ASAP7_75t_L g933 ( .A(n_729), .B(n_111), .Y(n_933) );
NAND2x1_ASAP7_75t_L g934 ( .A(n_828), .B(n_165), .Y(n_934) );
O2A1O1Ixp33_ASAP7_75t_L g935 ( .A1(n_815), .A2(n_112), .B(n_113), .C(n_114), .Y(n_935) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_728), .B(n_113), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_780), .Y(n_937) );
INVx3_ASAP7_75t_L g938 ( .A(n_776), .Y(n_938) );
O2A1O1Ixp33_ASAP7_75t_L g939 ( .A1(n_782), .A2(n_115), .B(n_167), .C(n_169), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_772), .A2(n_170), .B(n_171), .Y(n_940) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_762), .A2(n_174), .B1(n_180), .B2(n_181), .C(n_183), .Y(n_941) );
HB1xp67_ASAP7_75t_L g942 ( .A(n_791), .Y(n_942) );
BUFx2_ASAP7_75t_L g943 ( .A(n_807), .Y(n_943) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_783), .A2(n_185), .B1(n_187), .B2(n_188), .Y(n_944) );
OAI21x1_ASAP7_75t_L g945 ( .A1(n_784), .A2(n_191), .B(n_193), .Y(n_945) );
AOI22xp5_ASAP7_75t_L g946 ( .A1(n_747), .A2(n_194), .B1(n_195), .B2(n_198), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_776), .Y(n_947) );
BUFx3_ASAP7_75t_L g948 ( .A(n_763), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_775), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_763), .A2(n_200), .B1(n_201), .B2(n_202), .Y(n_950) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_776), .Y(n_951) );
OAI22x1_ASAP7_75t_L g952 ( .A1(n_807), .A2(n_203), .B1(n_204), .B2(n_207), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_749), .A2(n_218), .B1(n_219), .B2(n_220), .Y(n_953) );
OAI21x1_ASAP7_75t_L g954 ( .A1(n_784), .A2(n_222), .B(n_223), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g955 ( .A1(n_795), .A2(n_224), .B1(n_230), .B2(n_231), .Y(n_955) );
INVx4_ASAP7_75t_L g956 ( .A(n_705), .Y(n_956) );
AOI221x1_ASAP7_75t_L g957 ( .A1(n_802), .A2(n_232), .B1(n_233), .B2(n_234), .C(n_235), .Y(n_957) );
AOI21xp33_ASAP7_75t_L g958 ( .A1(n_788), .A2(n_244), .B(n_248), .Y(n_958) );
AO31x2_ASAP7_75t_L g959 ( .A1(n_733), .A2(n_249), .A3(n_250), .B(n_252), .Y(n_959) );
AND2x2_ASAP7_75t_L g960 ( .A(n_701), .B(n_254), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_705), .Y(n_961) );
INVx5_ASAP7_75t_L g962 ( .A(n_708), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g963 ( .A1(n_787), .A2(n_255), .B1(n_257), .B2(n_259), .Y(n_963) );
AOI21xp5_ASAP7_75t_L g964 ( .A1(n_777), .A2(n_262), .B(n_263), .Y(n_964) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_795), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_795), .A2(n_264), .B1(n_265), .B2(n_266), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g967 ( .A1(n_786), .A2(n_268), .B(n_271), .Y(n_967) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_708), .Y(n_968) );
O2A1O1Ixp33_ASAP7_75t_SL g969 ( .A1(n_800), .A2(n_272), .B(n_273), .C(n_274), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_759), .Y(n_970) );
O2A1O1Ixp33_ASAP7_75t_SL g971 ( .A1(n_801), .A2(n_275), .B(n_276), .C(n_277), .Y(n_971) );
AO32x2_ASAP7_75t_L g972 ( .A1(n_823), .A2(n_278), .A3(n_279), .B1(n_281), .B2(n_282), .Y(n_972) );
AOI21xp5_ASAP7_75t_L g973 ( .A1(n_823), .A2(n_287), .B(n_289), .Y(n_973) );
A2O1A1Ixp33_ASAP7_75t_L g974 ( .A1(n_774), .A2(n_290), .B(n_291), .C(n_293), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_779), .Y(n_975) );
CKINVDCx5p33_ASAP7_75t_R g976 ( .A(n_736), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_723), .B(n_296), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_724), .B(n_297), .Y(n_978) );
AOI221x1_ASAP7_75t_L g979 ( .A1(n_808), .A2(n_298), .B1(n_300), .B2(n_301), .C(n_303), .Y(n_979) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_823), .A2(n_810), .B(n_744), .Y(n_980) );
AND2x4_ASAP7_75t_L g981 ( .A(n_708), .B(n_327), .Y(n_981) );
OA21x2_ASAP7_75t_L g982 ( .A1(n_765), .A2(n_304), .B(n_305), .Y(n_982) );
A2O1A1Ixp33_ASAP7_75t_L g983 ( .A1(n_757), .A2(n_306), .B(n_308), .C(n_310), .Y(n_983) );
A2O1A1Ixp33_ASAP7_75t_L g984 ( .A1(n_814), .A2(n_311), .B(n_753), .C(n_760), .Y(n_984) );
NAND3xp33_ASAP7_75t_SL g985 ( .A(n_809), .B(n_753), .C(n_760), .Y(n_985) );
BUFx6f_ASAP7_75t_L g986 ( .A(n_761), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_761), .B(n_739), .Y(n_987) );
OAI21x1_ASAP7_75t_L g988 ( .A1(n_761), .A2(n_811), .B(n_684), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_727), .Y(n_989) );
NAND3xp33_ASAP7_75t_L g990 ( .A(n_741), .B(n_717), .C(n_769), .Y(n_990) );
O2A1O1Ixp33_ASAP7_75t_L g991 ( .A1(n_721), .A2(n_704), .B(n_825), .C(n_771), .Y(n_991) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_711), .B(n_613), .Y(n_992) );
BUFx8_ASAP7_75t_L g993 ( .A(n_719), .Y(n_993) );
AO31x2_ASAP7_75t_L g994 ( .A1(n_845), .A2(n_835), .A3(n_980), .B(n_979), .Y(n_994) );
AO31x2_ASAP7_75t_L g995 ( .A1(n_973), .A2(n_957), .A3(n_970), .B(n_975), .Y(n_995) );
OAI21x1_ASAP7_75t_L g996 ( .A1(n_988), .A2(n_954), .B(n_945), .Y(n_996) );
AO21x2_ASAP7_75t_L g997 ( .A1(n_833), .A2(n_985), .B(n_862), .Y(n_997) );
BUFx3_ASAP7_75t_L g998 ( .A(n_843), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_937), .B(n_908), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_942), .B(n_834), .Y(n_1000) );
AND2x2_ASAP7_75t_SL g1001 ( .A(n_943), .B(n_842), .Y(n_1001) );
OA21x2_ASAP7_75t_L g1002 ( .A1(n_892), .A2(n_882), .B(n_873), .Y(n_1002) );
INVx4_ASAP7_75t_SL g1003 ( .A(n_878), .Y(n_1003) );
INVx8_ASAP7_75t_L g1004 ( .A(n_883), .Y(n_1004) );
OAI22xp33_ASAP7_75t_L g1005 ( .A1(n_855), .A2(n_897), .B1(n_840), .B2(n_837), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_906), .B(n_929), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_869), .A2(n_990), .B1(n_992), .B2(n_856), .Y(n_1007) );
AOI21xp5_ASAP7_75t_L g1008 ( .A1(n_991), .A2(n_931), .B(n_949), .Y(n_1008) );
AO21x2_ASAP7_75t_L g1009 ( .A1(n_832), .A2(n_913), .B(n_866), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_838), .B(n_849), .Y(n_1010) );
A2O1A1Ixp33_ASAP7_75t_L g1011 ( .A1(n_922), .A2(n_936), .B(n_870), .C(n_887), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_872), .A2(n_889), .B1(n_847), .B2(n_987), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_876), .B(n_989), .Y(n_1013) );
A2O1A1Ixp33_ASAP7_75t_L g1014 ( .A1(n_853), .A2(n_901), .B(n_935), .C(n_907), .Y(n_1014) );
INVx1_ASAP7_75t_SL g1015 ( .A(n_875), .Y(n_1015) );
OA21x2_ASAP7_75t_L g1016 ( .A1(n_932), .A2(n_890), .B(n_852), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_880), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_859), .A2(n_863), .B(n_898), .Y(n_1018) );
INVx2_ASAP7_75t_L g1019 ( .A(n_888), .Y(n_1019) );
INVx1_ASAP7_75t_L g1020 ( .A(n_842), .Y(n_1020) );
OA21x2_ASAP7_75t_L g1021 ( .A1(n_918), .A2(n_984), .B(n_974), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_905), .B(n_927), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g1023 ( .A(n_993), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_861), .B(n_915), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_896), .B(n_881), .Y(n_1025) );
INVx1_ASAP7_75t_L g1026 ( .A(n_926), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1027 ( .A(n_865), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_926), .A2(n_893), .B1(n_965), .B2(n_902), .Y(n_1028) );
OA21x2_ASAP7_75t_L g1029 ( .A1(n_877), .A2(n_900), .B(n_912), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1030 ( .A(n_841), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_917), .B(n_851), .Y(n_1031) );
OAI21x1_ASAP7_75t_L g1032 ( .A1(n_934), .A2(n_928), .B(n_982), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g1033 ( .A(n_911), .Y(n_1033) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_836), .A2(n_871), .B1(n_831), .B2(n_874), .C(n_903), .Y(n_1034) );
AO31x2_ASAP7_75t_L g1035 ( .A1(n_854), .A2(n_923), .A3(n_952), .B(n_867), .Y(n_1035) );
INVx4_ASAP7_75t_L g1036 ( .A(n_883), .Y(n_1036) );
NOR2xp33_ASAP7_75t_L g1037 ( .A(n_909), .B(n_914), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_948), .B(n_875), .Y(n_1038) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_921), .Y(n_1039) );
OR2x6_ASAP7_75t_L g1040 ( .A(n_925), .B(n_868), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1041 ( .A(n_864), .B(n_876), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_930), .Y(n_1042) );
AND2x4_ASAP7_75t_L g1043 ( .A(n_883), .B(n_895), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_895), .B(n_962), .Y(n_1044) );
OAI221xp5_ASAP7_75t_L g1045 ( .A1(n_879), .A2(n_919), .B1(n_848), .B2(n_830), .C(n_904), .Y(n_1045) );
BUFx12f_ASAP7_75t_L g1046 ( .A(n_993), .Y(n_1046) );
NAND2xp5_ASAP7_75t_SL g1047 ( .A(n_895), .B(n_962), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_864), .B(n_899), .Y(n_1048) );
BUFx3_ASAP7_75t_L g1049 ( .A(n_962), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_977), .B(n_978), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_947), .B(n_961), .Y(n_1051) );
AOI21xp5_ASAP7_75t_L g1052 ( .A1(n_969), .A2(n_971), .B(n_941), .Y(n_1052) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_968), .B(n_951), .Y(n_1053) );
AOI22xp33_ASAP7_75t_SL g1054 ( .A1(n_920), .A2(n_916), .B1(n_858), .B2(n_966), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g1055 ( .A(n_976), .Y(n_1055) );
OR2x2_ASAP7_75t_L g1056 ( .A(n_894), .B(n_938), .Y(n_1056) );
AOI222xp33_ASAP7_75t_L g1057 ( .A1(n_933), .A2(n_955), .B1(n_844), .B2(n_960), .C1(n_944), .C2(n_981), .Y(n_1057) );
OAI21xp5_ASAP7_75t_L g1058 ( .A1(n_964), .A2(n_967), .B(n_946), .Y(n_1058) );
OAI21x1_ASAP7_75t_L g1059 ( .A1(n_940), .A2(n_953), .B(n_950), .Y(n_1059) );
AO31x2_ASAP7_75t_L g1060 ( .A1(n_983), .A2(n_860), .A3(n_839), .B(n_956), .Y(n_1060) );
AO31x2_ASAP7_75t_L g1061 ( .A1(n_860), .A2(n_956), .A3(n_972), .B(n_857), .Y(n_1061) );
AO21x2_ASAP7_75t_L g1062 ( .A1(n_958), .A2(n_981), .B(n_972), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1063 ( .A1(n_963), .A2(n_986), .B1(n_910), .B2(n_878), .C(n_884), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_884), .Y(n_1064) );
INVx2_ASAP7_75t_L g1065 ( .A(n_857), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g1066 ( .A(n_878), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_924), .Y(n_1067) );
OR2x6_ASAP7_75t_L g1068 ( .A(n_910), .B(n_986), .Y(n_1068) );
OA21x2_ASAP7_75t_L g1069 ( .A1(n_972), .A2(n_857), .B(n_891), .Y(n_1069) );
NOR3xp33_ASAP7_75t_L g1070 ( .A(n_891), .B(n_850), .C(n_885), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_986), .B(n_910), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_894), .B(n_924), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_894), .B(n_885), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_850), .A2(n_886), .B1(n_885), .B2(n_959), .Y(n_1074) );
OA21x2_ASAP7_75t_L g1075 ( .A1(n_959), .A2(n_886), .B(n_850), .Y(n_1075) );
AO21x1_ASAP7_75t_L g1076 ( .A1(n_886), .A2(n_939), .B(n_935), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g1077 ( .A(n_921), .Y(n_1077) );
BUFx3_ASAP7_75t_L g1078 ( .A(n_843), .Y(n_1078) );
CKINVDCx6p67_ASAP7_75t_R g1079 ( .A(n_841), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_942), .Y(n_1080) );
OAI22xp33_ASAP7_75t_L g1081 ( .A1(n_855), .A2(n_739), .B1(n_612), .B2(n_621), .Y(n_1081) );
BUFx3_ASAP7_75t_L g1082 ( .A(n_843), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_838), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_942), .B(n_612), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_937), .B(n_721), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_833), .A2(n_663), .B(n_980), .Y(n_1086) );
AND2x2_ASAP7_75t_SL g1087 ( .A(n_834), .B(n_943), .Y(n_1087) );
A2O1A1Ixp33_ASAP7_75t_L g1088 ( .A1(n_991), .A2(n_990), .B(n_740), .C(n_922), .Y(n_1088) );
AOI22xp33_ASAP7_75t_SL g1089 ( .A1(n_834), .A2(n_739), .B1(n_612), .B2(n_842), .Y(n_1089) );
NAND3xp33_ASAP7_75t_L g1090 ( .A(n_990), .B(n_845), .C(n_741), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_834), .B(n_637), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_834), .B(n_637), .Y(n_1092) );
OA21x2_ASAP7_75t_L g1093 ( .A1(n_945), .A2(n_954), .B(n_980), .Y(n_1093) );
AOI21x1_ASAP7_75t_L g1094 ( .A1(n_980), .A2(n_973), .B(n_846), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_937), .B(n_721), .Y(n_1095) );
INVx3_ASAP7_75t_L g1096 ( .A(n_875), .Y(n_1096) );
OAI21xp5_ASAP7_75t_L g1097 ( .A1(n_845), .A2(n_695), .B(n_738), .Y(n_1097) );
INVx2_ASAP7_75t_L g1098 ( .A(n_838), .Y(n_1098) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_942), .B(n_612), .Y(n_1099) );
INVx1_ASAP7_75t_L g1100 ( .A(n_838), .Y(n_1100) );
AOI21xp5_ASAP7_75t_L g1101 ( .A1(n_833), .A2(n_663), .B(n_980), .Y(n_1101) );
AOI21xp5_ASAP7_75t_L g1102 ( .A1(n_833), .A2(n_663), .B(n_980), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g1103 ( .A(n_992), .B(n_739), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_937), .B(n_721), .Y(n_1104) );
INVx2_ASAP7_75t_L g1105 ( .A(n_838), .Y(n_1105) );
NOR2xp33_ASAP7_75t_L g1106 ( .A(n_992), .B(n_739), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_838), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_834), .B(n_637), .Y(n_1108) );
INVxp67_ASAP7_75t_L g1109 ( .A(n_842), .Y(n_1109) );
A2O1A1Ixp33_ASAP7_75t_L g1110 ( .A1(n_991), .A2(n_990), .B(n_740), .C(n_922), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_937), .B(n_721), .Y(n_1111) );
INVx4_ASAP7_75t_L g1112 ( .A(n_883), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_937), .B(n_721), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_838), .Y(n_1114) );
INVx4_ASAP7_75t_L g1115 ( .A(n_883), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_838), .Y(n_1116) );
A2O1A1Ixp33_ASAP7_75t_L g1117 ( .A1(n_991), .A2(n_990), .B(n_740), .C(n_922), .Y(n_1117) );
CKINVDCx11_ASAP7_75t_R g1118 ( .A(n_841), .Y(n_1118) );
INVx1_ASAP7_75t_SL g1119 ( .A(n_834), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_937), .B(n_721), .Y(n_1120) );
BUFx8_ASAP7_75t_L g1121 ( .A(n_841), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g1122 ( .A(n_942), .Y(n_1122) );
BUFx6f_ASAP7_75t_L g1123 ( .A(n_878), .Y(n_1123) );
NAND2xp5_ASAP7_75t_SL g1124 ( .A(n_834), .B(n_943), .Y(n_1124) );
BUFx4f_ASAP7_75t_SL g1125 ( .A(n_841), .Y(n_1125) );
OAI21x1_ASAP7_75t_L g1126 ( .A1(n_988), .A2(n_980), .B(n_954), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_838), .Y(n_1127) );
INVx2_ASAP7_75t_SL g1128 ( .A(n_875), .Y(n_1128) );
INVx2_ASAP7_75t_L g1129 ( .A(n_838), .Y(n_1129) );
OAI21xp33_ASAP7_75t_L g1130 ( .A1(n_869), .A2(n_639), .B(n_717), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_838), .Y(n_1131) );
HB1xp67_ASAP7_75t_L g1132 ( .A(n_942), .Y(n_1132) );
OA21x2_ASAP7_75t_L g1133 ( .A1(n_945), .A2(n_954), .B(n_980), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_937), .B(n_721), .Y(n_1134) );
INVx2_ASAP7_75t_L g1135 ( .A(n_838), .Y(n_1135) );
INVx2_ASAP7_75t_L g1136 ( .A(n_838), .Y(n_1136) );
OA21x2_ASAP7_75t_L g1137 ( .A1(n_945), .A2(n_954), .B(n_980), .Y(n_1137) );
NAND2xp5_ASAP7_75t_SL g1138 ( .A(n_1005), .B(n_1001), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1041), .Y(n_1139) );
OAI21xp5_ASAP7_75t_L g1140 ( .A1(n_1088), .A2(n_1117), .B(n_1110), .Y(n_1140) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1041), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_999), .B(n_1024), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_999), .B(n_1024), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1006), .B(n_1019), .Y(n_1144) );
AO21x2_ASAP7_75t_L g1145 ( .A1(n_1086), .A2(n_1102), .B(n_1101), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1146 ( .A(n_1004), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1098), .B(n_1105), .Y(n_1147) );
INVx2_ASAP7_75t_L g1148 ( .A(n_1065), .Y(n_1148) );
INVx3_ASAP7_75t_L g1149 ( .A(n_1004), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1067), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1151 ( .A1(n_1007), .A2(n_1130), .B1(n_1034), .B2(n_1089), .C(n_1103), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_1080), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_1031), .A2(n_1106), .B1(n_1034), .B2(n_1081), .Y(n_1153) );
NAND2xp5_ASAP7_75t_SL g1154 ( .A(n_1028), .B(n_1087), .Y(n_1154) );
INVx2_ASAP7_75t_SL g1155 ( .A(n_1004), .Y(n_1155) );
AND2x4_ASAP7_75t_SL g1156 ( .A(n_1079), .B(n_1044), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1085), .B(n_1095), .Y(n_1157) );
AO21x2_ASAP7_75t_L g1158 ( .A1(n_1072), .A2(n_1073), .B(n_1070), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1042), .Y(n_1159) );
AO21x2_ASAP7_75t_L g1160 ( .A1(n_1072), .A2(n_1073), .B(n_1094), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1048), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1048), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1163 ( .A(n_1109), .B(n_1084), .Y(n_1163) );
INVx2_ASAP7_75t_SL g1164 ( .A(n_1044), .Y(n_1164) );
INVx3_ASAP7_75t_L g1165 ( .A(n_1043), .Y(n_1165) );
OA21x2_ASAP7_75t_L g1166 ( .A1(n_1126), .A2(n_1074), .B(n_996), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1129), .B(n_1135), .Y(n_1167) );
AOI21xp5_ASAP7_75t_SL g1168 ( .A1(n_1028), .A2(n_1063), .B(n_1062), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1136), .B(n_1017), .Y(n_1169) );
INVx3_ASAP7_75t_L g1170 ( .A(n_1043), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1064), .Y(n_1171) );
OR2x6_ASAP7_75t_L g1172 ( .A(n_1036), .B(n_1112), .Y(n_1172) );
OA21x2_ASAP7_75t_L g1173 ( .A1(n_1076), .A2(n_1097), .B(n_1032), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1085), .B(n_1095), .Y(n_1174) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_1045), .A2(n_1012), .B1(n_1054), .B2(n_1099), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1056), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1083), .B(n_1100), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1178 ( .A1(n_1104), .A2(n_1134), .B1(n_1113), .B2(n_1111), .C(n_1120), .Y(n_1178) );
AO21x2_ASAP7_75t_L g1179 ( .A1(n_1097), .A2(n_1090), .B(n_997), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1010), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1107), .B(n_1114), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1182 ( .A(n_1010), .B(n_1104), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1116), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1111), .B(n_1113), .Y(n_1184) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1127), .Y(n_1185) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1068), .Y(n_1186) );
BUFx3_ASAP7_75t_L g1187 ( .A(n_1125), .Y(n_1187) );
HB1xp67_ASAP7_75t_L g1188 ( .A(n_1122), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1003), .B(n_1071), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1131), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1075), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1120), .B(n_1134), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g1193 ( .A1(n_1050), .A2(n_1020), .B1(n_1045), .B2(n_1026), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_1011), .A2(n_1014), .B1(n_1025), .B2(n_1050), .C(n_1119), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1195 ( .A(n_1068), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1053), .B(n_1022), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1008), .B(n_1013), .Y(n_1197) );
BUFx3_ASAP7_75t_L g1198 ( .A(n_1030), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1069), .Y(n_1199) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1123), .Y(n_1200) );
INVx2_ASAP7_75t_L g1201 ( .A(n_1069), .Y(n_1201) );
OA21x2_ASAP7_75t_L g1202 ( .A1(n_1090), .A2(n_1018), .B(n_1052), .Y(n_1202) );
INVx2_ASAP7_75t_SL g1203 ( .A(n_1049), .Y(n_1203) );
AO21x2_ASAP7_75t_L g1204 ( .A1(n_997), .A2(n_1062), .B(n_1009), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1205 ( .A1(n_1025), .A2(n_1037), .B1(n_1132), .B2(n_1022), .C(n_1119), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1013), .B(n_1091), .Y(n_1206) );
AOI222xp33_ASAP7_75t_L g1207 ( .A1(n_1046), .A2(n_1039), .B1(n_1121), .B2(n_1124), .C1(n_1092), .C2(n_1108), .Y(n_1207) );
AOI22xp33_ASAP7_75t_L g1208 ( .A1(n_1057), .A2(n_1033), .B1(n_1000), .B2(n_1027), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1061), .Y(n_1209) );
INVx4_ASAP7_75t_L g1210 ( .A(n_1036), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_995), .Y(n_1211) );
INVx2_ASAP7_75t_L g1212 ( .A(n_995), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1040), .B(n_1053), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1040), .B(n_1051), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1040), .B(n_1051), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1035), .B(n_1015), .Y(n_1216) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1061), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1061), .Y(n_1218) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1071), .Y(n_1219) );
OR2x6_ASAP7_75t_L g1220 ( .A(n_1112), .B(n_1115), .Y(n_1220) );
INVx3_ASAP7_75t_SL g1221 ( .A(n_1023), .Y(n_1221) );
BUFx2_ASAP7_75t_L g1222 ( .A(n_1068), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g1223 ( .A1(n_1057), .A2(n_1058), .B1(n_1082), .B2(n_998), .C(n_1078), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_995), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1035), .B(n_1015), .Y(n_1225) );
AO21x2_ASAP7_75t_L g1226 ( .A1(n_1059), .A2(n_994), .B(n_1060), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1038), .B(n_1128), .Y(n_1227) );
AO21x2_ASAP7_75t_L g1228 ( .A1(n_994), .A2(n_1060), .B(n_1066), .Y(n_1228) );
AO21x2_ASAP7_75t_L g1229 ( .A1(n_994), .A2(n_1060), .B(n_1133), .Y(n_1229) );
OR2x2_ASAP7_75t_L g1230 ( .A(n_1096), .B(n_1115), .Y(n_1230) );
INVxp33_ASAP7_75t_L g1231 ( .A(n_1118), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1035), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1003), .B(n_1047), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1234 ( .A(n_1002), .B(n_1137), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1093), .Y(n_1235) );
AOI21xp5_ASAP7_75t_SL g1236 ( .A1(n_1021), .A2(n_1016), .B(n_1029), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1055), .B(n_1121), .Y(n_1237) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1003), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1016), .Y(n_1239) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1152), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1150), .Y(n_1241) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1201), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1142), .B(n_1077), .Y(n_1243) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1150), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1143), .B(n_1176), .Y(n_1245) );
AOI22xp33_ASAP7_75t_SL g1246 ( .A1(n_1175), .A2(n_1151), .B1(n_1223), .B2(n_1188), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1143), .B(n_1176), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1216), .B(n_1225), .Y(n_1248) );
BUFx2_ASAP7_75t_L g1249 ( .A(n_1195), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1180), .B(n_1178), .Y(n_1250) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1196), .B(n_1182), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1216), .B(n_1225), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1144), .B(n_1232), .Y(n_1253) );
OR2x6_ASAP7_75t_L g1254 ( .A(n_1168), .B(n_1154), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1144), .B(n_1232), .Y(n_1255) );
AO21x2_ASAP7_75t_L g1256 ( .A1(n_1236), .A2(n_1239), .B(n_1224), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1219), .B(n_1139), .Y(n_1257) );
INVxp67_ASAP7_75t_L g1258 ( .A(n_1214), .Y(n_1258) );
OAI22xp5_ASAP7_75t_L g1259 ( .A1(n_1153), .A2(n_1138), .B1(n_1182), .B2(n_1192), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1196), .B(n_1141), .Y(n_1260) );
BUFx2_ASAP7_75t_L g1261 ( .A(n_1195), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1141), .B(n_1161), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_1194), .A2(n_1208), .B1(n_1197), .B2(n_1140), .Y(n_1263) );
BUFx2_ASAP7_75t_L g1264 ( .A(n_1222), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1183), .B(n_1185), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1161), .B(n_1162), .Y(n_1266) );
INVxp67_ASAP7_75t_SL g1267 ( .A(n_1148), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1183), .B(n_1185), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1162), .B(n_1147), .Y(n_1269) );
INVx4_ASAP7_75t_L g1270 ( .A(n_1210), .Y(n_1270) );
BUFx2_ASAP7_75t_L g1271 ( .A(n_1222), .Y(n_1271) );
AND2x4_ASAP7_75t_L g1272 ( .A(n_1159), .B(n_1197), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1147), .B(n_1167), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1167), .B(n_1177), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1177), .B(n_1181), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1190), .B(n_1157), .Y(n_1276) );
OAI33xp33_ASAP7_75t_L g1277 ( .A1(n_1190), .A2(n_1184), .A3(n_1174), .B1(n_1227), .B2(n_1230), .B3(n_1199), .Y(n_1277) );
HB1xp67_ASAP7_75t_L g1278 ( .A(n_1213), .Y(n_1278) );
AND2x4_ASAP7_75t_L g1279 ( .A(n_1199), .B(n_1191), .Y(n_1279) );
BUFx3_ASAP7_75t_L g1280 ( .A(n_1172), .Y(n_1280) );
NOR2xp33_ASAP7_75t_L g1281 ( .A(n_1198), .B(n_1221), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1282 ( .A(n_1213), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1181), .B(n_1171), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_1214), .Y(n_1284) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_1156), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1171), .B(n_1169), .Y(n_1286) );
INVxp67_ASAP7_75t_L g1287 ( .A(n_1215), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1193), .B(n_1169), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1215), .B(n_1158), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1290 ( .A(n_1189), .Y(n_1290) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1209), .Y(n_1291) );
BUFx3_ASAP7_75t_L g1292 ( .A(n_1172), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1179), .B(n_1228), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1217), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1230), .B(n_1160), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1228), .B(n_1206), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1248), .B(n_1218), .Y(n_1297) );
OAI221xp5_ASAP7_75t_L g1298 ( .A1(n_1246), .A2(n_1205), .B1(n_1163), .B2(n_1168), .C(n_1146), .Y(n_1298) );
INVx2_ASAP7_75t_L g1299 ( .A(n_1242), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1291), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1291), .Y(n_1301) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1295), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1294), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1248), .B(n_1252), .Y(n_1304) );
NAND4xp25_ASAP7_75t_SL g1305 ( .A(n_1246), .B(n_1207), .C(n_1237), .D(n_1206), .Y(n_1305) );
INVxp67_ASAP7_75t_SL g1306 ( .A(n_1267), .Y(n_1306) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_1270), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1296), .B(n_1226), .Y(n_1308) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1283), .B(n_1211), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1279), .B(n_1226), .Y(n_1310) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_1243), .B(n_1231), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_1286), .B(n_1250), .Y(n_1312) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1286), .B(n_1212), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1253), .B(n_1226), .Y(n_1314) );
NOR2x1_ASAP7_75t_L g1315 ( .A(n_1270), .B(n_1210), .Y(n_1315) );
OR2x2_ASAP7_75t_L g1316 ( .A(n_1253), .B(n_1145), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1279), .B(n_1229), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1318 ( .A(n_1255), .B(n_1145), .Y(n_1318) );
NAND2xp5_ASAP7_75t_SL g1319 ( .A(n_1270), .B(n_1210), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1255), .B(n_1145), .Y(n_1320) );
AND2x4_ASAP7_75t_L g1321 ( .A(n_1272), .B(n_1235), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1275), .B(n_1229), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1250), .B(n_1212), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1275), .B(n_1229), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1272), .B(n_1204), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1272), .B(n_1204), .Y(n_1326) );
HB1xp67_ASAP7_75t_L g1327 ( .A(n_1295), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1289), .B(n_1234), .Y(n_1328) );
INVx1_ASAP7_75t_SL g1329 ( .A(n_1290), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1279), .B(n_1173), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1262), .B(n_1204), .Y(n_1331) );
OAI33xp33_ASAP7_75t_L g1332 ( .A1(n_1259), .A2(n_1234), .A3(n_1238), .B1(n_1198), .B2(n_1221), .B3(n_1200), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1279), .B(n_1173), .Y(n_1333) );
NAND2xp5_ASAP7_75t_SL g1334 ( .A(n_1270), .B(n_1155), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1262), .B(n_1202), .Y(n_1335) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_1289), .B(n_1173), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1272), .B(n_1173), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1293), .B(n_1166), .Y(n_1338) );
NAND2xp5_ASAP7_75t_SL g1339 ( .A(n_1285), .B(n_1155), .Y(n_1339) );
NAND2x1p5_ASAP7_75t_L g1340 ( .A(n_1280), .B(n_1189), .Y(n_1340) );
INVx3_ASAP7_75t_L g1341 ( .A(n_1256), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1266), .B(n_1202), .Y(n_1342) );
NAND2x1p5_ASAP7_75t_L g1343 ( .A(n_1280), .B(n_1189), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1312), .B(n_1274), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1345 ( .A(n_1304), .B(n_1274), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1300), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1304), .B(n_1251), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1300), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1301), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1323), .B(n_1245), .Y(n_1350) );
INVx2_ASAP7_75t_L g1351 ( .A(n_1299), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1297), .B(n_1278), .Y(n_1352) );
HB1xp67_ASAP7_75t_L g1353 ( .A(n_1302), .Y(n_1353) );
INVx3_ASAP7_75t_L g1354 ( .A(n_1307), .Y(n_1354) );
NAND2x1p5_ASAP7_75t_L g1355 ( .A(n_1315), .B(n_1285), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1297), .B(n_1251), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g1357 ( .A1(n_1305), .A2(n_1259), .B1(n_1263), .B2(n_1254), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1312), .B(n_1273), .Y(n_1358) );
AND2x2_ASAP7_75t_SL g1359 ( .A(n_1321), .B(n_1156), .Y(n_1359) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1322), .B(n_1282), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1361 ( .A(n_1322), .B(n_1273), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1362 ( .A(n_1307), .B(n_1290), .Y(n_1362) );
NOR2x1_ASAP7_75t_L g1363 ( .A(n_1315), .B(n_1281), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1324), .B(n_1284), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1324), .B(n_1247), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1366 ( .A(n_1313), .B(n_1240), .Y(n_1366) );
AOI22xp5_ASAP7_75t_L g1367 ( .A1(n_1305), .A2(n_1288), .B1(n_1254), .B2(n_1243), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1313), .B(n_1247), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1314), .B(n_1269), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1301), .Y(n_1370) );
NOR2xp33_ASAP7_75t_L g1371 ( .A(n_1311), .B(n_1221), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1309), .B(n_1260), .Y(n_1372) );
OR2x6_ASAP7_75t_L g1373 ( .A(n_1307), .B(n_1254), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1331), .B(n_1257), .Y(n_1374) );
OAI31xp33_ASAP7_75t_L g1375 ( .A1(n_1298), .A2(n_1146), .A3(n_1149), .B(n_1292), .Y(n_1375) );
CKINVDCx5p33_ASAP7_75t_R g1376 ( .A(n_1319), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1331), .B(n_1241), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1339), .B(n_1187), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1302), .B(n_1241), .Y(n_1379) );
NOR2xp33_ASAP7_75t_L g1380 ( .A(n_1334), .B(n_1187), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1327), .B(n_1244), .Y(n_1381) );
INVx1_ASAP7_75t_L g1382 ( .A(n_1303), .Y(n_1382) );
OR2x2_ASAP7_75t_L g1383 ( .A(n_1309), .B(n_1260), .Y(n_1383) );
OAI21xp33_ASAP7_75t_L g1384 ( .A1(n_1298), .A2(n_1254), .B(n_1293), .Y(n_1384) );
NAND2x1p5_ASAP7_75t_L g1385 ( .A(n_1329), .B(n_1280), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1353), .Y(n_1386) );
AOI22xp5_ASAP7_75t_L g1387 ( .A1(n_1357), .A2(n_1332), .B1(n_1288), .B2(n_1258), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1365), .B(n_1317), .Y(n_1388) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1361), .B(n_1328), .Y(n_1389) );
NAND2xp5_ASAP7_75t_L g1390 ( .A(n_1374), .B(n_1308), .Y(n_1390) );
INVx1_ASAP7_75t_SL g1391 ( .A(n_1363), .Y(n_1391) );
HB1xp67_ASAP7_75t_L g1392 ( .A(n_1366), .Y(n_1392) );
INVx2_ASAP7_75t_L g1393 ( .A(n_1351), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1374), .B(n_1308), .Y(n_1394) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1346), .Y(n_1395) );
INVx2_ASAP7_75t_SL g1396 ( .A(n_1355), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1360), .B(n_1317), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1364), .B(n_1317), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1350), .B(n_1308), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1348), .Y(n_1400) );
AOI221xp5_ASAP7_75t_L g1401 ( .A1(n_1384), .A2(n_1332), .B1(n_1277), .B2(n_1258), .C(n_1287), .Y(n_1401) );
OR2x2_ASAP7_75t_L g1402 ( .A(n_1345), .B(n_1328), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1350), .B(n_1314), .Y(n_1403) );
INVx2_ASAP7_75t_L g1404 ( .A(n_1349), .Y(n_1404) );
INVx2_ASAP7_75t_L g1405 ( .A(n_1370), .Y(n_1405) );
INVxp67_ASAP7_75t_L g1406 ( .A(n_1371), .Y(n_1406) );
AOI21xp33_ASAP7_75t_SL g1407 ( .A1(n_1375), .A2(n_1343), .B(n_1340), .Y(n_1407) );
NAND3xp33_ASAP7_75t_SL g1408 ( .A(n_1375), .B(n_1343), .C(n_1340), .Y(n_1408) );
NOR2xp33_ASAP7_75t_L g1409 ( .A(n_1344), .B(n_1203), .Y(n_1409) );
OAI21xp5_ASAP7_75t_L g1410 ( .A1(n_1355), .A2(n_1306), .B(n_1254), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1369), .B(n_1330), .Y(n_1411) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_1358), .B(n_1203), .Y(n_1412) );
AOI22xp5_ASAP7_75t_L g1413 ( .A1(n_1359), .A2(n_1287), .B1(n_1277), .B2(n_1269), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1352), .B(n_1330), .Y(n_1414) );
OR2x2_ASAP7_75t_L g1415 ( .A(n_1347), .B(n_1316), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1368), .B(n_1330), .Y(n_1416) );
INVxp67_ASAP7_75t_L g1417 ( .A(n_1392), .Y(n_1417) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1386), .Y(n_1418) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_1406), .B(n_1367), .Y(n_1419) );
INVx2_ASAP7_75t_L g1420 ( .A(n_1393), .Y(n_1420) );
INVxp67_ASAP7_75t_SL g1421 ( .A(n_1396), .Y(n_1421) );
OAI211xp5_ASAP7_75t_L g1422 ( .A1(n_1407), .A2(n_1376), .B(n_1380), .C(n_1378), .Y(n_1422) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1386), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1424 ( .A(n_1415), .B(n_1356), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1411), .B(n_1377), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1411), .B(n_1377), .Y(n_1426) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_1415), .B(n_1372), .Y(n_1427) );
AOI21xp33_ASAP7_75t_L g1428 ( .A1(n_1391), .A2(n_1379), .B(n_1381), .Y(n_1428) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_1408), .A2(n_1373), .B1(n_1326), .B2(n_1325), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1389), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1389), .B(n_1383), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1395), .Y(n_1432) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1395), .Y(n_1433) );
INVxp67_ASAP7_75t_L g1434 ( .A(n_1409), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1400), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1416), .B(n_1338), .Y(n_1436) );
AOI222xp33_ASAP7_75t_L g1437 ( .A1(n_1401), .A2(n_1333), .B1(n_1276), .B2(n_1310), .C1(n_1325), .C2(n_1326), .Y(n_1437) );
OAI31xp33_ASAP7_75t_L g1438 ( .A1(n_1396), .A2(n_1354), .A3(n_1362), .B(n_1329), .Y(n_1438) );
INVx1_ASAP7_75t_L g1439 ( .A(n_1400), .Y(n_1439) );
AOI222xp33_ASAP7_75t_L g1440 ( .A1(n_1417), .A2(n_1412), .B1(n_1410), .B2(n_1399), .C1(n_1394), .C2(n_1390), .Y(n_1440) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_1419), .A2(n_1387), .B1(n_1413), .B2(n_1403), .Y(n_1441) );
OAI22xp5_ASAP7_75t_L g1442 ( .A1(n_1429), .A2(n_1407), .B1(n_1387), .B2(n_1402), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1424), .Y(n_1443) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_1428), .A2(n_1416), .B1(n_1397), .B2(n_1398), .C(n_1410), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1424), .Y(n_1445) );
NAND2x1p5_ASAP7_75t_L g1446 ( .A(n_1431), .B(n_1354), .Y(n_1446) );
AOI21xp33_ASAP7_75t_SL g1447 ( .A1(n_1437), .A2(n_1373), .B(n_1402), .Y(n_1447) );
INVxp67_ASAP7_75t_L g1448 ( .A(n_1419), .Y(n_1448) );
AOI221x1_ASAP7_75t_L g1449 ( .A1(n_1418), .A2(n_1341), .B1(n_1405), .B2(n_1404), .C(n_1382), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1450 ( .A(n_1430), .B(n_1388), .Y(n_1450) );
AO22x1_ASAP7_75t_L g1451 ( .A1(n_1421), .A2(n_1362), .B1(n_1292), .B2(n_1306), .Y(n_1451) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1427), .Y(n_1452) );
NOR2xp33_ASAP7_75t_L g1453 ( .A(n_1434), .B(n_1388), .Y(n_1453) );
OAI21xp5_ASAP7_75t_L g1454 ( .A1(n_1429), .A2(n_1373), .B(n_1385), .Y(n_1454) );
XNOR2xp5_ASAP7_75t_L g1455 ( .A(n_1422), .B(n_1414), .Y(n_1455) );
OAI211xp5_ASAP7_75t_SL g1456 ( .A1(n_1448), .A2(n_1438), .B(n_1423), .C(n_1431), .Y(n_1456) );
AOI221xp5_ASAP7_75t_L g1457 ( .A1(n_1447), .A2(n_1439), .B1(n_1432), .B2(n_1435), .C(n_1433), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1443), .Y(n_1458) );
OAI221xp5_ASAP7_75t_SL g1459 ( .A1(n_1455), .A2(n_1426), .B1(n_1425), .B2(n_1320), .C(n_1316), .Y(n_1459) );
NAND5xp2_ASAP7_75t_L g1460 ( .A(n_1454), .B(n_1343), .C(n_1340), .D(n_1385), .E(n_1233), .Y(n_1460) );
AOI221xp5_ASAP7_75t_L g1461 ( .A1(n_1442), .A2(n_1436), .B1(n_1420), .B2(n_1397), .C(n_1398), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1441), .B(n_1414), .Y(n_1462) );
OAI211xp5_ASAP7_75t_SL g1463 ( .A1(n_1440), .A2(n_1276), .B(n_1420), .C(n_1341), .Y(n_1463) );
AOI22xp5_ASAP7_75t_L g1464 ( .A1(n_1444), .A2(n_1333), .B1(n_1310), .B2(n_1337), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1465 ( .A(n_1445), .B(n_1404), .Y(n_1465) );
OAI221xp5_ASAP7_75t_L g1466 ( .A1(n_1446), .A2(n_1405), .B1(n_1318), .B2(n_1320), .C(n_1340), .Y(n_1466) );
OAI211xp5_ASAP7_75t_SL g1467 ( .A1(n_1457), .A2(n_1452), .B(n_1453), .C(n_1450), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1462), .B(n_1451), .Y(n_1468) );
OAI321xp33_ASAP7_75t_L g1469 ( .A1(n_1456), .A2(n_1446), .A3(n_1343), .B1(n_1318), .B2(n_1342), .C(n_1335), .Y(n_1469) );
OAI211xp5_ASAP7_75t_L g1470 ( .A1(n_1461), .A2(n_1449), .B(n_1149), .C(n_1292), .Y(n_1470) );
NOR3xp33_ASAP7_75t_SL g1471 ( .A(n_1459), .B(n_1265), .C(n_1268), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1472 ( .A(n_1458), .B(n_1393), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1473 ( .A(n_1465), .B(n_1336), .Y(n_1473) );
AND2x4_ASAP7_75t_L g1474 ( .A(n_1468), .B(n_1464), .Y(n_1474) );
NOR3xp33_ASAP7_75t_L g1475 ( .A(n_1470), .B(n_1463), .C(n_1460), .Y(n_1475) );
NAND2xp5_ASAP7_75t_SL g1476 ( .A(n_1469), .B(n_1149), .Y(n_1476) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_1467), .B(n_1466), .Y(n_1477) );
NAND5xp2_ASAP7_75t_L g1478 ( .A(n_1471), .B(n_1271), .C(n_1249), .D(n_1261), .E(n_1264), .Y(n_1478) );
NOR2xp67_ASAP7_75t_L g1479 ( .A(n_1476), .B(n_1472), .Y(n_1479) );
NOR3xp33_ASAP7_75t_L g1480 ( .A(n_1477), .B(n_1473), .C(n_1170), .Y(n_1480) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1474), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1478), .Y(n_1482) );
NAND3xp33_ASAP7_75t_L g1483 ( .A(n_1481), .B(n_1475), .C(n_1220), .Y(n_1483) );
OAI22x1_ASAP7_75t_L g1484 ( .A1(n_1482), .A2(n_1164), .B1(n_1170), .B2(n_1165), .Y(n_1484) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1483), .Y(n_1485) );
OAI22xp5_ASAP7_75t_SL g1486 ( .A1(n_1485), .A2(n_1484), .B1(n_1480), .B2(n_1479), .Y(n_1486) );
AOI22xp5_ASAP7_75t_L g1487 ( .A1(n_1486), .A2(n_1220), .B1(n_1172), .B2(n_1164), .Y(n_1487) );
OAI21xp5_ASAP7_75t_L g1488 ( .A1(n_1487), .A2(n_1186), .B(n_1189), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_1488), .A2(n_1341), .B1(n_1310), .B2(n_1321), .Y(n_1489) );
endmodule