module real_jpeg_8336_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_1),
.A2(n_40),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_138)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_63),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_3),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_70),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_4),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_10),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_10),
.A2(n_53),
.B(n_65),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_10),
.A2(n_63),
.B1(n_69),
.B2(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_10),
.B(n_157),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_10),
.A2(n_38),
.B(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_10),
.B(n_38),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_210),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_10),
.A2(n_52),
.B(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_10),
.B(n_52),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_11),
.A2(n_63),
.B1(n_69),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_11),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_90),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_90),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_90),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_12),
.A2(n_63),
.B1(n_69),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_12),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_72),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_72),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_14),
.A2(n_63),
.B1(n_69),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_14),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_130),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_130),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_130),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_58),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_58),
.B1(n_63),
.B2(n_69),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_16),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_17),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_17),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_115),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_94),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_21),
.B(n_94),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_74),
.C(n_80),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_22),
.A2(n_23),
.B1(n_74),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_24),
.B(n_60),
.C(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_25),
.B(n_36),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_26),
.A2(n_33),
.B(n_34),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_26),
.A2(n_33),
.B1(n_83),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_26),
.A2(n_33),
.B1(n_193),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_33),
.B1(n_195),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_26),
.A2(n_33),
.B1(n_226),
.B2(n_241),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_27),
.A2(n_28),
.B1(n_138),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_27),
.A2(n_28),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_30),
.B1(n_42),
.B2(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_29),
.B(n_45),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_29),
.B(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_30),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_33),
.B(n_134),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_85),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_39),
.B1(n_51),
.B2(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_38),
.B(n_56),
.Y(n_238)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_39),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_44),
.B1(n_46),
.B2(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_41),
.A2(n_44),
.B1(n_78),
.B2(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_41),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_41),
.A2(n_44),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_41),
.A2(n_44),
.B1(n_201),
.B2(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_41),
.A2(n_44),
.B1(n_224),
.B2(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_41),
.A2(n_44),
.B1(n_160),
.B2(n_231),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_42),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_43),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_44),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_44),
.B(n_134),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_60),
.B1(n_61),
.B2(n_73),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_55),
.B1(n_57),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_55),
.B1(n_59),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_50),
.A2(n_55),
.B1(n_93),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_50),
.A2(n_55),
.B1(n_125),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_50),
.A2(n_55),
.B1(n_153),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_50),
.A2(n_55),
.B1(n_179),
.B2(n_233),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_67)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_55),
.B(n_134),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_67),
.B1(n_68),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_67),
.B1(n_71),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_62),
.A2(n_67),
.B1(n_89),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.Y(n_66)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_64),
.B(n_134),
.C(n_135),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_67),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_74),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_75),
.A2(n_76),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_77),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_80),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.C(n_91),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_84),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_86),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_111),
.B2(n_112),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_102),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_100),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_106),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_111),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_142),
.B(n_265),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_139),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_117),
.B(n_139),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.C(n_121),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_120),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_121),
.A2(n_122),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_126),
.C(n_131),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_129),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_136),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_184),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_166),
.B(n_183),
.Y(n_144)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_145),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_163),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_163),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_154),
.C(n_158),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_152),
.B1(n_158),
.B2(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_158),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_167),
.B(n_169),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_175),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_170),
.B(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_173),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.C(n_181),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_178),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_180),
.B(n_181),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_182),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_263),
.C(n_264),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_257),
.B(n_262),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_243),
.B(n_256),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_228),
.B(n_242),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_218),
.B(n_227),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_207),
.B(n_217),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_191),
.B(n_196),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_202),
.B2(n_206),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_197),
.B(n_206),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_202),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_219),
.B(n_220),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_221),
.B(n_229),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_223),
.CI(n_225),
.CON(n_221),
.SN(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_229),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_232),
.CI(n_235),
.CON(n_229),
.SN(n_229)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_236),
.B(n_240),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_245),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_253),
.C(n_254),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_258),
.B(n_259),
.Y(n_262)
);


endmodule