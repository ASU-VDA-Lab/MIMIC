module real_jpeg_14234_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_2),
.B(n_30),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_44),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_2),
.B(n_61),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_2),
.B(n_71),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_2),
.B(n_75),
.Y(n_271)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_5),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_5),
.B(n_30),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_5),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_5),
.B(n_61),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_5),
.B(n_75),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_52),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_6),
.B(n_34),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_30),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_6),
.B(n_44),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_6),
.B(n_61),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_6),
.B(n_26),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_6),
.B(n_71),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_6),
.B(n_75),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_7),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_44),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_7),
.B(n_71),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_7),
.B(n_61),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_7),
.B(n_26),
.Y(n_106)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_7),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_75),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_10),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_10),
.B(n_30),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_10),
.B(n_44),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_10),
.B(n_61),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_10),
.B(n_26),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_12),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_61),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_12),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_12),
.B(n_71),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_52),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_13),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_13),
.B(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_14),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_14),
.B(n_26),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_14),
.B(n_52),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_14),
.B(n_30),
.Y(n_148)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_168),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_166),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_19),
.B(n_129),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_84),
.C(n_99),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_20),
.B(n_84),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_63),
.B2(n_64),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_21),
.B(n_65),
.C(n_77),
.Y(n_165)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_40),
.C(n_57),
.Y(n_133)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_25),
.B(n_29),
.C(n_32),
.Y(n_164)
);

INVx5_ASAP7_75t_SL g186 ( 
.A(n_26),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_33),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_33),
.B(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_36),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_36),
.B(n_120),
.Y(n_257)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_55),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_43),
.B(n_51),
.C(n_53),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_44),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_47),
.A2(n_53),
.B1(n_106),
.B2(n_210),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_SL g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_49),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_49),
.B(n_108),
.Y(n_289)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_51),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_54),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_67),
.C(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_51),
.A2(n_54),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_51),
.B(n_259),
.Y(n_269)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_106),
.C(n_107),
.Y(n_105)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_60),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_58),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_62),
.B(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_77),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_74),
.C(n_76),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_69),
.A2(n_70),
.B1(n_180),
.B2(n_181),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_70),
.B(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_72),
.B(n_124),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_72),
.B(n_108),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_76),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_78),
.B(n_80),
.C(n_82),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_81),
.A2(n_82),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_81),
.A2(n_82),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_81),
.A2(n_82),
.B1(n_96),
.B2(n_116),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_82),
.B(n_96),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.C(n_94),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_85),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_89),
.B(n_94),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.C(n_93),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_90),
.A2(n_91),
.B1(n_93),
.B2(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_92),
.A2(n_158),
.B1(n_159),
.B2(n_162),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_92),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_92),
.A2(n_162),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_93),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.C(n_97),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_99),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_113),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_100),
.B(n_104),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_111),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_105),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_107),
.B(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_109),
.A2(n_111),
.B1(n_112),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_113),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.C(n_125),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_114),
.B(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_117),
.A2(n_118),
.B1(n_125),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_118),
.A2(n_119),
.B(n_122),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_120),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_124),
.B(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_125)
);

FAx1_ASAP7_75t_SL g178 ( 
.A(n_126),
.B(n_127),
.CI(n_128),
.CON(n_178),
.SN(n_178)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_165),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_145),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_144),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_143),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_148),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_163),
.B2(n_164),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_160),
.A2(n_161),
.B1(n_183),
.B2(n_184),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_183),
.C(n_185),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_196),
.B(n_327),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_194),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_170),
.B(n_194),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.C(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_171),
.B(n_173),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.C(n_190),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_202),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.C(n_182),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_177),
.A2(n_178),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_178),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_179),
.B(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_185),
.B(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_244),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_221),
.B(n_243),
.Y(n_198)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_199),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_219),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_219),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_207),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_204),
.B1(n_207),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_218),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_211),
.CI(n_218),
.CON(n_227),
.SN(n_227)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.C(n_216),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_212),
.A2(n_213),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_222),
.B(n_225),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.C(n_232),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_226),
.A2(n_227),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_227),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_228),
.A2(n_229),
.B1(n_232),
.B2(n_233),
.Y(n_323)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_234),
.B(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_236),
.B(n_237),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.C(n_241),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR3xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_325),
.C(n_326),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_319),
.B(n_324),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_304),
.B(n_318),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_274),
.B(n_303),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_261),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_249),
.B(n_261),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.C(n_258),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_250),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_300),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_252),
.CI(n_253),
.CON(n_250),
.SN(n_250)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_254),
.A2(n_255),
.B1(n_258),
.B2(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_268),
.B2(n_273),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_267),
.C(n_273),
.Y(n_305)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_297),
.B(n_302),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_287),
.B(n_296),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_291),
.B(n_295),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_289),
.B(n_290),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_305),
.B(n_306),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_310),
.B2(n_311),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_312),
.C(n_317),
.Y(n_320)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_316),
.B2(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_321),
.Y(n_324)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);


endmodule