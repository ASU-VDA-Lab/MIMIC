module fake_ibex_665_n_4247 (n_151, n_85, n_599, n_778, n_822, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_583, n_887, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_861, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_158, n_859, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_875, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_373, n_854, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_898, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_835, n_168, n_526, n_785, n_155, n_824, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_838, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_852, n_789, n_880, n_654, n_656, n_724, n_437, n_731, n_602, n_904, n_842, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_851, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_844, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_847, n_830, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_834, n_257, n_77, n_869, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_882, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_905, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_894, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_815, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_485, n_870, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_572, n_867, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_424, n_565, n_823, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_895, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_4247);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_583;
input n_887;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_861;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_158;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_875;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_854;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_851;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_844;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_847;
input n_830;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_869;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_882;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_815;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_867;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_424;
input n_565;
input n_823;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;

output n_4247;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_2017;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3272;
wire n_3255;
wire n_3674;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4179;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_1782;
wire n_963;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3904;
wire n_3135;
wire n_3440;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_2565;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_1981;
wire n_1195;
wire n_3353;
wire n_2918;
wire n_3976;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_3747;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3884;
wire n_3881;
wire n_3507;
wire n_3949;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1910;
wire n_1496;
wire n_2436;
wire n_1663;
wire n_2333;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_3711;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_3699;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3910;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3769;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_4067;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_971;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2928;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_1988;
wire n_1132;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2444;
wire n_1742;
wire n_2350;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_3241;
wire n_2746;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3733;
wire n_3626;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2573;
wire n_1793;
wire n_1237;
wire n_2424;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_3849;
wire n_965;
wire n_1109;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3529;
wire n_1711;
wire n_3222;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3855;
wire n_4033;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_4215;
wire n_2434;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_1115;
wire n_998;
wire n_1729;
wire n_1395;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_3460;
wire n_2905;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3646;
wire n_2635;
wire n_3477;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4077;
wire n_3897;
wire n_3074;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2654;
wire n_2463;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_2990;
wire n_3449;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2923;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1683;
wire n_1185;
wire n_3575;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_3284;
wire n_2524;
wire n_2875;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_3902;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_4133;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_3314;
wire n_2997;
wire n_991;
wire n_1349;
wire n_1223;
wire n_1331;
wire n_961;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4142;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3828;
wire n_3240;
wire n_3336;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2683;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1991;
wire n_1025;
wire n_1177;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_3356;
wire n_1191;
wire n_2004;
wire n_4099;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_2274;
wire n_2698;
wire n_3899;
wire n_1617;
wire n_1839;
wire n_3930;
wire n_4149;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3462;
wire n_3424;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1946;
wire n_1726;
wire n_3111;
wire n_1938;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_4068;
wire n_1063;
wire n_3021;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3647;
wire n_3623;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3928;
wire n_3349;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_2348;
wire n_2576;
wire n_2417;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_4229;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1433;
wire n_1314;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3648;
wire n_3234;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_946;
wire n_1586;
wire n_1542;
wire n_1362;
wire n_3497;
wire n_4178;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_3561;
wire n_956;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_3102;
wire n_2872;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_3305;
wire n_1635;
wire n_1572;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_3163;
wire n_2929;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1912;
wire n_1297;
wire n_1369;
wire n_3143;
wire n_3655;
wire n_1734;
wire n_3543;
wire n_3791;
wire n_3742;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_1811;
wire n_928;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3919;
wire n_3683;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_980;
wire n_1193;
wire n_3067;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3483;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1721;
wire n_1379;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1904;
wire n_1262;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_2357;
wire n_2653;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2961;
wire n_2770;
wire n_2704;
wire n_2996;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2749;
wire n_2378;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_1525;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

INVx2_ASAP7_75t_L g909 ( 
.A(n_452),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_835),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_213),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_793),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_434),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_666),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_115),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_851),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_880),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_45),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_413),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_891),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_8),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_366),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_812),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_212),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_898),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_671),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_30),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_204),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_393),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_301),
.Y(n_930)
);

CKINVDCx16_ASAP7_75t_R g931 ( 
.A(n_803),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_548),
.Y(n_932)
);

CKINVDCx14_ASAP7_75t_R g933 ( 
.A(n_10),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_227),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_194),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_810),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_82),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_149),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_333),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_12),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_366),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_525),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_881),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_569),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_802),
.Y(n_945)
);

CKINVDCx16_ASAP7_75t_R g946 ( 
.A(n_157),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_478),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_793),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_646),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_831),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_429),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_815),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_58),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_513),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_771),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_785),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_870),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_839),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_634),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_404),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_663),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_774),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_866),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_130),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_523),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_27),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_70),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_66),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_478),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_600),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_115),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_72),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_476),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_797),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_29),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_259),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_890),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_595),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_264),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_14),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_864),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_717),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_113),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_744),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_894),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_877),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_856),
.Y(n_987)
);

BUFx8_ASAP7_75t_SL g988 ( 
.A(n_788),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_685),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_39),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_861),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_765),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_872),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_833),
.Y(n_994)
);

CKINVDCx16_ASAP7_75t_R g995 ( 
.A(n_884),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_353),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_898),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_248),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_801),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_892),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_606),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_422),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_632),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_804),
.Y(n_1004)
);

CKINVDCx14_ASAP7_75t_R g1005 ( 
.A(n_791),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_454),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_44),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_501),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_830),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_522),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_673),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_539),
.Y(n_1012)
);

CKINVDCx14_ASAP7_75t_R g1013 ( 
.A(n_250),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_538),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_119),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_846),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_638),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_337),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_557),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_818),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_879),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_733),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_899),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_907),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_697),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_776),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_185),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_70),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_504),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_826),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_867),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_707),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_908),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_245),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_389),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_855),
.Y(n_1036)
);

CKINVDCx20_ASAP7_75t_R g1037 ( 
.A(n_365),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_188),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_23),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_761),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_741),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_147),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_347),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_40),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_552),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_170),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_431),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_521),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_610),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_707),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_729),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_895),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_628),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_601),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_896),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_826),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_653),
.Y(n_1057)
);

CKINVDCx20_ASAP7_75t_R g1058 ( 
.A(n_725),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_785),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_418),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_654),
.Y(n_1061)
);

CKINVDCx20_ASAP7_75t_R g1062 ( 
.A(n_120),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_710),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_203),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_485),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_364),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_187),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_136),
.Y(n_1068)
);

BUFx10_ASAP7_75t_L g1069 ( 
.A(n_577),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_759),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_841),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_405),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_711),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_508),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_822),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_873),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_538),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_878),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_818),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_519),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_19),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_347),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_702),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_448),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_415),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_378),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_798),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_389),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_862),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_811),
.Y(n_1090)
);

BUFx10_ASAP7_75t_L g1091 ( 
.A(n_528),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_158),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_231),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_640),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_658),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_140),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_676),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_198),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_140),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_61),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_490),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_96),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_624),
.Y(n_1103)
);

CKINVDCx20_ASAP7_75t_R g1104 ( 
.A(n_807),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_489),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_821),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_579),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_615),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_610),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_879),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_346),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_901),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_179),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_782),
.Y(n_1114)
);

INVxp67_ASAP7_75t_L g1115 ( 
.A(n_421),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_419),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_828),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_906),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_795),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_259),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_829),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_14),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_838),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_380),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_215),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_486),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_17),
.Y(n_1127)
);

BUFx10_ASAP7_75t_L g1128 ( 
.A(n_150),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_674),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_127),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_267),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_813),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_800),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_178),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_743),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_572),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_779),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_500),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_36),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_372),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_472),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_88),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_888),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_6),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_883),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_561),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_623),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_876),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_296),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_357),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_816),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_72),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_256),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_849),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_403),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_482),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_26),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_688),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_18),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_634),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_289),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_711),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_420),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_868),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_219),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_834),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_554),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_413),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_41),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_687),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_163),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_320),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_631),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_542),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_SL g1175 ( 
.A(n_306),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_25),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_827),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_715),
.Y(n_1178)
);

CKINVDCx16_ASAP7_75t_R g1179 ( 
.A(n_403),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_874),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_600),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_461),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_289),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_878),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_843),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_88),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_903),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_37),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_373),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_377),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_791),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_121),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_842),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_392),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_204),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_832),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_260),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_428),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_712),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_605),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_623),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_869),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_794),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_823),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_820),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_568),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_752),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_864),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_606),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_15),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_245),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_856),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_77),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_140),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_846),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_799),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_484),
.Y(n_1217)
);

CKINVDCx14_ASAP7_75t_R g1218 ( 
.A(n_805),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_478),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_860),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_133),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_161),
.Y(n_1222)
);

CKINVDCx16_ASAP7_75t_R g1223 ( 
.A(n_246),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_65),
.Y(n_1224)
);

BUFx2_ASAP7_75t_L g1225 ( 
.A(n_139),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_458),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_839),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_819),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_436),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_206),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_492),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_781),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_528),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_489),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_847),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_215),
.Y(n_1236)
);

BUFx5_ASAP7_75t_L g1237 ( 
.A(n_796),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_21),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_842),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_425),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_322),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_905),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_545),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_668),
.Y(n_1244)
);

CKINVDCx14_ASAP7_75t_R g1245 ( 
.A(n_825),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_393),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_806),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_713),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_593),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_857),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_625),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_614),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_534),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_498),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_13),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_850),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_190),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_95),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_701),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_401),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_814),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_792),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_651),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_572),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_594),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_635),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_198),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_680),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_528),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_89),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_896),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_368),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_309),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_395),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_90),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_808),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_696),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_422),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_806),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_181),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_863),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_377),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_353),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_344),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_845),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_252),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_886),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_512),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_103),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_875),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_905),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_459),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_824),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_134),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_168),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_114),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_829),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_871),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_293),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_523),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_245),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_378),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_188),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_213),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_786),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_750),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_615),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_854),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_771),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_570),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_54),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_628),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_510),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_552),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_754),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_608),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_844),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_897),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_56),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_412),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_858),
.Y(n_1321)
);

BUFx8_ASAP7_75t_SL g1322 ( 
.A(n_58),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_797),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_744),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_562),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_375),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_660),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_853),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_885),
.Y(n_1329)
);

HB1xp67_ASAP7_75t_L g1330 ( 
.A(n_110),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_904),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_490),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_817),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_852),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_840),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_789),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_505),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_355),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_899),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_130),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_475),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_343),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_782),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_882),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_467),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_154),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_848),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_160),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_890),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_141),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_190),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_458),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_43),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_749),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_572),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_557),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_859),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_53),
.Y(n_1358)
);

CKINVDCx16_ASAP7_75t_R g1359 ( 
.A(n_836),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_445),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_887),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_540),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_459),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_902),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_734),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_299),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_576),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_450),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_900),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_586),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_325),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_115),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_647),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_383),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_790),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_719),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_301),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_663),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_20),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_121),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_336),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_345),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_836),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_893),
.Y(n_1384)
);

CKINVDCx14_ASAP7_75t_R g1385 ( 
.A(n_825),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_377),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_3),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_467),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_113),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_22),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_394),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_161),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_706),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_257),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_271),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_641),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_820),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_787),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_889),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_88),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_658),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_238),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_566),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_837),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_625),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_289),
.Y(n_1406)
);

BUFx10_ASAP7_75t_L g1407 ( 
.A(n_284),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_349),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_614),
.Y(n_1409)
);

BUFx2_ASAP7_75t_SL g1410 ( 
.A(n_304),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_63),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_865),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_809),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_121),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_660),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_718),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_530),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_732),
.Y(n_1418)
);

INVx1_ASAP7_75t_SL g1419 ( 
.A(n_861),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_933),
.Y(n_1420)
);

CKINVDCx14_ASAP7_75t_R g1421 ( 
.A(n_933),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1322),
.Y(n_1422)
);

INVxp67_ASAP7_75t_SL g1423 ( 
.A(n_1039),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_L g1424 ( 
.A(n_1051),
.B(n_0),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1013),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_SL g1426 ( 
.A(n_1069),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1013),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1092),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1005),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_981),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_981),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1317),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1317),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_942),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1010),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_915),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1139),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1005),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1052),
.B(n_0),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1218),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1218),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1159),
.Y(n_1442)
);

INVxp67_ASAP7_75t_SL g1443 ( 
.A(n_1001),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_915),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_1037),
.Y(n_1445)
);

INVxp67_ASAP7_75t_SL g1446 ( 
.A(n_1001),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1237),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1245),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1037),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1161),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1346),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1107),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1062),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1089),
.B(n_0),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1237),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1113),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1062),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_944),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1385),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1127),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1149),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1225),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_988),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1126),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_992),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1237),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1313),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_988),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_946),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1149),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1330),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1179),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_918),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1223),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_940),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_941),
.Y(n_1476)
);

CKINVDCx20_ASAP7_75t_R g1477 ( 
.A(n_1198),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_953),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1198),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_954),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_969),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1219),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_R g1483 ( 
.A(n_911),
.B(n_1),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_970),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1294),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1219),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1383),
.B(n_1),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1230),
.Y(n_1488)
);

INVxp67_ASAP7_75t_SL g1489 ( 
.A(n_1027),
.Y(n_1489)
);

CKINVDCx20_ASAP7_75t_R g1490 ( 
.A(n_1230),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1027),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1241),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1086),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_913),
.Y(n_1494)
);

CKINVDCx20_ASAP7_75t_R g1495 ( 
.A(n_1241),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_976),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1273),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1273),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_919),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1283),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1283),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1086),
.Y(n_1502)
);

CKINVDCx16_ASAP7_75t_R g1503 ( 
.A(n_1069),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_978),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1316),
.Y(n_1505)
);

BUFx3_ASAP7_75t_L g1506 ( 
.A(n_992),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1374),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_983),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1012),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1237),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1018),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_921),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1041),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1035),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1316),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_924),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1097),
.B(n_2),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1038),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1237),
.Y(n_1519)
);

CKINVDCx16_ASAP7_75t_R g1520 ( 
.A(n_1069),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1042),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1043),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1054),
.Y(n_1523)
);

NOR2xp67_ASAP7_75t_L g1524 ( 
.A(n_1123),
.B(n_1135),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_927),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_929),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1064),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_930),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1374),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1065),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_932),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1072),
.Y(n_1532)
);

CKINVDCx16_ASAP7_75t_R g1533 ( 
.A(n_1091),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_928),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1074),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1406),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1115),
.Y(n_1537)
);

NOR2xp67_ASAP7_75t_L g1538 ( 
.A(n_1184),
.B(n_2),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1465),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1458),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1503),
.B(n_1091),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1420),
.B(n_1041),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1513),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1428),
.B(n_1091),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1428),
.B(n_931),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1489),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1430),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1427),
.B(n_934),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1458),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1489),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1447),
.A2(n_1466),
.B(n_1455),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1491),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1431),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1510),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1458),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1519),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1534),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1432),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1433),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1520),
.B(n_1128),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1443),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1434),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1458),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1493),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1502),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1502),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1435),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1437),
.Y(n_1569)
);

BUFx8_ASAP7_75t_L g1570 ( 
.A(n_1426),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1442),
.B(n_1450),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1446),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1451),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1473),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1423),
.B(n_935),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1533),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1423),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1475),
.Y(n_1578)
);

AND2x4_ASAP7_75t_L g1579 ( 
.A(n_1452),
.B(n_1263),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1421),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1476),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1478),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1456),
.B(n_1263),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1537),
.B(n_938),
.Y(n_1584)
);

BUFx8_ASAP7_75t_L g1585 ( 
.A(n_1426),
.Y(n_1585)
);

BUFx6f_ASAP7_75t_L g1586 ( 
.A(n_1480),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1481),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1494),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1484),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1496),
.Y(n_1590)
);

AND3x2_ASAP7_75t_L g1591 ( 
.A(n_1424),
.B(n_1175),
.C(n_1299),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1504),
.Y(n_1592)
);

AND3x2_ASAP7_75t_L g1593 ( 
.A(n_1439),
.B(n_996),
.C(n_909),
.Y(n_1593)
);

INVx3_ASAP7_75t_L g1594 ( 
.A(n_1508),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1509),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1511),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1425),
.B(n_939),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1499),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1512),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1464),
.B(n_947),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1514),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1518),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1429),
.Y(n_1603)
);

INVx6_ASAP7_75t_L g1604 ( 
.A(n_1524),
.Y(n_1604)
);

INVxp67_ASAP7_75t_L g1605 ( 
.A(n_1516),
.Y(n_1605)
);

NOR2x1_ASAP7_75t_L g1606 ( 
.A(n_1467),
.B(n_1102),
.Y(n_1606)
);

BUFx3_ASAP7_75t_L g1607 ( 
.A(n_1525),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1460),
.B(n_1462),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1521),
.Y(n_1609)
);

BUFx6f_ASAP7_75t_L g1610 ( 
.A(n_1522),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1523),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1527),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1471),
.B(n_1128),
.Y(n_1613)
);

OAI22x1_ASAP7_75t_R g1614 ( 
.A1(n_1436),
.A2(n_1406),
.B1(n_998),
.B2(n_979),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1530),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1532),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1438),
.B(n_995),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1535),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1526),
.B(n_1128),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1517),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1528),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1454),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1531),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1538),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1487),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1448),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1459),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1469),
.Y(n_1629)
);

BUFx6f_ASAP7_75t_L g1630 ( 
.A(n_1472),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1474),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1485),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1463),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1483),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1468),
.B(n_1102),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1444),
.B(n_960),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1422),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1445),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1449),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1453),
.Y(n_1640)
);

CKINVDCx8_ASAP7_75t_R g1641 ( 
.A(n_1457),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1461),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1470),
.Y(n_1643)
);

INVxp67_ASAP7_75t_L g1644 ( 
.A(n_1477),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1479),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1482),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1486),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1488),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1490),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1492),
.B(n_1163),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1495),
.B(n_964),
.Y(n_1651)
);

OA21x2_ASAP7_75t_L g1652 ( 
.A1(n_1497),
.A2(n_996),
.B(n_909),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1498),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1500),
.B(n_1236),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1501),
.B(n_1236),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1505),
.B(n_965),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1507),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1515),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1529),
.B(n_1359),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1536),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1489),
.Y(n_1661)
);

BUFx2_ASAP7_75t_L g1662 ( 
.A(n_1420),
.Y(n_1662)
);

INVx3_ASAP7_75t_L g1663 ( 
.A(n_1465),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1447),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1428),
.B(n_1236),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1465),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1489),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1465),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1489),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1420),
.B(n_966),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1489),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1465),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1447),
.A2(n_1081),
.B(n_1044),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1420),
.B(n_967),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1489),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1465),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1458),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1458),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1447),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1428),
.B(n_1300),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1489),
.Y(n_1681)
);

INVx3_ASAP7_75t_L g1682 ( 
.A(n_1465),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1465),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1428),
.B(n_1300),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1420),
.B(n_968),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1420),
.B(n_971),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1503),
.B(n_1300),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1428),
.B(n_1407),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1489),
.Y(n_1689)
);

INVx6_ASAP7_75t_L g1690 ( 
.A(n_1465),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1465),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1489),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1428),
.B(n_1407),
.Y(n_1693)
);

INVx3_ASAP7_75t_L g1694 ( 
.A(n_1465),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1465),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1420),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1465),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1465),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1420),
.B(n_972),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1420),
.B(n_1163),
.Y(n_1700)
);

AOI22x1_ASAP7_75t_SL g1701 ( 
.A1(n_1436),
.A2(n_1020),
.B1(n_1025),
.B2(n_1017),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1489),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1420),
.B(n_973),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1489),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1489),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1465),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1420),
.B(n_975),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1458),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1420),
.B(n_980),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1465),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1420),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1458),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1465),
.Y(n_1713)
);

BUFx6f_ASAP7_75t_L g1714 ( 
.A(n_1458),
.Y(n_1714)
);

OR2x6_ASAP7_75t_L g1715 ( 
.A(n_1428),
.B(n_1410),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1489),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1489),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1465),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1489),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1447),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1465),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1465),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1503),
.B(n_990),
.Y(n_1723)
);

BUFx2_ASAP7_75t_L g1724 ( 
.A(n_1420),
.Y(n_1724)
);

NOR2x1_ASAP7_75t_L g1725 ( 
.A(n_1464),
.B(n_1167),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1420),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1489),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1465),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1465),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1458),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1503),
.B(n_1006),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1489),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1420),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1620),
.B(n_1007),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1613),
.B(n_1044),
.Y(n_1735)
);

AOI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1545),
.A2(n_1014),
.B1(n_1015),
.B2(n_1008),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1665),
.B(n_1081),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1563),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1715),
.B(n_914),
.Y(n_1739)
);

BUFx6f_ASAP7_75t_L g1740 ( 
.A(n_1607),
.Y(n_1740)
);

BUFx10_ASAP7_75t_L g1741 ( 
.A(n_1715),
.Y(n_1741)
);

BUFx10_ASAP7_75t_L g1742 ( 
.A(n_1635),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1626),
.B(n_1019),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1570),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1673),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1549),
.B(n_1028),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1574),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1594),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1680),
.B(n_1222),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1636),
.B(n_937),
.C(n_922),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1684),
.B(n_1222),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1602),
.B(n_1029),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1568),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1569),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1670),
.B(n_1046),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1574),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1558),
.B(n_1075),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1688),
.A2(n_1048),
.B1(n_1049),
.B2(n_1047),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1586),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1634),
.A2(n_1066),
.B1(n_1067),
.B2(n_1060),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1573),
.Y(n_1761)
);

INVx8_ASAP7_75t_L g1762 ( 
.A(n_1576),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1693),
.B(n_1229),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1586),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1690),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1610),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1674),
.B(n_1068),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1685),
.B(n_1077),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_L g1769 ( 
.A1(n_1547),
.A2(n_1181),
.B1(n_1214),
.B2(n_1174),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1610),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1634),
.A2(n_1084),
.B1(n_1085),
.B2(n_1080),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1686),
.B(n_1088),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1616),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1570),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1616),
.Y(n_1775)
);

NAND2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1588),
.B(n_1598),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1585),
.B(n_1017),
.Y(n_1777)
);

INVxp67_ASAP7_75t_SL g1778 ( 
.A(n_1711),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1552),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1699),
.B(n_1093),
.Y(n_1780)
);

INVx2_ASAP7_75t_SL g1781 ( 
.A(n_1662),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1662),
.B(n_1696),
.Y(n_1782)
);

INVx1_ASAP7_75t_SL g1783 ( 
.A(n_1696),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1539),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1573),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1544),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1666),
.Y(n_1787)
);

AND2x6_ASAP7_75t_L g1788 ( 
.A(n_1619),
.B(n_1214),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1566),
.B(n_1099),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1548),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1724),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1668),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_SL g1793 ( 
.A(n_1638),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_SL g1794 ( 
.A(n_1597),
.B(n_1229),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1672),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1567),
.B(n_1100),
.Y(n_1796)
);

OR2x6_ASAP7_75t_L g1797 ( 
.A(n_1598),
.B(n_1409),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1554),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1559),
.Y(n_1799)
);

INVx6_ASAP7_75t_L g1800 ( 
.A(n_1585),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1551),
.A2(n_1325),
.B1(n_1340),
.B2(n_1289),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1703),
.B(n_1101),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1560),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1724),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1661),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1541),
.Y(n_1806)
);

INVx3_ASAP7_75t_L g1807 ( 
.A(n_1663),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1683),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1726),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1709),
.B(n_1105),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1695),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1667),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1623),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1669),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1671),
.Y(n_1815)
);

BUFx10_ASAP7_75t_L g1816 ( 
.A(n_1635),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1700),
.B(n_916),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1675),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1681),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1689),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1676),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1692),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_SL g1823 ( 
.A(n_1577),
.B(n_1260),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1702),
.Y(n_1824)
);

AND2x6_ASAP7_75t_L g1825 ( 
.A(n_1704),
.B(n_1705),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1698),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1706),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1621),
.Y(n_1828)
);

BUFx4f_ASAP7_75t_L g1829 ( 
.A(n_1630),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1546),
.B(n_951),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_L g1831 ( 
.A(n_1584),
.B(n_1109),
.C(n_1108),
.Y(n_1831)
);

HB1xp67_ASAP7_75t_L g1832 ( 
.A(n_1733),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1716),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1710),
.Y(n_1834)
);

CKINVDCx20_ASAP7_75t_R g1835 ( 
.A(n_1621),
.Y(n_1835)
);

BUFx10_ASAP7_75t_L g1836 ( 
.A(n_1630),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1623),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1682),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1717),
.A2(n_1325),
.B1(n_1340),
.B2(n_1289),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1713),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1719),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1562),
.B(n_1116),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1727),
.A2(n_1732),
.B1(n_1572),
.B2(n_1575),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1718),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1707),
.B(n_1120),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1700),
.B(n_1122),
.Y(n_1846)
);

OR2x6_ASAP7_75t_L g1847 ( 
.A(n_1654),
.B(n_1020),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1721),
.Y(n_1848)
);

OAI22x1_ASAP7_75t_L g1849 ( 
.A1(n_1644),
.A2(n_1125),
.B1(n_1130),
.B2(n_1124),
.Y(n_1849)
);

INVx2_ASAP7_75t_SL g1850 ( 
.A(n_1543),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1600),
.B(n_1260),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1581),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1728),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1650),
.Y(n_1854)
);

INVx3_ASAP7_75t_L g1855 ( 
.A(n_1691),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1582),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1587),
.Y(n_1857)
);

INVx4_ASAP7_75t_L g1858 ( 
.A(n_1694),
.Y(n_1858)
);

NOR2x1p5_ASAP7_75t_L g1859 ( 
.A(n_1639),
.B(n_1131),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1543),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1590),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1596),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1608),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1697),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1628),
.B(n_1134),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1601),
.Y(n_1866)
);

INVx4_ASAP7_75t_L g1867 ( 
.A(n_1722),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1729),
.Y(n_1868)
);

AO22x1_ASAP7_75t_L g1869 ( 
.A1(n_1606),
.A2(n_1138),
.B1(n_1141),
.B2(n_1136),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1571),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1725),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1578),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1589),
.Y(n_1873)
);

OR2x6_ASAP7_75t_L g1874 ( 
.A(n_1637),
.B(n_1025),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1553),
.B(n_1144),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1592),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1622),
.B(n_1275),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1723),
.A2(n_1070),
.B1(n_1104),
.B2(n_1058),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1595),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1565),
.B(n_1150),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1627),
.B(n_1152),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1731),
.B(n_1075),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_L g1883 ( 
.A(n_1617),
.B(n_1155),
.C(n_1153),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1580),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1624),
.B(n_1156),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1609),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1611),
.B(n_1612),
.Y(n_1887)
);

BUFx3_ASAP7_75t_L g1888 ( 
.A(n_1580),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1603),
.B(n_1165),
.Y(n_1889)
);

OR2x6_ASAP7_75t_L g1890 ( 
.A(n_1637),
.B(n_1058),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1615),
.B(n_1168),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1618),
.Y(n_1892)
);

OR2x6_ASAP7_75t_L g1893 ( 
.A(n_1650),
.B(n_1070),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1608),
.B(n_1169),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1579),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1579),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1583),
.B(n_1172),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1555),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1583),
.B(n_1338),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1652),
.A2(n_1379),
.B1(n_1370),
.B2(n_1096),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1599),
.B(n_1399),
.Y(n_1901)
);

INVx5_ASAP7_75t_L g1902 ( 
.A(n_1540),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1593),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1604),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1555),
.Y(n_1905)
);

BUFx3_ASAP7_75t_L g1906 ( 
.A(n_1633),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1557),
.Y(n_1907)
);

INVxp67_ASAP7_75t_SL g1908 ( 
.A(n_1605),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1557),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1664),
.Y(n_1910)
);

AND2x2_ASAP7_75t_SL g1911 ( 
.A(n_1659),
.B(n_1338),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1629),
.B(n_1395),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1679),
.Y(n_1913)
);

OR2x6_ASAP7_75t_L g1914 ( 
.A(n_1658),
.B(n_1104),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1720),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1542),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1632),
.A2(n_1098),
.B1(n_1111),
.B2(n_1082),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1540),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_SL g1919 ( 
.A(n_1638),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1561),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1687),
.B(n_1186),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1591),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1631),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1651),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1656),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1655),
.A2(n_1146),
.B1(n_1157),
.B2(n_1140),
.Y(n_1926)
);

AND2x6_ASAP7_75t_L g1927 ( 
.A(n_1643),
.B(n_1395),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1625),
.B(n_1408),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1642),
.Y(n_1929)
);

BUFx3_ASAP7_75t_L g1930 ( 
.A(n_1642),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1647),
.B(n_945),
.Y(n_1931)
);

OR2x6_ASAP7_75t_L g1932 ( 
.A(n_1645),
.B(n_1166),
.Y(n_1932)
);

AND3x2_ASAP7_75t_L g1933 ( 
.A(n_1640),
.B(n_1298),
.C(n_1166),
.Y(n_1933)
);

INVx5_ASAP7_75t_L g1934 ( 
.A(n_1550),
.Y(n_1934)
);

INVx5_ASAP7_75t_L g1935 ( 
.A(n_1556),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1564),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1564),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1677),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1677),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1641),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1678),
.Y(n_1941)
);

OR2x6_ASAP7_75t_L g1942 ( 
.A(n_1646),
.B(n_1298),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1648),
.B(n_1188),
.Y(n_1943)
);

AND2x2_ASAP7_75t_SL g1944 ( 
.A(n_1653),
.B(n_1171),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1678),
.Y(n_1945)
);

AOI22xp33_ASAP7_75t_L g1946 ( 
.A1(n_1643),
.A2(n_1183),
.B1(n_1189),
.B2(n_1176),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1708),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1646),
.B(n_1417),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1708),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1712),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1712),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1714),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1649),
.B(n_1190),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1657),
.B(n_1195),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1660),
.B(n_1197),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1714),
.B(n_1414),
.Y(n_1956)
);

OAI21xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1614),
.A2(n_1194),
.B(n_1192),
.Y(n_1957)
);

XOR2xp5_ASAP7_75t_L g1958 ( 
.A(n_1701),
.B(n_1305),
.Y(n_1958)
);

BUFx6f_ASAP7_75t_L g1959 ( 
.A(n_1730),
.Y(n_1959)
);

BUFx6f_ASAP7_75t_L g1960 ( 
.A(n_1701),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1613),
.B(n_1206),
.Y(n_1961)
);

INVx3_ASAP7_75t_L g1962 ( 
.A(n_1573),
.Y(n_1962)
);

INVx2_ASAP7_75t_SL g1963 ( 
.A(n_1662),
.Y(n_1963)
);

AND2x2_ASAP7_75t_SL g1964 ( 
.A(n_1723),
.B(n_1200),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1673),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1620),
.B(n_1211),
.Y(n_1966)
);

INVx2_ASAP7_75t_SL g1967 ( 
.A(n_1662),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1620),
.B(n_1213),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1594),
.B(n_1217),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1673),
.Y(n_1970)
);

AND2x6_ASAP7_75t_L g1971 ( 
.A(n_1613),
.B(n_944),
.Y(n_1971)
);

NAND2xp33_ASAP7_75t_R g1972 ( 
.A(n_1598),
.B(n_1221),
.Y(n_1972)
);

INVx2_ASAP7_75t_SL g1973 ( 
.A(n_1662),
.Y(n_1973)
);

AND2x6_ASAP7_75t_L g1974 ( 
.A(n_1613),
.B(n_944),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1558),
.B(n_1002),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1673),
.Y(n_1976)
);

NOR2x1p5_ASAP7_75t_L g1977 ( 
.A(n_1576),
.B(n_1224),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1594),
.B(n_1233),
.Y(n_1978)
);

INVx2_ASAP7_75t_SL g1979 ( 
.A(n_1662),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1563),
.Y(n_1980)
);

NAND2xp33_ASAP7_75t_L g1981 ( 
.A(n_1620),
.B(n_1237),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1673),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1673),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1563),
.Y(n_1984)
);

INVx2_ASAP7_75t_SL g1985 ( 
.A(n_1662),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1607),
.Y(n_1986)
);

AND3x2_ASAP7_75t_L g1987 ( 
.A(n_1723),
.B(n_1305),
.C(n_1003),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1563),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1673),
.Y(n_1989)
);

BUFx2_ASAP7_75t_L g1990 ( 
.A(n_1558),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1673),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1573),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1734),
.B(n_1240),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1805),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1809),
.B(n_1258),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1966),
.B(n_1246),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1968),
.B(n_1249),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1812),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1990),
.B(n_1252),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1990),
.B(n_1253),
.Y(n_2000)
);

INVx3_ASAP7_75t_L g2001 ( 
.A(n_1898),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1783),
.B(n_1399),
.Y(n_2002)
);

BUFx6f_ASAP7_75t_L g2003 ( 
.A(n_1959),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_1825),
.A2(n_1255),
.B1(n_1257),
.B2(n_1254),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1791),
.A2(n_1269),
.B1(n_1278),
.B2(n_1267),
.Y(n_2005)
);

NAND2x1_ASAP7_75t_L g2006 ( 
.A(n_1825),
.B(n_944),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1870),
.A2(n_1282),
.B1(n_1286),
.B2(n_1280),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1781),
.B(n_1292),
.Y(n_2008)
);

NAND2xp33_ASAP7_75t_L g2009 ( 
.A(n_1825),
.B(n_1314),
.Y(n_2009)
);

AOI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1924),
.A2(n_1303),
.B1(n_1304),
.B2(n_1296),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1804),
.Y(n_2011)
);

BUFx3_ASAP7_75t_L g2012 ( 
.A(n_1762),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1746),
.B(n_1310),
.Y(n_2013)
);

INVx2_ASAP7_75t_SL g2014 ( 
.A(n_1828),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1755),
.B(n_1319),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1963),
.B(n_1356),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1767),
.B(n_1320),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1967),
.B(n_1358),
.Y(n_2018)
);

HB1xp67_ASAP7_75t_L g2019 ( 
.A(n_1804),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1782),
.B(n_1399),
.Y(n_2020)
);

NOR2xp33_ASAP7_75t_SL g2021 ( 
.A(n_1964),
.B(n_1774),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_L g2022 ( 
.A(n_1830),
.B(n_1326),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1913),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1973),
.B(n_1979),
.Y(n_2024)
);

INVx4_ASAP7_75t_L g2025 ( 
.A(n_1813),
.Y(n_2025)
);

CKINVDCx5p33_ASAP7_75t_R g2026 ( 
.A(n_1835),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_1925),
.B(n_1332),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1985),
.B(n_1352),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1814),
.Y(n_2029)
);

BUFx2_ASAP7_75t_L g2030 ( 
.A(n_1832),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1925),
.B(n_1342),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1768),
.B(n_1345),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1750),
.A2(n_1351),
.B1(n_1353),
.B2(n_1350),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1742),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1772),
.B(n_1780),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1815),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_SL g2037 ( 
.A(n_1744),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1818),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1819),
.Y(n_2039)
);

BUFx3_ASAP7_75t_L g2040 ( 
.A(n_1800),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1820),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1863),
.B(n_1355),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_1742),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1802),
.B(n_1360),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1810),
.B(n_1362),
.Y(n_2045)
);

AOI22xp33_ASAP7_75t_L g2046 ( 
.A1(n_1743),
.A2(n_1366),
.B1(n_1367),
.B2(n_1363),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1923),
.A2(n_1737),
.B1(n_1751),
.B2(n_1749),
.Y(n_2047)
);

INVx3_ASAP7_75t_L g2048 ( 
.A(n_1761),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1975),
.B(n_1368),
.Y(n_2049)
);

NAND2xp33_ASAP7_75t_L g2050 ( 
.A(n_1788),
.B(n_1372),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1822),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1739),
.B(n_1371),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1959),
.Y(n_2053)
);

NOR2xp33_ASAP7_75t_L g2054 ( 
.A(n_1778),
.B(n_1381),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1873),
.Y(n_2055)
);

INVx2_ASAP7_75t_SL g2056 ( 
.A(n_1816),
.Y(n_2056)
);

NAND2xp33_ASAP7_75t_L g2057 ( 
.A(n_1788),
.B(n_1386),
.Y(n_2057)
);

OR2x2_ASAP7_75t_L g2058 ( 
.A(n_1797),
.B(n_1034),
.Y(n_2058)
);

NAND2xp33_ASAP7_75t_SL g2059 ( 
.A(n_1740),
.B(n_1387),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1879),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1776),
.B(n_1394),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1901),
.B(n_1402),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1886),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1739),
.B(n_1142),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1824),
.Y(n_2065)
);

INVx2_ASAP7_75t_SL g2066 ( 
.A(n_1816),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1889),
.B(n_1182),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1905),
.Y(n_2068)
);

NAND3xp33_ASAP7_75t_L g2069 ( 
.A(n_1845),
.B(n_912),
.C(n_910),
.Y(n_2069)
);

OR2x6_ASAP7_75t_L g2070 ( 
.A(n_1800),
.B(n_950),
.Y(n_2070)
);

INVxp67_ASAP7_75t_L g2071 ( 
.A(n_1972),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1882),
.B(n_1411),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1833),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1841),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1740),
.B(n_917),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1757),
.B(n_920),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1986),
.B(n_923),
.Y(n_2077)
);

NOR2xp33_ASAP7_75t_L g2078 ( 
.A(n_1920),
.B(n_925),
.Y(n_2078)
);

AOI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_1878),
.A2(n_1946),
.B1(n_1771),
.B2(n_1760),
.C(n_1894),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_1986),
.B(n_926),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1872),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1736),
.B(n_1758),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_SL g2083 ( 
.A(n_1831),
.B(n_936),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1887),
.B(n_1209),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1891),
.B(n_1210),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1907),
.Y(n_2086)
);

NAND2xp33_ASAP7_75t_L g2087 ( 
.A(n_1788),
.B(n_943),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1842),
.B(n_1403),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_1847),
.B(n_982),
.Y(n_2089)
);

INVx2_ASAP7_75t_SL g2090 ( 
.A(n_1884),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1876),
.B(n_1231),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1961),
.B(n_948),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1892),
.B(n_1234),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1909),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1763),
.A2(n_1243),
.B1(n_1264),
.B2(n_1238),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1738),
.B(n_1265),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_L g2097 ( 
.A(n_1875),
.B(n_952),
.C(n_949),
.Y(n_2097)
);

NOR2x1p5_ASAP7_75t_L g2098 ( 
.A(n_1940),
.B(n_997),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1850),
.B(n_956),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1753),
.B(n_1270),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1754),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1888),
.Y(n_2102)
);

BUFx3_ASAP7_75t_L g2103 ( 
.A(n_1813),
.Y(n_2103)
);

BUFx12f_ASAP7_75t_SL g2104 ( 
.A(n_1874),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1910),
.Y(n_2105)
);

BUFx12f_ASAP7_75t_SL g2106 ( 
.A(n_1890),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1915),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_1735),
.A2(n_1274),
.B1(n_1284),
.B2(n_1272),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1980),
.B(n_1288),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1984),
.B(n_1295),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1944),
.B(n_1419),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1988),
.B(n_1302),
.Y(n_2112)
);

NOR2xp33_ASAP7_75t_L g2113 ( 
.A(n_1860),
.B(n_958),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1856),
.Y(n_2114)
);

INVxp67_ASAP7_75t_L g2115 ( 
.A(n_1777),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1857),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_1908),
.B(n_959),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1852),
.B(n_1307),
.Y(n_2118)
);

NOR2x1_ASAP7_75t_L g2119 ( 
.A(n_1883),
.B(n_1311),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1861),
.B(n_1348),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1906),
.B(n_957),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_1916),
.B(n_962),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1862),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1752),
.B(n_1400),
.Y(n_2124)
);

NAND2x1p5_ASAP7_75t_L g2125 ( 
.A(n_1829),
.B(n_1837),
.Y(n_2125)
);

NOR3xp33_ASAP7_75t_L g2126 ( 
.A(n_1957),
.B(n_1869),
.C(n_1854),
.Y(n_2126)
);

AOI22xp33_ASAP7_75t_L g2127 ( 
.A1(n_1900),
.A2(n_1380),
.B1(n_1382),
.B2(n_1377),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1969),
.B(n_974),
.Y(n_2128)
);

O2A1O1Ixp33_ASAP7_75t_L g2129 ( 
.A1(n_1823),
.A2(n_1390),
.B(n_1391),
.C(n_1389),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1962),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_1971),
.A2(n_1392),
.B1(n_1226),
.B2(n_1301),
.Y(n_2131)
);

AOI22xp33_ASAP7_75t_L g2132 ( 
.A1(n_1971),
.A2(n_1226),
.B1(n_1301),
.B2(n_1045),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1866),
.Y(n_2133)
);

AND2x2_ASAP7_75t_SL g2134 ( 
.A(n_1960),
.B(n_950),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1978),
.B(n_977),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_1932),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1748),
.Y(n_2137)
);

NOR2xp33_ASAP7_75t_L g2138 ( 
.A(n_1846),
.B(n_985),
.Y(n_2138)
);

AND2x4_ASAP7_75t_L g2139 ( 
.A(n_1977),
.B(n_963),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1741),
.B(n_989),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_1741),
.B(n_991),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1931),
.B(n_1178),
.Y(n_2142)
);

A2O1A1Ixp33_ASAP7_75t_L g2143 ( 
.A1(n_1880),
.A2(n_986),
.B(n_987),
.C(n_984),
.Y(n_2143)
);

OR2x6_ASAP7_75t_L g2144 ( 
.A(n_1890),
.B(n_1009),
.Y(n_2144)
);

CKINVDCx5p33_ASAP7_75t_R g2145 ( 
.A(n_1793),
.Y(n_2145)
);

O2A1O1Ixp33_ASAP7_75t_L g2146 ( 
.A1(n_1897),
.A2(n_1899),
.B(n_1789),
.C(n_1796),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1917),
.B(n_1790),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1798),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1799),
.B(n_999),
.Y(n_2149)
);

INVx8_ASAP7_75t_L g2150 ( 
.A(n_1971),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1779),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1928),
.B(n_1865),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_1921),
.B(n_1004),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1803),
.B(n_1011),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1895),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1817),
.B(n_1016),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_1932),
.Y(n_2157)
);

INVxp33_ASAP7_75t_L g2158 ( 
.A(n_1943),
.Y(n_2158)
);

OR2x2_ASAP7_75t_L g2159 ( 
.A(n_1893),
.B(n_1378),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1955),
.B(n_1022),
.Y(n_2160)
);

INVxp67_ASAP7_75t_L g2161 ( 
.A(n_1942),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1784),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_1992),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1896),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1786),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1817),
.B(n_1021),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1787),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1974),
.B(n_1023),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1974),
.B(n_1030),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1931),
.B(n_1031),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1792),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1795),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1808),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_1881),
.A2(n_1033),
.B1(n_1036),
.B2(n_1032),
.Y(n_2174)
);

BUFx2_ASAP7_75t_L g2175 ( 
.A(n_1942),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1811),
.Y(n_2176)
);

NOR2xp33_ASAP7_75t_L g2177 ( 
.A(n_1953),
.B(n_1954),
.Y(n_2177)
);

AND2x6_ASAP7_75t_L g2178 ( 
.A(n_1903),
.B(n_1045),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1974),
.B(n_1040),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1769),
.B(n_1055),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_1836),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1826),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_SL g2183 ( 
.A(n_1801),
.B(n_1056),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1893),
.B(n_1057),
.Y(n_2184)
);

BUFx3_ASAP7_75t_L g2185 ( 
.A(n_1836),
.Y(n_2185)
);

NOR2xp67_ASAP7_75t_SL g2186 ( 
.A(n_1922),
.B(n_1063),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1851),
.B(n_1071),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1869),
.B(n_1073),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1827),
.Y(n_2189)
);

INVxp67_ASAP7_75t_L g2190 ( 
.A(n_1914),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_1914),
.B(n_1076),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_1834),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1840),
.Y(n_2193)
);

BUFx3_ASAP7_75t_L g2194 ( 
.A(n_1929),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_1927),
.A2(n_1226),
.B1(n_1301),
.B2(n_1045),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1844),
.Y(n_2196)
);

NAND2xp33_ASAP7_75t_SL g2197 ( 
.A(n_1859),
.B(n_1413),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_1794),
.B(n_1079),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1839),
.B(n_1083),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1885),
.B(n_1087),
.Y(n_2200)
);

BUFx3_ASAP7_75t_L g2201 ( 
.A(n_1930),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1926),
.B(n_1095),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_L g2203 ( 
.A1(n_1745),
.A2(n_1024),
.B(n_1009),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_SL g2204 ( 
.A(n_1956),
.B(n_1106),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_1911),
.B(n_1110),
.Y(n_2205)
);

NOR2xp67_ASAP7_75t_L g2206 ( 
.A(n_1871),
.B(n_3),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1848),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_1853),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_1912),
.A2(n_1877),
.B1(n_1849),
.B2(n_1981),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_1838),
.Y(n_2210)
);

NAND2xp33_ASAP7_75t_L g2211 ( 
.A(n_1965),
.B(n_1112),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_SL g2212 ( 
.A(n_1858),
.B(n_1114),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_1867),
.B(n_1117),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1806),
.B(n_1118),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1970),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_1948),
.B(n_993),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1807),
.B(n_1121),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1987),
.B(n_1129),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1785),
.Y(n_2219)
);

NAND2xp33_ASAP7_75t_L g2220 ( 
.A(n_1976),
.B(n_1132),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1821),
.B(n_1133),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1855),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1864),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1747),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_1756),
.B(n_1137),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1759),
.Y(n_2226)
);

NAND2xp33_ASAP7_75t_L g2227 ( 
.A(n_1982),
.B(n_1983),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_1868),
.A2(n_1148),
.B1(n_1151),
.B2(n_1143),
.Y(n_2228)
);

INVx3_ASAP7_75t_L g2229 ( 
.A(n_1764),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1989),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1765),
.B(n_1154),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_1919),
.Y(n_2232)
);

A2O1A1Ixp33_ASAP7_75t_L g2233 ( 
.A1(n_1991),
.A2(n_1000),
.B(n_1026),
.C(n_994),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1765),
.B(n_1158),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1766),
.B(n_1770),
.Y(n_2235)
);

NOR2xp33_ASAP7_75t_L g2236 ( 
.A(n_1904),
.B(n_1160),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_1773),
.B(n_1164),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1775),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1902),
.B(n_1170),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1902),
.B(n_1173),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_1902),
.B(n_1187),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1934),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1934),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_1933),
.B(n_1191),
.Y(n_2244)
);

INVx8_ASAP7_75t_L g2245 ( 
.A(n_1934),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_1958),
.A2(n_1201),
.B1(n_1202),
.B2(n_1196),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1935),
.B(n_1205),
.Y(n_2247)
);

NOR2xp67_ASAP7_75t_L g2248 ( 
.A(n_1935),
.B(n_3),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1935),
.Y(n_2249)
);

INVx2_ASAP7_75t_SL g2250 ( 
.A(n_1945),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_1937),
.B(n_1207),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1945),
.B(n_1208),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1947),
.B(n_1212),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1938),
.B(n_1216),
.Y(n_2254)
);

INVx4_ASAP7_75t_L g2255 ( 
.A(n_1918),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1939),
.B(n_1232),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1950),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1936),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1941),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_1949),
.B(n_1250),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_1951),
.B(n_1251),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1952),
.Y(n_2262)
);

HB1xp67_ASAP7_75t_L g2263 ( 
.A(n_1783),
.Y(n_2263)
);

AOI22xp33_ASAP7_75t_L g2264 ( 
.A1(n_1825),
.A2(n_1341),
.B1(n_1388),
.B2(n_1337),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1843),
.B(n_1259),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_1783),
.B(n_1266),
.Y(n_2266)
);

NAND3xp33_ASAP7_75t_L g2267 ( 
.A(n_1845),
.B(n_1271),
.C(n_1268),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1843),
.B(n_1279),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_1843),
.B(n_1281),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1843),
.B(n_1285),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1959),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1843),
.B(n_1291),
.Y(n_2272)
);

NAND2x1_ASAP7_75t_L g2273 ( 
.A(n_1825),
.B(n_1337),
.Y(n_2273)
);

NOR2xp33_ASAP7_75t_L g2274 ( 
.A(n_1990),
.B(n_1293),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1805),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1843),
.B(n_1297),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1843),
.B(n_1308),
.Y(n_2277)
);

INVxp67_ASAP7_75t_SL g2278 ( 
.A(n_1990),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_SL g2279 ( 
.A(n_1809),
.B(n_1315),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1843),
.B(n_1318),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1805),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_1809),
.B(n_1321),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1843),
.B(n_1323),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_1805),
.Y(n_2284)
);

NOR2xp33_ASAP7_75t_L g2285 ( 
.A(n_1990),
.B(n_1324),
.Y(n_2285)
);

NOR2xp67_ASAP7_75t_L g2286 ( 
.A(n_1831),
.B(n_4),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1843),
.B(n_1334),
.Y(n_2287)
);

OAI21xp33_ASAP7_75t_L g2288 ( 
.A1(n_1734),
.A2(n_1398),
.B(n_1397),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1805),
.Y(n_2289)
);

AO22x2_ASAP7_75t_L g2290 ( 
.A1(n_1958),
.A2(n_1050),
.B1(n_1059),
.B2(n_1053),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_1809),
.B(n_1335),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1843),
.B(n_1336),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1805),
.Y(n_2293)
);

INVx4_ASAP7_75t_L g2294 ( 
.A(n_1762),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_1825),
.A2(n_1388),
.B1(n_1341),
.B2(n_1090),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_1809),
.B(n_1339),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_1990),
.B(n_1343),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_SL g2298 ( 
.A(n_1809),
.B(n_1349),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_1843),
.B(n_1357),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1805),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1805),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1843),
.B(n_1365),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_1843),
.B(n_1373),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_1990),
.B(n_1396),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_1809),
.B(n_1415),
.Y(n_2305)
);

AOI22xp33_ASAP7_75t_L g2306 ( 
.A1(n_1825),
.A2(n_1388),
.B1(n_1341),
.B2(n_1119),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_L g2307 ( 
.A1(n_2227),
.A2(n_1145),
.B(n_1103),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2278),
.B(n_1364),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_2104),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2049),
.B(n_1369),
.Y(n_2310)
);

AOI21xp5_ASAP7_75t_L g2311 ( 
.A1(n_2215),
.A2(n_1177),
.B(n_1162),
.Y(n_2311)
);

OAI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_2084),
.A2(n_1193),
.B1(n_1204),
.B2(n_1180),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2081),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1994),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2082),
.B(n_1404),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_1998),
.Y(n_2316)
);

AOI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2126),
.A2(n_1227),
.B1(n_1228),
.B2(n_1215),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2230),
.A2(n_1239),
.B(n_1235),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2022),
.B(n_1344),
.Y(n_2319)
);

NOR2xp67_ASAP7_75t_L g2320 ( 
.A(n_2294),
.B(n_2263),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2029),
.B(n_1347),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2036),
.B(n_1354),
.Y(n_2322)
);

BUFx8_ASAP7_75t_L g2323 ( 
.A(n_2037),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2038),
.Y(n_2324)
);

O2A1O1Ixp33_ASAP7_75t_L g2325 ( 
.A1(n_2143),
.A2(n_1244),
.B(n_1247),
.C(n_1242),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2039),
.B(n_1384),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2245),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_2203),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2041),
.Y(n_2329)
);

AOI21x1_ASAP7_75t_L g2330 ( 
.A1(n_2151),
.A2(n_1061),
.B(n_1024),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_2158),
.B(n_1393),
.Y(n_2331)
);

AOI21xp5_ASAP7_75t_L g2332 ( 
.A1(n_2152),
.A2(n_1256),
.B(n_1248),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2051),
.B(n_1405),
.Y(n_2333)
);

BUFx4f_ASAP7_75t_L g2334 ( 
.A(n_2144),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2065),
.B(n_1412),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2011),
.B(n_1416),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2073),
.B(n_1262),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2146),
.A2(n_1277),
.B(n_1276),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2106),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_2030),
.B(n_955),
.Y(n_2340)
);

OAI22xp5_ASAP7_75t_L g2341 ( 
.A1(n_2147),
.A2(n_1290),
.B1(n_1306),
.B2(n_1287),
.Y(n_2341)
);

O2A1O1Ixp33_ASAP7_75t_L g2342 ( 
.A1(n_2233),
.A2(n_1312),
.B(n_1328),
.C(n_1309),
.Y(n_2342)
);

AOI21x1_ASAP7_75t_L g2343 ( 
.A1(n_2248),
.A2(n_1078),
.B(n_1061),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2074),
.B(n_1375),
.Y(n_2344)
);

AO21x1_ASAP7_75t_L g2345 ( 
.A1(n_2211),
.A2(n_1331),
.B(n_1329),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2102),
.B(n_955),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2275),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2297),
.B(n_1401),
.Y(n_2348)
);

A2O1A1Ixp33_ASAP7_75t_L g2349 ( 
.A1(n_2129),
.A2(n_1361),
.B(n_1376),
.C(n_1333),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2190),
.B(n_1078),
.Y(n_2350)
);

AOI21xp5_ASAP7_75t_L g2351 ( 
.A1(n_2088),
.A2(n_1147),
.B(n_1094),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2281),
.B(n_1094),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2284),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_SL g2354 ( 
.A(n_2003),
.B(n_2053),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2289),
.B(n_1147),
.Y(n_2355)
);

AOI21xp5_ASAP7_75t_L g2356 ( 
.A1(n_2085),
.A2(n_1220),
.B(n_1199),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2293),
.Y(n_2357)
);

NOR2xp67_ASAP7_75t_L g2358 ( 
.A(n_2115),
.B(n_2),
.Y(n_2358)
);

AOI21xp5_ASAP7_75t_L g2359 ( 
.A1(n_2124),
.A2(n_1220),
.B(n_1199),
.Y(n_2359)
);

AOI22x1_ASAP7_75t_L g2360 ( 
.A1(n_2003),
.A2(n_1261),
.B1(n_961),
.B2(n_1185),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2300),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2301),
.B(n_1261),
.Y(n_2362)
);

INVxp67_ASAP7_75t_L g2363 ( 
.A(n_2019),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_2012),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2061),
.B(n_4),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2055),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2027),
.B(n_4),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2068),
.Y(n_2368)
);

NAND3xp33_ASAP7_75t_L g2369 ( 
.A(n_2209),
.B(n_1203),
.C(n_1185),
.Y(n_2369)
);

BUFx12f_ASAP7_75t_L g2370 ( 
.A(n_2145),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2031),
.B(n_5),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1999),
.B(n_5),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2005),
.B(n_1203),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2000),
.B(n_6),
.Y(n_2374)
);

BUFx4f_ASAP7_75t_L g2375 ( 
.A(n_2144),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2020),
.B(n_7),
.Y(n_2376)
);

INVx4_ASAP7_75t_L g2377 ( 
.A(n_2245),
.Y(n_2377)
);

AOI21xp5_ASAP7_75t_L g2378 ( 
.A1(n_2235),
.A2(n_1327),
.B(n_1203),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2060),
.Y(n_2379)
);

NAND2x1p5_ASAP7_75t_L g2380 ( 
.A(n_2025),
.B(n_1327),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2091),
.A2(n_1418),
.B(n_1327),
.Y(n_2381)
);

OAI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2023),
.A2(n_1418),
.B(n_7),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_2054),
.B(n_7),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2142),
.B(n_8),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2003),
.B(n_1418),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2093),
.A2(n_9),
.B(n_10),
.Y(n_2386)
);

INVxp67_ASAP7_75t_L g2387 ( 
.A(n_2266),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_L g2388 ( 
.A(n_2052),
.B(n_9),
.Y(n_2388)
);

HB1xp67_ASAP7_75t_L g2389 ( 
.A(n_2026),
.Y(n_2389)
);

BUFx6f_ASAP7_75t_L g2390 ( 
.A(n_2053),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2086),
.Y(n_2391)
);

AOI21xp5_ASAP7_75t_L g2392 ( 
.A1(n_2013),
.A2(n_10),
.B(n_11),
.Y(n_2392)
);

O2A1O1Ixp5_ASAP7_75t_L g2393 ( 
.A1(n_2006),
.A2(n_14),
.B(n_11),
.C(n_12),
.Y(n_2393)
);

AOI21xp5_ASAP7_75t_L g2394 ( 
.A1(n_2015),
.A2(n_11),
.B(n_12),
.Y(n_2394)
);

OAI321xp33_ASAP7_75t_L g2395 ( 
.A1(n_2127),
.A2(n_17),
.A3(n_19),
.B1(n_15),
.B2(n_16),
.C(n_18),
.Y(n_2395)
);

BUFx2_ASAP7_75t_L g2396 ( 
.A(n_2070),
.Y(n_2396)
);

O2A1O1Ixp33_ASAP7_75t_L g2397 ( 
.A1(n_1993),
.A2(n_1996),
.B(n_1997),
.C(n_2017),
.Y(n_2397)
);

AOI21xp33_ASAP7_75t_L g2398 ( 
.A1(n_2062),
.A2(n_15),
.B(n_16),
.Y(n_2398)
);

INVx3_ASAP7_75t_L g2399 ( 
.A(n_2242),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2053),
.B(n_19),
.Y(n_2400)
);

NAND2x1p5_ASAP7_75t_L g2401 ( 
.A(n_2025),
.B(n_17),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2007),
.B(n_20),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2095),
.B(n_20),
.Y(n_2403)
);

AOI21xp5_ASAP7_75t_L g2404 ( 
.A1(n_2032),
.A2(n_21),
.B(n_22),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2111),
.B(n_21),
.Y(n_2405)
);

AOI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2044),
.A2(n_22),
.B(n_23),
.Y(n_2406)
);

INVx3_ASAP7_75t_L g2407 ( 
.A(n_2242),
.Y(n_2407)
);

INVxp67_ASAP7_75t_L g2408 ( 
.A(n_2058),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2274),
.B(n_23),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2045),
.A2(n_24),
.B(n_25),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2137),
.A2(n_24),
.B(n_25),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2285),
.B(n_24),
.Y(n_2412)
);

NOR2xp33_ASAP7_75t_L g2413 ( 
.A(n_2205),
.B(n_26),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2304),
.B(n_26),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2128),
.A2(n_27),
.B(n_28),
.Y(n_2415)
);

INVx1_ASAP7_75t_SL g2416 ( 
.A(n_2185),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2010),
.B(n_28),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2063),
.Y(n_2418)
);

OAI21xp33_ASAP7_75t_L g2419 ( 
.A1(n_2160),
.A2(n_28),
.B(n_29),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2108),
.B(n_29),
.Y(n_2420)
);

OAI21xp33_ASAP7_75t_L g2421 ( 
.A1(n_2076),
.A2(n_30),
.B(n_31),
.Y(n_2421)
);

INVx3_ASAP7_75t_SL g2422 ( 
.A(n_2070),
.Y(n_2422)
);

AOI21xp5_ASAP7_75t_L g2423 ( 
.A1(n_2135),
.A2(n_30),
.B(n_31),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_2271),
.B(n_32),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2271),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2094),
.A2(n_31),
.B(n_32),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_L g2427 ( 
.A(n_2161),
.B(n_32),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2105),
.Y(n_2428)
);

AOI21xp5_ASAP7_75t_L g2429 ( 
.A1(n_2107),
.A2(n_33),
.B(n_34),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2170),
.B(n_33),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_2149),
.A2(n_34),
.B(n_35),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2047),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2154),
.A2(n_35),
.B(n_36),
.Y(n_2433)
);

AND2x2_ASAP7_75t_L g2434 ( 
.A(n_2002),
.B(n_37),
.Y(n_2434)
);

INVx3_ASAP7_75t_L g2435 ( 
.A(n_2242),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2101),
.B(n_38),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2148),
.B(n_40),
.Y(n_2437)
);

INVxp67_ASAP7_75t_L g2438 ( 
.A(n_2175),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2001),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2046),
.B(n_41),
.Y(n_2440)
);

OAI21xp5_ASAP7_75t_L g2441 ( 
.A1(n_2123),
.A2(n_42),
.B(n_43),
.Y(n_2441)
);

BUFx6f_ASAP7_75t_L g2442 ( 
.A(n_2271),
.Y(n_2442)
);

AND2x4_ASAP7_75t_L g2443 ( 
.A(n_2210),
.B(n_42),
.Y(n_2443)
);

INVx3_ASAP7_75t_L g2444 ( 
.A(n_2249),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_SL g2445 ( 
.A(n_2090),
.B(n_43),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2072),
.B(n_42),
.Y(n_2446)
);

AOI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2252),
.A2(n_44),
.B(n_45),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2177),
.B(n_2303),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2001),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_2449)
);

BUFx6f_ASAP7_75t_L g2450 ( 
.A(n_2249),
.Y(n_2450)
);

OAI21xp33_ASAP7_75t_L g2451 ( 
.A1(n_2153),
.A2(n_46),
.B(n_47),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2021),
.B(n_48),
.Y(n_2452)
);

INVx2_ASAP7_75t_SL g2453 ( 
.A(n_2040),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2004),
.B(n_48),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2121),
.B(n_47),
.Y(n_2455)
);

AOI21xp5_ASAP7_75t_L g2456 ( 
.A1(n_2067),
.A2(n_47),
.B(n_49),
.Y(n_2456)
);

A2O1A1Ixp33_ASAP7_75t_L g2457 ( 
.A1(n_2286),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2265),
.B(n_50),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2114),
.A2(n_50),
.B(n_51),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2268),
.B(n_51),
.Y(n_2460)
);

INVx2_ASAP7_75t_SL g2461 ( 
.A(n_2103),
.Y(n_2461)
);

AOI21xp5_ASAP7_75t_L g2462 ( 
.A1(n_2116),
.A2(n_52),
.B(n_53),
.Y(n_2462)
);

OAI22xp5_ASAP7_75t_L g2463 ( 
.A1(n_2096),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2463)
);

NOR2xp33_ASAP7_75t_L g2464 ( 
.A(n_2064),
.B(n_52),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2133),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_2249),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2162),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2269),
.B(n_54),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2270),
.B(n_2302),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2272),
.B(n_55),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2100),
.Y(n_2471)
);

AOI21xp5_ASAP7_75t_L g2472 ( 
.A1(n_2220),
.A2(n_55),
.B(n_56),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2165),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2109),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2121),
.B(n_55),
.Y(n_2475)
);

AOI21xp5_ASAP7_75t_L g2476 ( 
.A1(n_2254),
.A2(n_56),
.B(n_57),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2136),
.Y(n_2477)
);

BUFx4f_ASAP7_75t_L g2478 ( 
.A(n_2150),
.Y(n_2478)
);

AOI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2009),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2479)
);

INVx2_ASAP7_75t_SL g2480 ( 
.A(n_2181),
.Y(n_2480)
);

BUFx8_ASAP7_75t_SL g2481 ( 
.A(n_2037),
.Y(n_2481)
);

O2A1O1Ixp5_ASAP7_75t_L g2482 ( 
.A1(n_2273),
.A2(n_60),
.B(n_57),
.C(n_59),
.Y(n_2482)
);

AOI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2256),
.A2(n_59),
.B(n_60),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2276),
.B(n_60),
.Y(n_2484)
);

A2O1A1Ixp33_ASAP7_75t_L g2485 ( 
.A1(n_2286),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_2485)
);

AOI21xp5_ASAP7_75t_L g2486 ( 
.A1(n_2250),
.A2(n_61),
.B(n_62),
.Y(n_2486)
);

AND2x2_ASAP7_75t_L g2487 ( 
.A(n_2033),
.B(n_62),
.Y(n_2487)
);

NOR2xp33_ASAP7_75t_L g2488 ( 
.A(n_2191),
.B(n_63),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2290),
.B(n_64),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_SL g2490 ( 
.A(n_2034),
.B(n_2043),
.Y(n_2490)
);

OAI22xp5_ASAP7_75t_L g2491 ( 
.A1(n_2110),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2491)
);

AOI22xp5_ASAP7_75t_L g2492 ( 
.A1(n_2216),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2492)
);

BUFx12f_ASAP7_75t_L g2493 ( 
.A(n_2125),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2277),
.B(n_67),
.Y(n_2494)
);

OAI21xp5_ASAP7_75t_L g2495 ( 
.A1(n_2119),
.A2(n_67),
.B(n_68),
.Y(n_2495)
);

AOI21x1_ASAP7_75t_L g2496 ( 
.A1(n_2248),
.A2(n_67),
.B(n_68),
.Y(n_2496)
);

AOI21xp5_ASAP7_75t_L g2497 ( 
.A1(n_2219),
.A2(n_68),
.B(n_69),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2171),
.Y(n_2498)
);

AOI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_2008),
.A2(n_69),
.B(n_70),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_2024),
.B(n_69),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_L g2501 ( 
.A(n_1995),
.B(n_71),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2290),
.B(n_71),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2280),
.B(n_71),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2172),
.Y(n_2504)
);

NAND2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2210),
.B(n_72),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2194),
.Y(n_2506)
);

OAI321xp33_ASAP7_75t_L g2507 ( 
.A1(n_2089),
.A2(n_75),
.A3(n_77),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_2507)
);

AOI21xp5_ASAP7_75t_L g2508 ( 
.A1(n_2016),
.A2(n_73),
.B(n_74),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2283),
.B(n_73),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_2056),
.B(n_75),
.Y(n_2510)
);

OAI22xp5_ASAP7_75t_L g2511 ( 
.A1(n_2112),
.A2(n_2120),
.B1(n_2118),
.B2(n_2287),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2117),
.B(n_74),
.Y(n_2512)
);

O2A1O1Ixp33_ASAP7_75t_L g2513 ( 
.A1(n_2292),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2173),
.Y(n_2514)
);

AND2x2_ASAP7_75t_SL g2515 ( 
.A(n_2134),
.B(n_76),
.Y(n_2515)
);

AOI21xp5_ASAP7_75t_L g2516 ( 
.A1(n_2018),
.A2(n_78),
.B(n_79),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2299),
.B(n_78),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2157),
.Y(n_2518)
);

NOR2xp33_ASAP7_75t_L g2519 ( 
.A(n_2184),
.B(n_78),
.Y(n_2519)
);

AOI21xp5_ASAP7_75t_L g2520 ( 
.A1(n_2028),
.A2(n_79),
.B(n_80),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2182),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2138),
.B(n_79),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2122),
.B(n_80),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2216),
.B(n_2042),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2206),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2119),
.B(n_81),
.Y(n_2526)
);

AOI33xp33_ASAP7_75t_L g2527 ( 
.A1(n_2139),
.A2(n_83),
.A3(n_85),
.B1(n_81),
.B2(n_82),
.B3(n_84),
.Y(n_2527)
);

BUFx2_ASAP7_75t_L g2528 ( 
.A(n_2201),
.Y(n_2528)
);

AOI21x1_ASAP7_75t_L g2529 ( 
.A1(n_2206),
.A2(n_83),
.B(n_84),
.Y(n_2529)
);

NOR2xp33_ASAP7_75t_L g2530 ( 
.A(n_2071),
.B(n_83),
.Y(n_2530)
);

AOI21xp5_ASAP7_75t_L g2531 ( 
.A1(n_2192),
.A2(n_84),
.B(n_85),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2167),
.Y(n_2532)
);

AOI33xp33_ASAP7_75t_L g2533 ( 
.A1(n_2139),
.A2(n_2218),
.A3(n_2164),
.B1(n_2155),
.B2(n_2246),
.B3(n_2174),
.Y(n_2533)
);

NOR2xp33_ASAP7_75t_L g2534 ( 
.A(n_2159),
.B(n_85),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2202),
.B(n_2200),
.Y(n_2535)
);

AOI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2193),
.A2(n_86),
.B(n_87),
.Y(n_2536)
);

OAI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2069),
.A2(n_89),
.B1(n_86),
.B2(n_87),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_L g2538 ( 
.A(n_2092),
.B(n_86),
.Y(n_2538)
);

AOI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2050),
.A2(n_91),
.B1(n_87),
.B2(n_90),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2066),
.B(n_91),
.Y(n_2540)
);

AOI21xp5_ASAP7_75t_L g2541 ( 
.A1(n_2196),
.A2(n_90),
.B(n_91),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2176),
.Y(n_2542)
);

A2O1A1Ixp33_ASAP7_75t_L g2543 ( 
.A1(n_2288),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_2543)
);

OR2x2_ASAP7_75t_L g2544 ( 
.A(n_2156),
.B(n_92),
.Y(n_2544)
);

BUFx2_ASAP7_75t_L g2545 ( 
.A(n_2059),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2199),
.B(n_92),
.Y(n_2546)
);

AOI22xp5_ASAP7_75t_L g2547 ( 
.A1(n_2057),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_2547)
);

AOI22xp5_ASAP7_75t_L g2548 ( 
.A1(n_2087),
.A2(n_96),
.B1(n_93),
.B2(n_95),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_R g2549 ( 
.A(n_2197),
.B(n_96),
.Y(n_2549)
);

INVx2_ASAP7_75t_L g2550 ( 
.A(n_2208),
.Y(n_2550)
);

AOI21xp5_ASAP7_75t_L g2551 ( 
.A1(n_2189),
.A2(n_97),
.B(n_98),
.Y(n_2551)
);

INVxp67_ASAP7_75t_L g2552 ( 
.A(n_2166),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2228),
.B(n_97),
.Y(n_2553)
);

NOR3xp33_ASAP7_75t_L g2554 ( 
.A(n_2244),
.B(n_99),
.C(n_98),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2099),
.B(n_97),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2207),
.Y(n_2556)
);

OAI22xp5_ASAP7_75t_L g2557 ( 
.A1(n_2267),
.A2(n_100),
.B1(n_98),
.B2(n_99),
.Y(n_2557)
);

AOI21xp5_ASAP7_75t_L g2558 ( 
.A1(n_2238),
.A2(n_100),
.B(n_101),
.Y(n_2558)
);

AOI21xp5_ASAP7_75t_L g2559 ( 
.A1(n_2204),
.A2(n_101),
.B(n_102),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_2279),
.B(n_102),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_L g2561 ( 
.A(n_2282),
.B(n_102),
.Y(n_2561)
);

BUFx8_ASAP7_75t_L g2562 ( 
.A(n_2243),
.Y(n_2562)
);

HB1xp67_ASAP7_75t_L g2563 ( 
.A(n_2232),
.Y(n_2563)
);

AOI21xp5_ASAP7_75t_L g2564 ( 
.A1(n_2257),
.A2(n_103),
.B(n_104),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2188),
.B(n_105),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2237),
.Y(n_2566)
);

AOI21xp5_ASAP7_75t_L g2567 ( 
.A1(n_2187),
.A2(n_105),
.B(n_106),
.Y(n_2567)
);

AOI21x1_ASAP7_75t_L g2568 ( 
.A1(n_2083),
.A2(n_105),
.B(n_106),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_2198),
.B(n_2097),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2262),
.A2(n_106),
.B(n_107),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2078),
.B(n_2291),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_2098),
.B(n_107),
.Y(n_2572)
);

OAI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2150),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2296),
.B(n_108),
.Y(n_2574)
);

AOI21xp5_ASAP7_75t_L g2575 ( 
.A1(n_2258),
.A2(n_109),
.B(n_110),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2113),
.B(n_109),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2298),
.B(n_111),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_2150),
.Y(n_2578)
);

AOI21xp5_ASAP7_75t_L g2579 ( 
.A1(n_2259),
.A2(n_111),
.B(n_112),
.Y(n_2579)
);

A2O1A1Ixp33_ASAP7_75t_L g2580 ( 
.A1(n_2295),
.A2(n_2306),
.B(n_2264),
.C(n_2261),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2239),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_SL g2582 ( 
.A(n_2213),
.B(n_113),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2180),
.A2(n_112),
.B(n_114),
.Y(n_2583)
);

NOR2xp33_ASAP7_75t_L g2584 ( 
.A(n_2305),
.B(n_114),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2224),
.Y(n_2585)
);

O2A1O1Ixp33_ASAP7_75t_L g2586 ( 
.A1(n_2183),
.A2(n_118),
.B(n_116),
.C(n_117),
.Y(n_2586)
);

AOI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2214),
.A2(n_116),
.B(n_117),
.Y(n_2587)
);

OAI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_2195),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_2588)
);

AOI21xp5_ASAP7_75t_L g2589 ( 
.A1(n_2217),
.A2(n_119),
.B(n_120),
.Y(n_2589)
);

AO21x1_ASAP7_75t_L g2590 ( 
.A1(n_2255),
.A2(n_626),
.B(n_624),
.Y(n_2590)
);

AOI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2251),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_2591)
);

AND2x2_ASAP7_75t_L g2592 ( 
.A(n_2221),
.B(n_122),
.Y(n_2592)
);

NOR2x1_ASAP7_75t_L g2593 ( 
.A(n_2140),
.B(n_122),
.Y(n_2593)
);

BUFx12f_ASAP7_75t_L g2594 ( 
.A(n_2178),
.Y(n_2594)
);

AOI21xp5_ASAP7_75t_L g2595 ( 
.A1(n_2253),
.A2(n_123),
.B(n_124),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2212),
.A2(n_124),
.B(n_125),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2226),
.A2(n_124),
.B(n_125),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2222),
.B(n_125),
.Y(n_2598)
);

AO21x2_ASAP7_75t_L g2599 ( 
.A1(n_2168),
.A2(n_126),
.B(n_127),
.Y(n_2599)
);

OAI22x1_ASAP7_75t_L g2600 ( 
.A1(n_2141),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_2600)
);

BUFx8_ASAP7_75t_L g2601 ( 
.A(n_2223),
.Y(n_2601)
);

BUFx8_ASAP7_75t_SL g2602 ( 
.A(n_2231),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2186),
.B(n_126),
.Y(n_2603)
);

NAND2xp33_ASAP7_75t_SL g2604 ( 
.A(n_2169),
.B(n_128),
.Y(n_2604)
);

INVx4_ASAP7_75t_L g2605 ( 
.A(n_2178),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2179),
.B(n_130),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2226),
.A2(n_129),
.B(n_131),
.Y(n_2607)
);

OR2x2_ASAP7_75t_L g2608 ( 
.A(n_2234),
.B(n_129),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2236),
.B(n_129),
.Y(n_2609)
);

AOI21xp5_ASAP7_75t_L g2610 ( 
.A1(n_2229),
.A2(n_131),
.B(n_132),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2229),
.A2(n_131),
.B(n_132),
.Y(n_2611)
);

A2O1A1Ixp33_ASAP7_75t_L g2612 ( 
.A1(n_2260),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2612)
);

INVx2_ASAP7_75t_SL g2613 ( 
.A(n_2075),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2240),
.B(n_134),
.Y(n_2614)
);

BUFx6f_ASAP7_75t_L g2615 ( 
.A(n_2178),
.Y(n_2615)
);

OAI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_2131),
.A2(n_133),
.B(n_135),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2225),
.B(n_135),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_SL g2618 ( 
.A(n_2241),
.B(n_137),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2255),
.Y(n_2619)
);

CKINVDCx8_ASAP7_75t_R g2620 ( 
.A(n_2178),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2077),
.B(n_136),
.Y(n_2621)
);

INVx2_ASAP7_75t_SL g2622 ( 
.A(n_2080),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2048),
.B(n_2130),
.Y(n_2623)
);

INVx4_ASAP7_75t_L g2624 ( 
.A(n_2048),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_SL g2625 ( 
.A(n_2247),
.B(n_139),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2130),
.Y(n_2626)
);

AOI21xp5_ASAP7_75t_L g2627 ( 
.A1(n_2163),
.A2(n_138),
.B(n_139),
.Y(n_2627)
);

BUFx6f_ASAP7_75t_L g2628 ( 
.A(n_2163),
.Y(n_2628)
);

INVx3_ASAP7_75t_L g2629 ( 
.A(n_2132),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2081),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2081),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2278),
.B(n_138),
.Y(n_2632)
);

BUFx12f_ASAP7_75t_L g2633 ( 
.A(n_2145),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2278),
.B(n_141),
.Y(n_2634)
);

INVx5_ASAP7_75t_L g2635 ( 
.A(n_2294),
.Y(n_2635)
);

AOI21xp33_ASAP7_75t_L g2636 ( 
.A1(n_2158),
.A2(n_141),
.B(n_142),
.Y(n_2636)
);

OAI22xp5_ASAP7_75t_L g2637 ( 
.A1(n_2084),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2203),
.Y(n_2638)
);

AOI21xp5_ASAP7_75t_L g2639 ( 
.A1(n_2227),
.A2(n_142),
.B(n_144),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2294),
.Y(n_2640)
);

AOI21xp5_ASAP7_75t_L g2641 ( 
.A1(n_2227),
.A2(n_144),
.B(n_145),
.Y(n_2641)
);

NOR2xp33_ASAP7_75t_L g2642 ( 
.A(n_2158),
.B(n_145),
.Y(n_2642)
);

AOI21x1_ASAP7_75t_L g2643 ( 
.A1(n_2203),
.A2(n_146),
.B(n_147),
.Y(n_2643)
);

NOR2xp33_ASAP7_75t_L g2644 ( 
.A(n_2158),
.B(n_146),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2278),
.B(n_146),
.Y(n_2645)
);

AOI21xp5_ASAP7_75t_L g2646 ( 
.A1(n_2227),
.A2(n_148),
.B(n_149),
.Y(n_2646)
);

AOI21xp5_ASAP7_75t_L g2647 ( 
.A1(n_2227),
.A2(n_148),
.B(n_149),
.Y(n_2647)
);

AOI21xp5_ASAP7_75t_L g2648 ( 
.A1(n_2227),
.A2(n_148),
.B(n_150),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2084),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_2649)
);

BUFx2_ASAP7_75t_L g2650 ( 
.A(n_2263),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2081),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_SL g2652 ( 
.A(n_2003),
.B(n_151),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2081),
.Y(n_2653)
);

AOI21xp5_ASAP7_75t_L g2654 ( 
.A1(n_2227),
.A2(n_151),
.B(n_152),
.Y(n_2654)
);

OAI21xp5_ASAP7_75t_L g2655 ( 
.A1(n_2035),
.A2(n_152),
.B(n_153),
.Y(n_2655)
);

NAND2xp5_ASAP7_75t_L g2656 ( 
.A(n_2278),
.B(n_153),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2278),
.B(n_153),
.Y(n_2657)
);

O2A1O1Ixp33_ASAP7_75t_L g2658 ( 
.A1(n_2143),
.A2(n_156),
.B(n_154),
.C(n_155),
.Y(n_2658)
);

OR2x2_ASAP7_75t_L g2659 ( 
.A(n_2263),
.B(n_154),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2278),
.B(n_155),
.Y(n_2660)
);

AOI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2079),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_2661)
);

AOI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2227),
.A2(n_156),
.B(n_157),
.Y(n_2662)
);

AND2x4_ASAP7_75t_SL g2663 ( 
.A(n_2294),
.B(n_158),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2278),
.B(n_159),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2203),
.Y(n_2665)
);

AOI21xp5_ASAP7_75t_L g2666 ( 
.A1(n_2227),
.A2(n_159),
.B(n_160),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2158),
.B(n_161),
.Y(n_2667)
);

AOI21xp5_ASAP7_75t_L g2668 ( 
.A1(n_2227),
.A2(n_162),
.B(n_163),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2158),
.B(n_162),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2003),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_SL g2671 ( 
.A(n_2014),
.B(n_164),
.Y(n_2671)
);

BUFx2_ASAP7_75t_L g2672 ( 
.A(n_2263),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2014),
.B(n_164),
.Y(n_2673)
);

AOI21x1_ASAP7_75t_L g2674 ( 
.A1(n_2203),
.A2(n_163),
.B(n_164),
.Y(n_2674)
);

INVx3_ASAP7_75t_L g2675 ( 
.A(n_2245),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2081),
.Y(n_2676)
);

O2A1O1Ixp5_ASAP7_75t_L g2677 ( 
.A1(n_2006),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2278),
.B(n_165),
.Y(n_2678)
);

AOI21xp5_ASAP7_75t_L g2679 ( 
.A1(n_2227),
.A2(n_166),
.B(n_167),
.Y(n_2679)
);

INVx4_ASAP7_75t_L g2680 ( 
.A(n_2294),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2049),
.B(n_168),
.Y(n_2681)
);

AO21x1_ASAP7_75t_L g2682 ( 
.A1(n_2227),
.A2(n_627),
.B(n_626),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2081),
.Y(n_2683)
);

AOI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2227),
.A2(n_168),
.B(n_169),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2278),
.B(n_169),
.Y(n_2685)
);

NOR2xp33_ASAP7_75t_R g2686 ( 
.A(n_2104),
.B(n_169),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_2014),
.B(n_170),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2203),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2278),
.B(n_171),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2278),
.B(n_172),
.Y(n_2690)
);

AOI21xp5_ASAP7_75t_L g2691 ( 
.A1(n_2227),
.A2(n_172),
.B(n_173),
.Y(n_2691)
);

OAI21xp5_ASAP7_75t_L g2692 ( 
.A1(n_2035),
.A2(n_172),
.B(n_173),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2278),
.B(n_173),
.Y(n_2693)
);

NOR2xp33_ASAP7_75t_L g2694 ( 
.A(n_2158),
.B(n_174),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_SL g2695 ( 
.A(n_2003),
.B(n_174),
.Y(n_2695)
);

AOI21xp5_ASAP7_75t_L g2696 ( 
.A1(n_2227),
.A2(n_174),
.B(n_175),
.Y(n_2696)
);

BUFx4f_ASAP7_75t_L g2697 ( 
.A(n_2144),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2158),
.B(n_175),
.Y(n_2698)
);

OAI21xp5_ASAP7_75t_L g2699 ( 
.A1(n_2035),
.A2(n_175),
.B(n_176),
.Y(n_2699)
);

AOI21xp5_ASAP7_75t_L g2700 ( 
.A1(n_2227),
.A2(n_176),
.B(n_177),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2278),
.B(n_176),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2263),
.Y(n_2702)
);

AO21x2_ASAP7_75t_L g2703 ( 
.A1(n_2227),
.A2(n_177),
.B(n_178),
.Y(n_2703)
);

AOI21xp5_ASAP7_75t_L g2704 ( 
.A1(n_2227),
.A2(n_177),
.B(n_178),
.Y(n_2704)
);

AOI21xp5_ASAP7_75t_L g2705 ( 
.A1(n_2227),
.A2(n_179),
.B(n_180),
.Y(n_2705)
);

BUFx3_ASAP7_75t_L g2706 ( 
.A(n_2012),
.Y(n_2706)
);

OAI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2084),
.A2(n_181),
.B1(n_179),
.B2(n_180),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_2003),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2278),
.B(n_180),
.Y(n_2709)
);

O2A1O1Ixp33_ASAP7_75t_L g2710 ( 
.A1(n_2143),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2278),
.B(n_182),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2081),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2294),
.B(n_182),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2278),
.B(n_183),
.Y(n_2714)
);

AOI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2227),
.A2(n_183),
.B(n_184),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2278),
.B(n_184),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2278),
.B(n_184),
.Y(n_2717)
);

BUFx12f_ASAP7_75t_L g2718 ( 
.A(n_2145),
.Y(n_2718)
);

O2A1O1Ixp33_ASAP7_75t_L g2719 ( 
.A1(n_2143),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_2719)
);

AOI21xp5_ASAP7_75t_L g2720 ( 
.A1(n_2227),
.A2(n_185),
.B(n_186),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2081),
.Y(n_2721)
);

AOI21xp5_ASAP7_75t_L g2722 ( 
.A1(n_2227),
.A2(n_186),
.B(n_188),
.Y(n_2722)
);

OAI21xp5_ASAP7_75t_L g2723 ( 
.A1(n_2035),
.A2(n_189),
.B(n_190),
.Y(n_2723)
);

INVx4_ASAP7_75t_L g2724 ( 
.A(n_2294),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2278),
.B(n_189),
.Y(n_2725)
);

OAI321xp33_ASAP7_75t_L g2726 ( 
.A1(n_2144),
.A2(n_192),
.A3(n_194),
.B1(n_189),
.B2(n_191),
.C(n_193),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2081),
.Y(n_2727)
);

AOI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2227),
.A2(n_191),
.B(n_192),
.Y(n_2728)
);

INVx2_ASAP7_75t_SL g2729 ( 
.A(n_2294),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2049),
.B(n_191),
.Y(n_2730)
);

INVx2_ASAP7_75t_SL g2731 ( 
.A(n_2294),
.Y(n_2731)
);

OAI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2035),
.A2(n_192),
.B(n_193),
.Y(n_2732)
);

NOR2xp33_ASAP7_75t_L g2733 ( 
.A(n_2158),
.B(n_193),
.Y(n_2733)
);

NAND2xp33_ASAP7_75t_L g2734 ( 
.A(n_2003),
.B(n_195),
.Y(n_2734)
);

AOI21xp5_ASAP7_75t_L g2735 ( 
.A1(n_2227),
.A2(n_194),
.B(n_195),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2158),
.B(n_195),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2227),
.A2(n_196),
.B(n_197),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_SL g2738 ( 
.A(n_2014),
.B(n_197),
.Y(n_2738)
);

AOI21xp5_ASAP7_75t_L g2739 ( 
.A1(n_2227),
.A2(n_196),
.B(n_197),
.Y(n_2739)
);

AOI21xp5_ASAP7_75t_L g2740 ( 
.A1(n_2227),
.A2(n_196),
.B(n_198),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2081),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2278),
.B(n_199),
.Y(n_2742)
);

AOI21xp5_ASAP7_75t_L g2743 ( 
.A1(n_2227),
.A2(n_199),
.B(n_200),
.Y(n_2743)
);

AOI22xp5_ASAP7_75t_L g2744 ( 
.A1(n_2079),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_SL g2745 ( 
.A(n_2014),
.B(n_201),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2104),
.Y(n_2746)
);

AOI21xp5_ASAP7_75t_L g2747 ( 
.A1(n_2227),
.A2(n_200),
.B(n_201),
.Y(n_2747)
);

BUFx2_ASAP7_75t_L g2748 ( 
.A(n_2263),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_L g2749 ( 
.A(n_2158),
.B(n_202),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2278),
.B(n_202),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2003),
.Y(n_2751)
);

OR2x6_ASAP7_75t_L g2752 ( 
.A(n_2294),
.B(n_202),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2081),
.Y(n_2753)
);

OR2x2_ASAP7_75t_L g2754 ( 
.A(n_2263),
.B(n_203),
.Y(n_2754)
);

AOI21xp5_ASAP7_75t_L g2755 ( 
.A1(n_2227),
.A2(n_204),
.B(n_205),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2278),
.B(n_205),
.Y(n_2756)
);

AOI21xp5_ASAP7_75t_L g2757 ( 
.A1(n_2227),
.A2(n_205),
.B(n_206),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_L g2758 ( 
.A(n_2278),
.B(n_206),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2203),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2227),
.A2(n_207),
.B(n_208),
.Y(n_2760)
);

AOI21xp5_ASAP7_75t_L g2761 ( 
.A1(n_2227),
.A2(n_207),
.B(n_208),
.Y(n_2761)
);

AOI22xp33_ASAP7_75t_L g2762 ( 
.A1(n_2030),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2278),
.B(n_209),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2227),
.A2(n_210),
.B(n_211),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_2014),
.B(n_211),
.Y(n_2765)
);

AOI21xp5_ASAP7_75t_L g2766 ( 
.A1(n_2227),
.A2(n_210),
.B(n_211),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2081),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2049),
.B(n_210),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2014),
.B(n_213),
.Y(n_2769)
);

AOI21xp5_ASAP7_75t_L g2770 ( 
.A1(n_2227),
.A2(n_212),
.B(n_214),
.Y(n_2770)
);

AOI21xp5_ASAP7_75t_L g2771 ( 
.A1(n_2227),
.A2(n_214),
.B(n_215),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2003),
.Y(n_2772)
);

A2O1A1Ixp33_ASAP7_75t_L g2773 ( 
.A1(n_2146),
.A2(n_217),
.B(n_214),
.C(n_216),
.Y(n_2773)
);

AND2x4_ASAP7_75t_L g2774 ( 
.A(n_2294),
.B(n_216),
.Y(n_2774)
);

OAI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2084),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2245),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2158),
.B(n_217),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2030),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.Y(n_2778)
);

NAND2x1_ASAP7_75t_L g2779 ( 
.A(n_2003),
.B(n_218),
.Y(n_2779)
);

AOI21xp5_ASAP7_75t_L g2780 ( 
.A1(n_2227),
.A2(n_219),
.B(n_220),
.Y(n_2780)
);

AOI21xp5_ASAP7_75t_L g2781 ( 
.A1(n_2227),
.A2(n_220),
.B(n_221),
.Y(n_2781)
);

BUFx4f_ASAP7_75t_L g2782 ( 
.A(n_2144),
.Y(n_2782)
);

INVx1_ASAP7_75t_SL g2783 ( 
.A(n_2263),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2203),
.Y(n_2784)
);

OAI22xp5_ASAP7_75t_L g2785 ( 
.A1(n_2084),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2081),
.Y(n_2786)
);

OAI21xp33_ASAP7_75t_L g2787 ( 
.A1(n_2035),
.A2(n_222),
.B(n_223),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2278),
.B(n_222),
.Y(n_2788)
);

AOI22xp33_ASAP7_75t_L g2789 ( 
.A1(n_2030),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_2789)
);

NOR2xp33_ASAP7_75t_L g2790 ( 
.A(n_2158),
.B(n_224),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2227),
.A2(n_225),
.B(n_226),
.Y(n_2791)
);

NOR2xp33_ASAP7_75t_L g2792 ( 
.A(n_2158),
.B(n_227),
.Y(n_2792)
);

INVx4_ASAP7_75t_L g2793 ( 
.A(n_2294),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2203),
.Y(n_2794)
);

BUFx2_ASAP7_75t_L g2795 ( 
.A(n_2263),
.Y(n_2795)
);

O2A1O1Ixp33_ASAP7_75t_L g2796 ( 
.A1(n_2143),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2203),
.Y(n_2797)
);

HB1xp67_ASAP7_75t_L g2798 ( 
.A(n_2263),
.Y(n_2798)
);

AOI21xp5_ASAP7_75t_L g2799 ( 
.A1(n_2227),
.A2(n_230),
.B(n_231),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2227),
.A2(n_232),
.B(n_233),
.Y(n_2800)
);

BUFx4f_ASAP7_75t_SL g2801 ( 
.A(n_2294),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2294),
.B(n_232),
.Y(n_2802)
);

OAI22xp5_ASAP7_75t_L g2803 ( 
.A1(n_2084),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_2803)
);

O2A1O1Ixp33_ASAP7_75t_L g2804 ( 
.A1(n_2143),
.A2(n_237),
.B(n_235),
.C(n_236),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2278),
.B(n_235),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2278),
.B(n_236),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2081),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2081),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2003),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2203),
.Y(n_2810)
);

NOR2xp33_ASAP7_75t_L g2811 ( 
.A(n_2158),
.B(n_239),
.Y(n_2811)
);

AOI33xp33_ASAP7_75t_L g2812 ( 
.A1(n_2033),
.A2(n_241),
.A3(n_243),
.B1(n_239),
.B2(n_240),
.B3(n_242),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_2245),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2245),
.Y(n_2814)
);

OAI21xp33_ASAP7_75t_L g2815 ( 
.A1(n_2035),
.A2(n_244),
.B(n_246),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_SL g2816 ( 
.A(n_2014),
.B(n_248),
.Y(n_2816)
);

OAI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2035),
.A2(n_247),
.B(n_249),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2081),
.Y(n_2818)
);

CKINVDCx8_ASAP7_75t_R g2819 ( 
.A(n_2145),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2081),
.Y(n_2820)
);

NOR3xp33_ASAP7_75t_L g2821 ( 
.A(n_2079),
.B(n_250),
.C(n_249),
.Y(n_2821)
);

O2A1O1Ixp33_ASAP7_75t_L g2822 ( 
.A1(n_2143),
.A2(n_253),
.B(n_251),
.C(n_252),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2278),
.B(n_252),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2081),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2278),
.B(n_253),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_SL g2826 ( 
.A(n_2014),
.B(n_254),
.Y(n_2826)
);

INVxp67_ASAP7_75t_L g2827 ( 
.A(n_2263),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2203),
.Y(n_2828)
);

NAND2x1p5_ASAP7_75t_L g2829 ( 
.A(n_2294),
.B(n_255),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2278),
.B(n_257),
.Y(n_2830)
);

BUFx2_ASAP7_75t_L g2831 ( 
.A(n_2263),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_SL g2832 ( 
.A(n_2014),
.B(n_260),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2227),
.A2(n_258),
.B(n_260),
.Y(n_2833)
);

OAI21xp5_ASAP7_75t_L g2834 ( 
.A1(n_2035),
.A2(n_261),
.B(n_262),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2227),
.A2(n_261),
.B(n_262),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2294),
.B(n_262),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2227),
.A2(n_263),
.B(n_264),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2278),
.B(n_263),
.Y(n_2838)
);

OAI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_2752),
.A2(n_265),
.B1(n_263),
.B2(n_264),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2471),
.B(n_265),
.Y(n_2840)
);

AOI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2397),
.A2(n_265),
.B(n_266),
.Y(n_2841)
);

INVx2_ASAP7_75t_L g2842 ( 
.A(n_2329),
.Y(n_2842)
);

BUFx4f_ASAP7_75t_L g2843 ( 
.A(n_2752),
.Y(n_2843)
);

OR2x6_ASAP7_75t_L g2844 ( 
.A(n_2752),
.B(n_266),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_2481),
.Y(n_2845)
);

OA21x2_ASAP7_75t_L g2846 ( 
.A1(n_2328),
.A2(n_267),
.B(n_268),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_SL g2847 ( 
.A(n_2334),
.B(n_629),
.Y(n_2847)
);

NOR2xp67_ASAP7_75t_SL g2848 ( 
.A(n_2620),
.B(n_268),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2474),
.B(n_269),
.Y(n_2849)
);

INVx1_ASAP7_75t_SL g2850 ( 
.A(n_2783),
.Y(n_2850)
);

OAI22xp5_ASAP7_75t_L g2851 ( 
.A1(n_2511),
.A2(n_271),
.B1(n_269),
.B2(n_270),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2638),
.A2(n_270),
.B(n_271),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2821),
.B(n_270),
.Y(n_2853)
);

AND3x1_ASAP7_75t_SL g2854 ( 
.A(n_2686),
.B(n_272),
.C(n_273),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2361),
.Y(n_2855)
);

NOR2xp33_ASAP7_75t_L g2856 ( 
.A(n_2387),
.B(n_272),
.Y(n_2856)
);

OAI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2661),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2831),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2313),
.Y(n_2859)
);

INVx6_ASAP7_75t_L g2860 ( 
.A(n_2635),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2314),
.Y(n_2861)
);

O2A1O1Ixp33_ASAP7_75t_SL g2862 ( 
.A1(n_2773),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_2375),
.B(n_629),
.Y(n_2863)
);

AOI21xp5_ASAP7_75t_L g2864 ( 
.A1(n_2665),
.A2(n_275),
.B(n_276),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2533),
.B(n_276),
.Y(n_2865)
);

BUFx6f_ASAP7_75t_L g2866 ( 
.A(n_2390),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2316),
.B(n_2324),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_2801),
.Y(n_2868)
);

INVx3_ASAP7_75t_L g2869 ( 
.A(n_2377),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2650),
.Y(n_2870)
);

OR2x6_ASAP7_75t_L g2871 ( 
.A(n_2377),
.B(n_277),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2347),
.B(n_278),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2635),
.B(n_278),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2353),
.Y(n_2874)
);

NOR2xp33_ASAP7_75t_SL g2875 ( 
.A(n_2819),
.B(n_279),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2368),
.Y(n_2876)
);

BUFx2_ASAP7_75t_L g2877 ( 
.A(n_2672),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2375),
.B(n_630),
.Y(n_2878)
);

INVx4_ASAP7_75t_L g2879 ( 
.A(n_2635),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2357),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2630),
.B(n_280),
.Y(n_2881)
);

BUFx6f_ASAP7_75t_L g2882 ( 
.A(n_2390),
.Y(n_2882)
);

AND2x4_ASAP7_75t_L g2883 ( 
.A(n_2680),
.B(n_280),
.Y(n_2883)
);

BUFx3_ASAP7_75t_L g2884 ( 
.A(n_2364),
.Y(n_2884)
);

BUFx4_ASAP7_75t_SL g2885 ( 
.A(n_2309),
.Y(n_2885)
);

A2O1A1Ixp33_ASAP7_75t_SL g2886 ( 
.A1(n_2609),
.A2(n_2382),
.B(n_2692),
.C(n_2655),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2631),
.B(n_280),
.Y(n_2887)
);

AOI21xp5_ASAP7_75t_L g2888 ( 
.A1(n_2688),
.A2(n_281),
.B(n_282),
.Y(n_2888)
);

AND2x6_ASAP7_75t_L g2889 ( 
.A(n_2615),
.B(n_282),
.Y(n_2889)
);

INVx3_ASAP7_75t_L g2890 ( 
.A(n_2724),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2391),
.Y(n_2891)
);

BUFx6f_ASAP7_75t_L g2892 ( 
.A(n_2390),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2428),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2759),
.A2(n_283),
.B(n_284),
.Y(n_2894)
);

OAI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2661),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_2408),
.B(n_2524),
.Y(n_2896)
);

OAI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2535),
.A2(n_285),
.B(n_286),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2552),
.B(n_285),
.Y(n_2898)
);

NOR2xp67_ASAP7_75t_SL g2899 ( 
.A(n_2594),
.B(n_287),
.Y(n_2899)
);

OAI21xp33_ASAP7_75t_L g2900 ( 
.A1(n_2451),
.A2(n_2421),
.B(n_2419),
.Y(n_2900)
);

O2A1O1Ixp33_ASAP7_75t_SL g2901 ( 
.A1(n_2525),
.A2(n_290),
.B(n_287),
.C(n_288),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2651),
.Y(n_2902)
);

INVx2_ASAP7_75t_L g2903 ( 
.A(n_2653),
.Y(n_2903)
);

INVx2_ASAP7_75t_L g2904 ( 
.A(n_2676),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2683),
.B(n_288),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2712),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2721),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2727),
.B(n_290),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_SL g2909 ( 
.A(n_2697),
.B(n_2782),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2744),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_2910)
);

OAI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2744),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_2911)
);

BUFx6f_ASAP7_75t_L g2912 ( 
.A(n_2425),
.Y(n_2912)
);

A2O1A1Ixp33_ASAP7_75t_L g2913 ( 
.A1(n_2419),
.A2(n_295),
.B(n_292),
.C(n_294),
.Y(n_2913)
);

NOR2xp33_ASAP7_75t_L g2914 ( 
.A(n_2396),
.B(n_294),
.Y(n_2914)
);

A2O1A1Ixp33_ASAP7_75t_L g2915 ( 
.A1(n_2451),
.A2(n_296),
.B(n_294),
.C(n_295),
.Y(n_2915)
);

AO32x2_ASAP7_75t_L g2916 ( 
.A1(n_2449),
.A2(n_297),
.A3(n_295),
.B1(n_296),
.B2(n_298),
.Y(n_2916)
);

OAI22x1_ASAP7_75t_L g2917 ( 
.A1(n_2829),
.A2(n_2422),
.B1(n_2492),
.B2(n_2572),
.Y(n_2917)
);

NOR3xp33_ASAP7_75t_SL g2918 ( 
.A(n_2339),
.B(n_2746),
.C(n_2519),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2741),
.B(n_297),
.Y(n_2919)
);

BUFx2_ASAP7_75t_L g2920 ( 
.A(n_2702),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2697),
.B(n_630),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_SL g2922 ( 
.A(n_2782),
.B(n_631),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2753),
.B(n_298),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2515),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2767),
.B(n_300),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_SL g2926 ( 
.A(n_2652),
.B(n_632),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2786),
.B(n_300),
.Y(n_2927)
);

BUFx6f_ASAP7_75t_L g2928 ( 
.A(n_2425),
.Y(n_2928)
);

OAI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2479),
.A2(n_304),
.B1(n_302),
.B2(n_303),
.Y(n_2929)
);

AOI21xp5_ASAP7_75t_L g2930 ( 
.A1(n_2784),
.A2(n_302),
.B(n_303),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2489),
.B(n_302),
.Y(n_2931)
);

BUFx3_ASAP7_75t_L g2932 ( 
.A(n_2706),
.Y(n_2932)
);

AOI22xp33_ASAP7_75t_L g2933 ( 
.A1(n_2413),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_2933)
);

NAND3xp33_ASAP7_75t_L g2934 ( 
.A(n_2543),
.B(n_305),
.C(n_306),
.Y(n_2934)
);

AND2x2_ASAP7_75t_L g2935 ( 
.A(n_2502),
.B(n_307),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2807),
.Y(n_2936)
);

AOI21xp5_ASAP7_75t_L g2937 ( 
.A1(n_2794),
.A2(n_307),
.B(n_308),
.Y(n_2937)
);

OA22x2_ASAP7_75t_L g2938 ( 
.A1(n_2663),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_2938)
);

O2A1O1Ixp33_ASAP7_75t_L g2939 ( 
.A1(n_2522),
.A2(n_310),
.B(n_308),
.C(n_309),
.Y(n_2939)
);

AOI21xp5_ASAP7_75t_L g2940 ( 
.A1(n_2797),
.A2(n_310),
.B(n_311),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2810),
.A2(n_310),
.B(n_311),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_L g2942 ( 
.A(n_2363),
.B(n_311),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2808),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2818),
.Y(n_2944)
);

AO22x1_ASAP7_75t_L g2945 ( 
.A1(n_2323),
.A2(n_314),
.B1(n_312),
.B2(n_313),
.Y(n_2945)
);

AO32x1_ASAP7_75t_L g2946 ( 
.A1(n_2573),
.A2(n_2432),
.A3(n_2557),
.B1(n_2537),
.B2(n_2637),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_SL g2947 ( 
.A(n_2652),
.B(n_2695),
.Y(n_2947)
);

AND2x4_ASAP7_75t_L g2948 ( 
.A(n_2724),
.B(n_313),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_SL g2949 ( 
.A(n_2695),
.B(n_633),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2828),
.A2(n_314),
.B(n_315),
.Y(n_2950)
);

BUFx6f_ASAP7_75t_L g2951 ( 
.A(n_2425),
.Y(n_2951)
);

AOI21xp5_ASAP7_75t_L g2952 ( 
.A1(n_2469),
.A2(n_315),
.B(n_316),
.Y(n_2952)
);

O2A1O1Ixp33_ASAP7_75t_L g2953 ( 
.A1(n_2372),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_2953)
);

BUFx6f_ASAP7_75t_L g2954 ( 
.A(n_2442),
.Y(n_2954)
);

A2O1A1Ixp33_ASAP7_75t_SL g2955 ( 
.A1(n_2699),
.A2(n_319),
.B(n_317),
.C(n_318),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_SL g2956 ( 
.A(n_2793),
.B(n_317),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2354),
.A2(n_318),
.B(n_319),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_SL g2958 ( 
.A(n_2549),
.B(n_633),
.Y(n_2958)
);

NOR2xp67_ASAP7_75t_SL g2959 ( 
.A(n_2793),
.B(n_320),
.Y(n_2959)
);

INVx3_ASAP7_75t_L g2960 ( 
.A(n_2493),
.Y(n_2960)
);

O2A1O1Ixp33_ASAP7_75t_L g2961 ( 
.A1(n_2383),
.A2(n_2409),
.B(n_2414),
.C(n_2412),
.Y(n_2961)
);

AOI21xp5_ASAP7_75t_L g2962 ( 
.A1(n_2354),
.A2(n_320),
.B(n_321),
.Y(n_2962)
);

NOR2xp33_ASAP7_75t_L g2963 ( 
.A(n_2389),
.B(n_2571),
.Y(n_2963)
);

AOI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2315),
.A2(n_321),
.B(n_322),
.Y(n_2964)
);

HB1xp67_ASAP7_75t_L g2965 ( 
.A(n_2748),
.Y(n_2965)
);

O2A1O1Ixp33_ASAP7_75t_L g2966 ( 
.A1(n_2319),
.A2(n_325),
.B(n_323),
.C(n_324),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2827),
.B(n_323),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2820),
.B(n_324),
.Y(n_2968)
);

A2O1A1Ixp33_ASAP7_75t_L g2969 ( 
.A1(n_2421),
.A2(n_2472),
.B(n_2732),
.C(n_2723),
.Y(n_2969)
);

BUFx6f_ASAP7_75t_L g2970 ( 
.A(n_2442),
.Y(n_2970)
);

BUFx2_ASAP7_75t_L g2971 ( 
.A(n_2795),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2824),
.B(n_324),
.Y(n_2972)
);

INVx4_ASAP7_75t_L g2973 ( 
.A(n_2478),
.Y(n_2973)
);

CKINVDCx14_ASAP7_75t_R g2974 ( 
.A(n_2370),
.Y(n_2974)
);

AOI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2488),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_SL g2976 ( 
.A(n_2320),
.B(n_635),
.Y(n_2976)
);

AOI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_2448),
.A2(n_326),
.B(n_327),
.Y(n_2977)
);

OAI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2479),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_2978)
);

AOI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2580),
.A2(n_328),
.B(n_329),
.Y(n_2979)
);

INVxp67_ASAP7_75t_L g2980 ( 
.A(n_2798),
.Y(n_2980)
);

AOI22xp5_ASAP7_75t_L g2981 ( 
.A1(n_2443),
.A2(n_2534),
.B1(n_2644),
.B2(n_2642),
.Y(n_2981)
);

OAI21x1_ASAP7_75t_L g2982 ( 
.A1(n_2343),
.A2(n_330),
.B(n_331),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2465),
.Y(n_2983)
);

AOI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_2365),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2984)
);

NAND3xp33_ASAP7_75t_SL g2985 ( 
.A(n_2829),
.B(n_330),
.C(n_331),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2438),
.B(n_332),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2532),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2327),
.B(n_2675),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2542),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2556),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2436),
.Y(n_2991)
);

BUFx6f_ASAP7_75t_L g2992 ( 
.A(n_2442),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2366),
.Y(n_2993)
);

BUFx2_ASAP7_75t_L g2994 ( 
.A(n_2713),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_L g2995 ( 
.A(n_2348),
.B(n_333),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2443),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2681),
.B(n_336),
.Y(n_2997)
);

A2O1A1Ixp33_ASAP7_75t_L g2998 ( 
.A1(n_2817),
.A2(n_339),
.B(n_337),
.C(n_338),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2730),
.B(n_337),
.Y(n_2999)
);

O2A1O1Ixp33_ASAP7_75t_L g3000 ( 
.A1(n_2398),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_3000)
);

AOI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2667),
.A2(n_340),
.B1(n_338),
.B2(n_339),
.Y(n_3001)
);

BUFx2_ASAP7_75t_L g3002 ( 
.A(n_2713),
.Y(n_3002)
);

AOI22xp33_ASAP7_75t_L g3003 ( 
.A1(n_2669),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.Y(n_3003)
);

OAI21xp5_ASAP7_75t_L g3004 ( 
.A1(n_2349),
.A2(n_341),
.B(n_342),
.Y(n_3004)
);

AND2x4_ASAP7_75t_L g3005 ( 
.A(n_2327),
.B(n_341),
.Y(n_3005)
);

INVx3_ASAP7_75t_L g3006 ( 
.A(n_2675),
.Y(n_3006)
);

INVxp67_ASAP7_75t_L g3007 ( 
.A(n_2774),
.Y(n_3007)
);

A2O1A1Ixp33_ASAP7_75t_L g3008 ( 
.A1(n_2834),
.A2(n_346),
.B(n_344),
.C(n_345),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2539),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_3009)
);

AOI21x1_ASAP7_75t_L g3010 ( 
.A1(n_2330),
.A2(n_348),
.B(n_349),
.Y(n_3010)
);

INVx3_ASAP7_75t_L g3011 ( 
.A(n_2776),
.Y(n_3011)
);

BUFx3_ASAP7_75t_L g3012 ( 
.A(n_2323),
.Y(n_3012)
);

NAND2x1p5_ASAP7_75t_L g3013 ( 
.A(n_2478),
.B(n_348),
.Y(n_3013)
);

BUFx6f_ASAP7_75t_L g3014 ( 
.A(n_2670),
.Y(n_3014)
);

OAI21x1_ASAP7_75t_L g3015 ( 
.A1(n_2643),
.A2(n_349),
.B(n_350),
.Y(n_3015)
);

OAI22xp5_ASAP7_75t_L g3016 ( 
.A1(n_2539),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_SL g3017 ( 
.A(n_2450),
.B(n_2605),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2581),
.B(n_350),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2437),
.Y(n_3019)
);

OAI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2547),
.A2(n_354),
.B1(n_351),
.B2(n_352),
.Y(n_3020)
);

O2A1O1Ixp5_ASAP7_75t_L g3021 ( 
.A1(n_2345),
.A2(n_354),
.B(n_351),
.C(n_352),
.Y(n_3021)
);

O2A1O1Ixp33_ASAP7_75t_L g3022 ( 
.A1(n_2523),
.A2(n_2582),
.B(n_2538),
.C(n_2612),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2450),
.B(n_636),
.Y(n_3023)
);

BUFx4f_ASAP7_75t_L g3024 ( 
.A(n_2633),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_SL g3025 ( 
.A(n_2450),
.B(n_637),
.Y(n_3025)
);

HB1xp67_ASAP7_75t_L g3026 ( 
.A(n_2416),
.Y(n_3026)
);

O2A1O1Ixp5_ASAP7_75t_L g3027 ( 
.A1(n_2346),
.A2(n_357),
.B(n_355),
.C(n_356),
.Y(n_3027)
);

A2O1A1Ixp33_ASAP7_75t_L g3028 ( 
.A1(n_2392),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_3028)
);

CKINVDCx5p33_ASAP7_75t_R g3029 ( 
.A(n_2718),
.Y(n_3029)
);

AOI22xp5_ASAP7_75t_L g3030 ( 
.A1(n_2694),
.A2(n_2733),
.B1(n_2736),
.B2(n_2698),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2768),
.B(n_356),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2379),
.Y(n_3032)
);

AOI21xp5_ASAP7_75t_L g3033 ( 
.A1(n_2569),
.A2(n_358),
.B(n_359),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_L g3034 ( 
.A1(n_2749),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_3034)
);

NOR2x1_ASAP7_75t_SL g3035 ( 
.A(n_2605),
.B(n_359),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2418),
.Y(n_3036)
);

O2A1O1Ixp5_ASAP7_75t_L g3037 ( 
.A1(n_2373),
.A2(n_362),
.B(n_360),
.C(n_361),
.Y(n_3037)
);

OR2x6_ASAP7_75t_L g3038 ( 
.A(n_2774),
.B(n_361),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_SL g3039 ( 
.A(n_2416),
.B(n_638),
.Y(n_3039)
);

OAI21xp5_ASAP7_75t_L g3040 ( 
.A1(n_2317),
.A2(n_363),
.B(n_364),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_SL g3041 ( 
.A(n_2802),
.B(n_639),
.Y(n_3041)
);

A2O1A1Ixp33_ASAP7_75t_L g3042 ( 
.A1(n_2394),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_L g3043 ( 
.A(n_2566),
.B(n_2477),
.Y(n_3043)
);

AOI21xp5_ASAP7_75t_L g3044 ( 
.A1(n_2546),
.A2(n_365),
.B(n_366),
.Y(n_3044)
);

AO21x1_ASAP7_75t_L g3045 ( 
.A1(n_2505),
.A2(n_640),
.B(n_639),
.Y(n_3045)
);

BUFx8_ASAP7_75t_L g3046 ( 
.A(n_2802),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2405),
.B(n_367),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2467),
.Y(n_3048)
);

AOI21x1_ASAP7_75t_L g3049 ( 
.A1(n_2674),
.A2(n_367),
.B(n_368),
.Y(n_3049)
);

AND2x2_ASAP7_75t_L g3050 ( 
.A(n_2455),
.B(n_367),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2527),
.Y(n_3051)
);

CKINVDCx5p33_ASAP7_75t_R g3052 ( 
.A(n_2602),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2812),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2317),
.B(n_369),
.Y(n_3054)
);

BUFx2_ASAP7_75t_L g3055 ( 
.A(n_2836),
.Y(n_3055)
);

OA21x2_ASAP7_75t_L g3056 ( 
.A1(n_2369),
.A2(n_369),
.B(n_370),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2367),
.B(n_370),
.Y(n_3057)
);

AOI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2777),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2659),
.Y(n_3059)
);

NOR2xp33_ASAP7_75t_L g3060 ( 
.A(n_2518),
.B(n_371),
.Y(n_3060)
);

OR2x6_ASAP7_75t_SL g3061 ( 
.A(n_2754),
.B(n_372),
.Y(n_3061)
);

OAI22xp5_ASAP7_75t_L g3062 ( 
.A1(n_2548),
.A2(n_2591),
.B1(n_2634),
.B2(n_2632),
.Y(n_3062)
);

NAND3xp33_ASAP7_75t_SL g3063 ( 
.A(n_2554),
.B(n_373),
.C(n_374),
.Y(n_3063)
);

BUFx3_ASAP7_75t_L g3064 ( 
.A(n_2562),
.Y(n_3064)
);

CKINVDCx5p33_ASAP7_75t_R g3065 ( 
.A(n_2601),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2401),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_SL g3067 ( 
.A(n_2836),
.B(n_641),
.Y(n_3067)
);

NAND2x1p5_ASAP7_75t_L g3068 ( 
.A(n_2813),
.B(n_2814),
.Y(n_3068)
);

OAI22xp5_ASAP7_75t_L g3069 ( 
.A1(n_2548),
.A2(n_378),
.B1(n_375),
.B2(n_376),
.Y(n_3069)
);

A2O1A1Ixp33_ASAP7_75t_L g3070 ( 
.A1(n_2404),
.A2(n_380),
.B(n_376),
.C(n_379),
.Y(n_3070)
);

BUFx6f_ASAP7_75t_L g3071 ( 
.A(n_2670),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_2430),
.B(n_379),
.Y(n_3072)
);

NOR2xp33_ASAP7_75t_L g3073 ( 
.A(n_2790),
.B(n_381),
.Y(n_3073)
);

BUFx6f_ASAP7_75t_L g3074 ( 
.A(n_2670),
.Y(n_3074)
);

INVx5_ASAP7_75t_L g3075 ( 
.A(n_2708),
.Y(n_3075)
);

OAI21x1_ASAP7_75t_L g3076 ( 
.A1(n_2378),
.A2(n_381),
.B(n_382),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2371),
.B(n_384),
.Y(n_3077)
);

AO22x1_ASAP7_75t_L g3078 ( 
.A1(n_2495),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2473),
.Y(n_3079)
);

OAI22xp5_ASAP7_75t_L g3080 ( 
.A1(n_2591),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_3080)
);

AOI222xp33_ASAP7_75t_L g3081 ( 
.A1(n_2310),
.A2(n_387),
.B1(n_390),
.B2(n_385),
.C1(n_386),
.C2(n_388),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2458),
.A2(n_387),
.B(n_388),
.Y(n_3082)
);

AOI21x1_ASAP7_75t_L g3083 ( 
.A1(n_2496),
.A2(n_388),
.B(n_390),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2475),
.B(n_2553),
.Y(n_3084)
);

INVx3_ASAP7_75t_L g3085 ( 
.A(n_2813),
.Y(n_3085)
);

BUFx2_ASAP7_75t_SL g3086 ( 
.A(n_2814),
.Y(n_3086)
);

AO32x1_ASAP7_75t_L g3087 ( 
.A1(n_2649),
.A2(n_392),
.A3(n_390),
.B1(n_391),
.B2(n_393),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2708),
.B(n_642),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2487),
.B(n_2434),
.Y(n_3089)
);

OAI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2460),
.A2(n_2470),
.B(n_2468),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2645),
.A2(n_394),
.B1(n_391),
.B2(n_392),
.Y(n_3091)
);

OAI21xp5_ASAP7_75t_L g3092 ( 
.A1(n_2484),
.A2(n_391),
.B(n_394),
.Y(n_3092)
);

BUFx2_ASAP7_75t_L g3093 ( 
.A(n_2601),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_SL g3094 ( 
.A(n_2708),
.B(n_2751),
.Y(n_3094)
);

AOI221x1_ASAP7_75t_L g3095 ( 
.A1(n_2787),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.C(n_398),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2401),
.Y(n_3096)
);

AO21x1_ASAP7_75t_L g3097 ( 
.A1(n_2441),
.A2(n_644),
.B(n_643),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2656),
.A2(n_398),
.B1(n_396),
.B2(n_397),
.Y(n_3098)
);

AOI21xp5_ASAP7_75t_L g3099 ( 
.A1(n_2494),
.A2(n_397),
.B(n_398),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2384),
.B(n_2374),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2498),
.Y(n_3101)
);

BUFx3_ASAP7_75t_L g3102 ( 
.A(n_2562),
.Y(n_3102)
);

AND2x4_ASAP7_75t_L g3103 ( 
.A(n_2640),
.B(n_399),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2544),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2503),
.A2(n_399),
.B(n_400),
.Y(n_3105)
);

INVx3_ASAP7_75t_L g3106 ( 
.A(n_2729),
.Y(n_3106)
);

NAND2xp5_ASAP7_75t_L g3107 ( 
.A(n_2341),
.B(n_399),
.Y(n_3107)
);

AND2x4_ASAP7_75t_L g3108 ( 
.A(n_2731),
.B(n_400),
.Y(n_3108)
);

AOI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2509),
.A2(n_400),
.B(n_401),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2504),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2402),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2514),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2512),
.B(n_402),
.Y(n_3113)
);

BUFx2_ASAP7_75t_L g3114 ( 
.A(n_2528),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2517),
.A2(n_402),
.B(n_403),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2312),
.B(n_402),
.Y(n_3116)
);

NAND2x1p5_ASAP7_75t_L g3117 ( 
.A(n_2578),
.B(n_404),
.Y(n_3117)
);

A2O1A1Ixp33_ASAP7_75t_L g3118 ( 
.A1(n_2406),
.A2(n_406),
.B(n_404),
.C(n_405),
.Y(n_3118)
);

NOR3xp33_ASAP7_75t_SL g3119 ( 
.A(n_2726),
.B(n_406),
.C(n_407),
.Y(n_3119)
);

A2O1A1Ixp33_ASAP7_75t_L g3120 ( 
.A1(n_2410),
.A2(n_2787),
.B(n_2815),
.C(n_2513),
.Y(n_3120)
);

AOI22xp5_ASAP7_75t_L g3121 ( 
.A1(n_2792),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_3121)
);

OAI21xp5_ASAP7_75t_L g3122 ( 
.A1(n_2332),
.A2(n_408),
.B(n_409),
.Y(n_3122)
);

AOI22xp33_ASAP7_75t_L g3123 ( 
.A1(n_2811),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_2657),
.Y(n_3124)
);

AOI21x1_ASAP7_75t_L g3125 ( 
.A1(n_2529),
.A2(n_410),
.B(n_411),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2325),
.B(n_410),
.Y(n_3126)
);

BUFx2_ASAP7_75t_L g3127 ( 
.A(n_2563),
.Y(n_3127)
);

OR2x2_ASAP7_75t_L g3128 ( 
.A(n_2308),
.B(n_411),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2555),
.B(n_412),
.Y(n_3129)
);

INVx3_ASAP7_75t_SL g3130 ( 
.A(n_2453),
.Y(n_3130)
);

INVx4_ASAP7_75t_L g3131 ( 
.A(n_2578),
.Y(n_3131)
);

BUFx6f_ASAP7_75t_L g3132 ( 
.A(n_2751),
.Y(n_3132)
);

NOR2xp33_ASAP7_75t_L g3133 ( 
.A(n_2331),
.B(n_414),
.Y(n_3133)
);

AOI21xp5_ASAP7_75t_L g3134 ( 
.A1(n_2381),
.A2(n_414),
.B(n_415),
.Y(n_3134)
);

CKINVDCx20_ASAP7_75t_R g3135 ( 
.A(n_2506),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2576),
.B(n_414),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2592),
.B(n_415),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_SL g3138 ( 
.A(n_2751),
.B(n_643),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2613),
.B(n_416),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2660),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2521),
.Y(n_3141)
);

BUFx3_ASAP7_75t_L g3142 ( 
.A(n_2480),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2550),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_2622),
.B(n_416),
.Y(n_3144)
);

AOI22xp5_ASAP7_75t_L g3145 ( 
.A1(n_2388),
.A2(n_419),
.B1(n_417),
.B2(n_418),
.Y(n_3145)
);

A2O1A1Ixp33_ASAP7_75t_SL g3146 ( 
.A1(n_2501),
.A2(n_420),
.B(n_417),
.C(n_419),
.Y(n_3146)
);

NOR3xp33_ASAP7_75t_SL g3147 ( 
.A(n_2726),
.B(n_420),
.C(n_421),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2664),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_L g3149 ( 
.A(n_2376),
.B(n_421),
.Y(n_3149)
);

A2O1A1Ixp33_ASAP7_75t_L g3150 ( 
.A1(n_2815),
.A2(n_424),
.B(n_422),
.C(n_423),
.Y(n_3150)
);

NOR2xp33_ASAP7_75t_L g3151 ( 
.A(n_2336),
.B(n_2464),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2446),
.B(n_423),
.Y(n_3152)
);

AND2x4_ASAP7_75t_L g3153 ( 
.A(n_2624),
.B(n_423),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_SL g3154 ( 
.A(n_2772),
.B(n_644),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2342),
.B(n_424),
.Y(n_3155)
);

AOI22xp5_ASAP7_75t_L g3156 ( 
.A1(n_2560),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_3156)
);

BUFx2_ASAP7_75t_L g3157 ( 
.A(n_2399),
.Y(n_3157)
);

AO22x1_ASAP7_75t_L g3158 ( 
.A1(n_2593),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2678),
.Y(n_3159)
);

AOI21xp5_ASAP7_75t_L g3160 ( 
.A1(n_2338),
.A2(n_428),
.B(n_429),
.Y(n_3160)
);

OAI22xp5_ASAP7_75t_L g3161 ( 
.A1(n_2685),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2689),
.Y(n_3162)
);

OR2x6_ASAP7_75t_L g3163 ( 
.A(n_2578),
.B(n_430),
.Y(n_3163)
);

BUFx6f_ASAP7_75t_L g3164 ( 
.A(n_2772),
.Y(n_3164)
);

O2A1O1Ixp33_ASAP7_75t_L g3165 ( 
.A1(n_2671),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2454),
.A2(n_2355),
.B(n_2352),
.Y(n_3166)
);

AOI21x1_ASAP7_75t_L g3167 ( 
.A1(n_2307),
.A2(n_432),
.B(n_433),
.Y(n_3167)
);

INVx1_ASAP7_75t_SL g3168 ( 
.A(n_2545),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_SL g3169 ( 
.A(n_2772),
.B(n_645),
.Y(n_3169)
);

A2O1A1Ixp33_ASAP7_75t_L g3170 ( 
.A1(n_2431),
.A2(n_434),
.B(n_432),
.C(n_433),
.Y(n_3170)
);

O2A1O1Ixp33_ASAP7_75t_SL g3171 ( 
.A1(n_2457),
.A2(n_437),
.B(n_435),
.C(n_436),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_2690),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2440),
.B(n_435),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2321),
.B(n_436),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2693),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2362),
.A2(n_437),
.B(n_438),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2322),
.B(n_2326),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2427),
.B(n_437),
.Y(n_3178)
);

OAI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2701),
.A2(n_2711),
.B1(n_2714),
.B2(n_2709),
.Y(n_3179)
);

INVx3_ASAP7_75t_L g3180 ( 
.A(n_2624),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2333),
.B(n_438),
.Y(n_3181)
);

INVx4_ASAP7_75t_L g3182 ( 
.A(n_2809),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_SL g3183 ( 
.A(n_2809),
.B(n_645),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2716),
.Y(n_3184)
);

INVx3_ASAP7_75t_L g3185 ( 
.A(n_2399),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2717),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_2703),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2734),
.A2(n_439),
.B(n_440),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2565),
.A2(n_439),
.B(n_440),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2335),
.B(n_440),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2351),
.A2(n_2356),
.B(n_2614),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2568),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2618),
.A2(n_441),
.B(n_442),
.Y(n_3193)
);

NOR3xp33_ASAP7_75t_SL g3194 ( 
.A(n_2507),
.B(n_441),
.C(n_442),
.Y(n_3194)
);

BUFx3_ASAP7_75t_L g3195 ( 
.A(n_2461),
.Y(n_3195)
);

BUFx6f_ASAP7_75t_L g3196 ( 
.A(n_2809),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2599),
.Y(n_3197)
);

INVx2_ASAP7_75t_SL g3198 ( 
.A(n_2407),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2337),
.B(n_441),
.Y(n_3199)
);

BUFx3_ASAP7_75t_L g3200 ( 
.A(n_2407),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2344),
.B(n_442),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2500),
.B(n_443),
.Y(n_3202)
);

BUFx6f_ASAP7_75t_L g3203 ( 
.A(n_2615),
.Y(n_3203)
);

NOR2xp33_ASAP7_75t_L g3204 ( 
.A(n_2608),
.B(n_443),
.Y(n_3204)
);

NOR2xp67_ASAP7_75t_L g3205 ( 
.A(n_2507),
.B(n_443),
.Y(n_3205)
);

BUFx12f_ASAP7_75t_L g3206 ( 
.A(n_2615),
.Y(n_3206)
);

AOI21xp33_ASAP7_75t_L g3207 ( 
.A1(n_2586),
.A2(n_444),
.B(n_445),
.Y(n_3207)
);

AOI21xp5_ASAP7_75t_L g3208 ( 
.A1(n_2625),
.A2(n_444),
.B(n_445),
.Y(n_3208)
);

BUFx6f_ASAP7_75t_L g3209 ( 
.A(n_2380),
.Y(n_3209)
);

OAI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_2725),
.A2(n_447),
.B1(n_444),
.B2(n_446),
.Y(n_3210)
);

BUFx6f_ASAP7_75t_L g3211 ( 
.A(n_2380),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2742),
.B(n_446),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_2750),
.Y(n_3213)
);

INVx1_ASAP7_75t_SL g3214 ( 
.A(n_2435),
.Y(n_3214)
);

BUFx4_ASAP7_75t_SL g3215 ( 
.A(n_2626),
.Y(n_3215)
);

NAND3xp33_ASAP7_75t_SL g3216 ( 
.A(n_2590),
.B(n_447),
.C(n_448),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_2756),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_2762),
.B(n_447),
.Y(n_3218)
);

BUFx2_ASAP7_75t_SL g3219 ( 
.A(n_2435),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_SL g3220 ( 
.A(n_2358),
.B(n_646),
.Y(n_3220)
);

BUFx2_ASAP7_75t_L g3221 ( 
.A(n_2444),
.Y(n_3221)
);

O2A1O1Ixp33_ASAP7_75t_L g3222 ( 
.A1(n_2673),
.A2(n_450),
.B(n_448),
.C(n_449),
.Y(n_3222)
);

OAI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_2758),
.A2(n_451),
.B1(n_449),
.B2(n_450),
.Y(n_3223)
);

INVxp67_ASAP7_75t_L g3224 ( 
.A(n_2561),
.Y(n_3224)
);

NOR2xp33_ASAP7_75t_L g3225 ( 
.A(n_2490),
.B(n_449),
.Y(n_3225)
);

NAND2xp33_ASAP7_75t_L g3226 ( 
.A(n_2628),
.B(n_451),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_SL g3227 ( 
.A(n_2444),
.B(n_648),
.Y(n_3227)
);

INVxp67_ASAP7_75t_L g3228 ( 
.A(n_2584),
.Y(n_3228)
);

OAI21x1_ASAP7_75t_L g3229 ( 
.A1(n_2360),
.A2(n_451),
.B(n_452),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_2599),
.Y(n_3230)
);

NOR2xp33_ASAP7_75t_L g3231 ( 
.A(n_2350),
.B(n_452),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2393),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2763),
.B(n_453),
.Y(n_3233)
);

O2A1O1Ixp33_ASAP7_75t_L g3234 ( 
.A1(n_2687),
.A2(n_455),
.B(n_453),
.C(n_454),
.Y(n_3234)
);

OAI21xp33_ASAP7_75t_SL g3235 ( 
.A1(n_2400),
.A2(n_455),
.B(n_456),
.Y(n_3235)
);

AO21x1_ASAP7_75t_L g3236 ( 
.A1(n_2639),
.A2(n_649),
.B(n_648),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2788),
.B(n_456),
.Y(n_3237)
);

AOI21x1_ASAP7_75t_L g3238 ( 
.A1(n_2682),
.A2(n_456),
.B(n_457),
.Y(n_3238)
);

INVx2_ASAP7_75t_L g3239 ( 
.A(n_2482),
.Y(n_3239)
);

HB1xp67_ASAP7_75t_L g3240 ( 
.A(n_2466),
.Y(n_3240)
);

INVx1_ASAP7_75t_SL g3241 ( 
.A(n_2466),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2805),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_SL g3243 ( 
.A(n_2628),
.B(n_649),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2806),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_SL g3245 ( 
.A(n_2628),
.B(n_650),
.Y(n_3245)
);

A2O1A1Ixp33_ASAP7_75t_L g3246 ( 
.A1(n_2433),
.A2(n_459),
.B(n_457),
.C(n_458),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2574),
.B(n_457),
.Y(n_3247)
);

O2A1O1Ixp33_ASAP7_75t_L g3248 ( 
.A1(n_2738),
.A2(n_462),
.B(n_460),
.C(n_461),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2677),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_2823),
.B(n_651),
.Y(n_3250)
);

NOR3xp33_ASAP7_75t_L g3251 ( 
.A(n_2452),
.B(n_460),
.C(n_462),
.Y(n_3251)
);

INVx3_ASAP7_75t_L g3252 ( 
.A(n_2619),
.Y(n_3252)
);

AOI22xp5_ASAP7_75t_SL g3253 ( 
.A1(n_2600),
.A2(n_463),
.B1(n_460),
.B2(n_462),
.Y(n_3253)
);

INVx2_ASAP7_75t_SL g3254 ( 
.A(n_2340),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_2439),
.B(n_463),
.Y(n_3255)
);

AOI21x1_ASAP7_75t_L g3256 ( 
.A1(n_2641),
.A2(n_463),
.B(n_464),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_2359),
.A2(n_2647),
.B(n_2646),
.Y(n_3257)
);

INVx4_ASAP7_75t_L g3258 ( 
.A(n_2585),
.Y(n_3258)
);

NOR2xp33_ASAP7_75t_SL g3259 ( 
.A(n_2616),
.B(n_2636),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2577),
.B(n_464),
.Y(n_3260)
);

O2A1O1Ixp33_ASAP7_75t_L g3261 ( 
.A1(n_2745),
.A2(n_466),
.B(n_464),
.C(n_465),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_2825),
.B(n_465),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2598),
.Y(n_3263)
);

AOI21xp5_ASAP7_75t_L g3264 ( 
.A1(n_2648),
.A2(n_465),
.B(n_466),
.Y(n_3264)
);

INVx2_ASAP7_75t_L g3265 ( 
.A(n_2779),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_SL g3266 ( 
.A(n_2830),
.B(n_652),
.Y(n_3266)
);

INVx6_ASAP7_75t_L g3267 ( 
.A(n_2445),
.Y(n_3267)
);

AOI21x1_ASAP7_75t_L g3268 ( 
.A1(n_2654),
.A2(n_466),
.B(n_467),
.Y(n_3268)
);

A2O1A1Ixp33_ASAP7_75t_L g3269 ( 
.A1(n_2447),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_3269)
);

O2A1O1Ixp33_ASAP7_75t_L g3270 ( 
.A1(n_2765),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_3270)
);

OAI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_2838),
.A2(n_470),
.B1(n_468),
.B2(n_469),
.Y(n_3271)
);

AOI21x1_ASAP7_75t_L g3272 ( 
.A1(n_2662),
.A2(n_471),
.B(n_472),
.Y(n_3272)
);

INVx5_ASAP7_75t_L g3273 ( 
.A(n_2629),
.Y(n_3273)
);

BUFx6f_ASAP7_75t_L g3274 ( 
.A(n_2623),
.Y(n_3274)
);

BUFx6f_ASAP7_75t_L g3275 ( 
.A(n_2385),
.Y(n_3275)
);

A2O1A1Ixp33_ASAP7_75t_L g3276 ( 
.A1(n_2476),
.A2(n_2483),
.B(n_2589),
.C(n_2587),
.Y(n_3276)
);

OA22x2_ASAP7_75t_L g3277 ( 
.A1(n_2510),
.A2(n_473),
.B1(n_471),
.B2(n_472),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2526),
.Y(n_3278)
);

OAI22x1_ASAP7_75t_L g3279 ( 
.A1(n_2769),
.A2(n_474),
.B1(n_471),
.B2(n_473),
.Y(n_3279)
);

INVxp67_ASAP7_75t_L g3280 ( 
.A(n_2530),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2403),
.B(n_473),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_2395),
.B(n_652),
.Y(n_3282)
);

A2O1A1Ixp33_ASAP7_75t_L g3283 ( 
.A1(n_2567),
.A2(n_476),
.B(n_474),
.C(n_475),
.Y(n_3283)
);

BUFx2_ASAP7_75t_L g3284 ( 
.A(n_2604),
.Y(n_3284)
);

INVx5_ASAP7_75t_L g3285 ( 
.A(n_2629),
.Y(n_3285)
);

BUFx6f_ASAP7_75t_L g3286 ( 
.A(n_2424),
.Y(n_3286)
);

NOR2xp67_ASAP7_75t_SL g3287 ( 
.A(n_2395),
.B(n_476),
.Y(n_3287)
);

O2A1O1Ixp33_ASAP7_75t_L g3288 ( 
.A1(n_2816),
.A2(n_480),
.B(n_477),
.C(n_479),
.Y(n_3288)
);

O2A1O1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_2826),
.A2(n_480),
.B(n_477),
.C(n_479),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_2778),
.A2(n_481),
.B1(n_477),
.B2(n_479),
.Y(n_3290)
);

OAI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_2789),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_3291)
);

NAND2xp33_ASAP7_75t_SL g3292 ( 
.A(n_2832),
.B(n_481),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_2420),
.B(n_482),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_2947),
.A2(n_2668),
.B(n_2666),
.Y(n_3294)
);

OAI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_2841),
.A2(n_2583),
.B(n_2423),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_2842),
.Y(n_3296)
);

O2A1O1Ixp33_ASAP7_75t_L g3297 ( 
.A1(n_3179),
.A2(n_2540),
.B(n_2485),
.C(n_2822),
.Y(n_3297)
);

OAI21x1_ASAP7_75t_L g3298 ( 
.A1(n_3192),
.A2(n_2684),
.B(n_2679),
.Y(n_3298)
);

A2O1A1Ixp33_ASAP7_75t_L g3299 ( 
.A1(n_2843),
.A2(n_2658),
.B(n_2719),
.C(n_2710),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3051),
.B(n_2417),
.Y(n_3300)
);

OAI21x1_ASAP7_75t_L g3301 ( 
.A1(n_3187),
.A2(n_2696),
.B(n_2691),
.Y(n_3301)
);

AOI21x1_ASAP7_75t_L g3302 ( 
.A1(n_3197),
.A2(n_2704),
.B(n_2700),
.Y(n_3302)
);

OAI21x1_ASAP7_75t_L g3303 ( 
.A1(n_3257),
.A2(n_2715),
.B(n_2705),
.Y(n_3303)
);

NAND2x1p5_ASAP7_75t_L g3304 ( 
.A(n_2868),
.B(n_2606),
.Y(n_3304)
);

O2A1O1Ixp33_ASAP7_75t_SL g3305 ( 
.A1(n_2886),
.A2(n_2707),
.B(n_2785),
.C(n_2775),
.Y(n_3305)
);

NAND2x1p5_ASAP7_75t_L g3306 ( 
.A(n_2960),
.B(n_2486),
.Y(n_3306)
);

OAI22xp5_ASAP7_75t_L g3307 ( 
.A1(n_2844),
.A2(n_2603),
.B1(n_2803),
.B2(n_2463),
.Y(n_3307)
);

AOI221x1_ASAP7_75t_L g3308 ( 
.A1(n_2917),
.A2(n_2915),
.B1(n_2913),
.B2(n_3216),
.C(n_3150),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_2961),
.A2(n_2722),
.B(n_2720),
.Y(n_3309)
);

OAI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_2844),
.A2(n_2491),
.B1(n_2735),
.B2(n_2728),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_2896),
.B(n_2456),
.Y(n_3311)
);

OAI21x1_ASAP7_75t_L g3312 ( 
.A1(n_3230),
.A2(n_3094),
.B(n_3232),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3151),
.B(n_2386),
.Y(n_3313)
);

AOI21xp33_ASAP7_75t_L g3314 ( 
.A1(n_3022),
.A2(n_2804),
.B(n_2796),
.Y(n_3314)
);

AND2x4_ASAP7_75t_L g3315 ( 
.A(n_2973),
.B(n_2621),
.Y(n_3315)
);

OAI21x1_ASAP7_75t_L g3316 ( 
.A1(n_3239),
.A2(n_2739),
.B(n_2737),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_2859),
.Y(n_3317)
);

OR2x6_ASAP7_75t_L g3318 ( 
.A(n_2871),
.B(n_2499),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2969),
.A2(n_2743),
.B(n_2740),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_3090),
.A2(n_2755),
.B(n_2747),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2861),
.Y(n_3321)
);

BUFx6f_ASAP7_75t_L g3322 ( 
.A(n_2884),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3120),
.A2(n_2760),
.B(n_2757),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3084),
.B(n_2617),
.Y(n_3324)
);

AND2x4_ASAP7_75t_L g3325 ( 
.A(n_2973),
.B(n_2508),
.Y(n_3325)
);

NAND2x1p5_ASAP7_75t_L g3326 ( 
.A(n_3064),
.B(n_2516),
.Y(n_3326)
);

OAI21x1_ASAP7_75t_L g3327 ( 
.A1(n_3249),
.A2(n_2764),
.B(n_2761),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_2931),
.B(n_483),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3053),
.B(n_2520),
.Y(n_3329)
);

O2A1O1Ixp33_ASAP7_75t_L g3330 ( 
.A1(n_3146),
.A2(n_2415),
.B(n_2596),
.C(n_2559),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_3276),
.A2(n_2770),
.B(n_2766),
.Y(n_3331)
);

BUFx3_ASAP7_75t_L g3332 ( 
.A(n_3135),
.Y(n_3332)
);

AO32x2_ASAP7_75t_L g3333 ( 
.A1(n_3062),
.A2(n_2839),
.A3(n_3080),
.B1(n_2978),
.B2(n_3009),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3166),
.A2(n_2780),
.B(n_2771),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3089),
.B(n_2311),
.Y(n_3335)
);

AO31x2_ASAP7_75t_L g3336 ( 
.A1(n_3095),
.A2(n_3097),
.A3(n_3236),
.B(n_3045),
.Y(n_3336)
);

INVxp67_ASAP7_75t_L g3337 ( 
.A(n_2870),
.Y(n_3337)
);

AOI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_3063),
.A2(n_2595),
.B1(n_2588),
.B2(n_2551),
.Y(n_3338)
);

OAI21x1_ASAP7_75t_L g3339 ( 
.A1(n_3015),
.A2(n_2791),
.B(n_2781),
.Y(n_3339)
);

NOR2xp33_ASAP7_75t_L g3340 ( 
.A(n_3007),
.B(n_2627),
.Y(n_3340)
);

NAND3xp33_ASAP7_75t_L g3341 ( 
.A(n_2956),
.B(n_2497),
.C(n_2429),
.Y(n_3341)
);

AOI21xp5_ASAP7_75t_L g3342 ( 
.A1(n_2900),
.A2(n_2800),
.B(n_2799),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_2935),
.B(n_483),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2874),
.Y(n_3344)
);

A2O1A1Ixp33_ASAP7_75t_L g3345 ( 
.A1(n_3040),
.A2(n_2897),
.B(n_3253),
.C(n_3004),
.Y(n_3345)
);

OR2x2_ASAP7_75t_L g3346 ( 
.A(n_2850),
.B(n_2426),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3111),
.B(n_2318),
.Y(n_3347)
);

INVx2_ASAP7_75t_SL g3348 ( 
.A(n_3102),
.Y(n_3348)
);

OAI21x1_ASAP7_75t_L g3349 ( 
.A1(n_2982),
.A2(n_2835),
.B(n_2833),
.Y(n_3349)
);

OAI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_2979),
.A2(n_2837),
.B(n_2607),
.Y(n_3350)
);

AOI21xp5_ASAP7_75t_L g3351 ( 
.A1(n_3191),
.A2(n_2575),
.B(n_2558),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3104),
.B(n_2570),
.Y(n_3352)
);

AND2x6_ASAP7_75t_L g3353 ( 
.A(n_3066),
.B(n_2411),
.Y(n_3353)
);

NAND3xp33_ASAP7_75t_L g3354 ( 
.A(n_3081),
.B(n_2564),
.C(n_2462),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2880),
.Y(n_3355)
);

AOI21xp5_ASAP7_75t_L g3356 ( 
.A1(n_2926),
.A2(n_2949),
.B(n_3259),
.Y(n_3356)
);

A2O1A1Ixp33_ASAP7_75t_L g3357 ( 
.A1(n_2998),
.A2(n_2531),
.B(n_2536),
.C(n_2459),
.Y(n_3357)
);

OAI21x1_ASAP7_75t_L g3358 ( 
.A1(n_3049),
.A2(n_2579),
.B(n_2541),
.Y(n_3358)
);

INVx2_ASAP7_75t_SL g3359 ( 
.A(n_2860),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3059),
.B(n_2597),
.Y(n_3360)
);

OAI22xp5_ASAP7_75t_L g3361 ( 
.A1(n_3038),
.A2(n_2611),
.B1(n_2610),
.B2(n_486),
.Y(n_3361)
);

AO31x2_ASAP7_75t_L g3362 ( 
.A1(n_2851),
.A2(n_486),
.A3(n_484),
.B(n_485),
.Y(n_3362)
);

OAI21x1_ASAP7_75t_SL g3363 ( 
.A1(n_3035),
.A2(n_3092),
.B(n_3016),
.Y(n_3363)
);

NOR2xp67_ASAP7_75t_L g3364 ( 
.A(n_2879),
.B(n_484),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_2981),
.A2(n_3163),
.B1(n_2994),
.B2(n_3055),
.Y(n_3365)
);

AO31x2_ASAP7_75t_L g3366 ( 
.A1(n_3008),
.A2(n_488),
.A3(n_485),
.B(n_487),
.Y(n_3366)
);

AOI21x1_ASAP7_75t_L g3367 ( 
.A1(n_3238),
.A2(n_654),
.B(n_653),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3209),
.B(n_487),
.Y(n_3368)
);

AO32x2_ASAP7_75t_L g3369 ( 
.A1(n_2929),
.A2(n_491),
.A3(n_488),
.B1(n_489),
.B2(n_492),
.Y(n_3369)
);

INVx2_ASAP7_75t_L g3370 ( 
.A(n_2903),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_2946),
.A2(n_3226),
.B(n_2955),
.Y(n_3371)
);

OAI21x1_ASAP7_75t_L g3372 ( 
.A1(n_3010),
.A2(n_3083),
.B(n_3125),
.Y(n_3372)
);

HB1xp67_ASAP7_75t_L g3373 ( 
.A(n_2877),
.Y(n_3373)
);

NAND2xp5_ASAP7_75t_L g3374 ( 
.A(n_2902),
.B(n_488),
.Y(n_3374)
);

A2O1A1Ixp33_ASAP7_75t_L g3375 ( 
.A1(n_2966),
.A2(n_493),
.B(n_491),
.C(n_492),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_SL g3376 ( 
.A(n_3209),
.B(n_491),
.Y(n_3376)
);

CKINVDCx16_ASAP7_75t_R g3377 ( 
.A(n_2909),
.Y(n_3377)
);

INVx5_ASAP7_75t_L g3378 ( 
.A(n_2871),
.Y(n_3378)
);

AOI21xp5_ASAP7_75t_L g3379 ( 
.A1(n_2946),
.A2(n_493),
.B(n_494),
.Y(n_3379)
);

O2A1O1Ixp33_ASAP7_75t_SL g3380 ( 
.A1(n_2985),
.A2(n_496),
.B(n_494),
.C(n_495),
.Y(n_3380)
);

AOI21x1_ASAP7_75t_L g3381 ( 
.A1(n_3284),
.A2(n_656),
.B(n_655),
.Y(n_3381)
);

NOR2xp33_ASAP7_75t_L g3382 ( 
.A(n_3224),
.B(n_495),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2906),
.Y(n_3383)
);

OAI21x1_ASAP7_75t_L g3384 ( 
.A1(n_3265),
.A2(n_497),
.B(n_496),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_2904),
.Y(n_3385)
);

NAND3xp33_ASAP7_75t_L g3386 ( 
.A(n_3030),
.B(n_495),
.C(n_496),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_2989),
.Y(n_3387)
);

AND2x4_ASAP7_75t_L g3388 ( 
.A(n_2869),
.B(n_497),
.Y(n_3388)
);

CKINVDCx5p33_ASAP7_75t_R g3389 ( 
.A(n_2885),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_2867),
.Y(n_3390)
);

NAND3xp33_ASAP7_75t_L g3391 ( 
.A(n_3073),
.B(n_498),
.C(n_499),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3043),
.B(n_499),
.Y(n_3392)
);

INVx4_ASAP7_75t_L g3393 ( 
.A(n_3065),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2907),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2963),
.B(n_499),
.Y(n_3395)
);

AOI22xp5_ASAP7_75t_L g3396 ( 
.A1(n_3133),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_3396)
);

O2A1O1Ixp33_ASAP7_75t_SL g3397 ( 
.A1(n_3282),
.A2(n_504),
.B(n_502),
.C(n_503),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2936),
.Y(n_3398)
);

INVx3_ASAP7_75t_L g3399 ( 
.A(n_2860),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_L g3400 ( 
.A(n_3228),
.B(n_502),
.Y(n_3400)
);

OAI21x1_ASAP7_75t_L g3401 ( 
.A1(n_3017),
.A2(n_506),
.B(n_505),
.Y(n_3401)
);

OAI21x1_ASAP7_75t_L g3402 ( 
.A1(n_3229),
.A2(n_508),
.B(n_507),
.Y(n_3402)
);

O2A1O1Ixp33_ASAP7_75t_L g3403 ( 
.A1(n_3177),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_SL g3404 ( 
.A1(n_3163),
.A2(n_2873),
.B(n_3020),
.Y(n_3404)
);

A2O1A1Ixp33_ASAP7_75t_L g3405 ( 
.A1(n_2953),
.A2(n_510),
.B(n_507),
.C(n_509),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3050),
.B(n_509),
.Y(n_3406)
);

OAI21x1_ASAP7_75t_L g3407 ( 
.A1(n_3076),
.A2(n_513),
.B(n_512),
.Y(n_3407)
);

AO31x2_ASAP7_75t_L g3408 ( 
.A1(n_3278),
.A2(n_513),
.A3(n_511),
.B(n_512),
.Y(n_3408)
);

NOR2xp33_ASAP7_75t_SL g3409 ( 
.A(n_3093),
.B(n_511),
.Y(n_3409)
);

NAND2x1p5_ASAP7_75t_L g3410 ( 
.A(n_3012),
.B(n_511),
.Y(n_3410)
);

OAI21xp5_ASAP7_75t_L g3411 ( 
.A1(n_3037),
.A2(n_514),
.B(n_515),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_2943),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2944),
.Y(n_3413)
);

AOI22xp5_ASAP7_75t_L g3414 ( 
.A1(n_2924),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3124),
.B(n_514),
.Y(n_3415)
);

AOI221x1_ASAP7_75t_L g3416 ( 
.A1(n_3069),
.A2(n_518),
.B1(n_516),
.B2(n_517),
.C(n_519),
.Y(n_3416)
);

OA21x2_ASAP7_75t_L g3417 ( 
.A1(n_2934),
.A2(n_517),
.B(n_518),
.Y(n_3417)
);

OAI21x1_ASAP7_75t_L g3418 ( 
.A1(n_3256),
.A2(n_3272),
.B(n_3268),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3140),
.B(n_517),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_3148),
.A2(n_518),
.B(n_519),
.Y(n_3420)
);

OAI21x1_ASAP7_75t_L g3421 ( 
.A1(n_3096),
.A2(n_522),
.B(n_521),
.Y(n_3421)
);

NAND2x1_ASAP7_75t_SL g3422 ( 
.A(n_3130),
.B(n_2873),
.Y(n_3422)
);

OAI21xp5_ASAP7_75t_L g3423 ( 
.A1(n_3072),
.A2(n_520),
.B(n_522),
.Y(n_3423)
);

NOR2xp33_ASAP7_75t_L g3424 ( 
.A(n_3002),
.B(n_523),
.Y(n_3424)
);

CKINVDCx20_ASAP7_75t_R g3425 ( 
.A(n_3052),
.Y(n_3425)
);

AOI21xp5_ASAP7_75t_L g3426 ( 
.A1(n_3159),
.A2(n_524),
.B(n_525),
.Y(n_3426)
);

AOI21xp33_ASAP7_75t_L g3427 ( 
.A1(n_3162),
.A2(n_524),
.B(n_525),
.Y(n_3427)
);

AOI31xp67_ASAP7_75t_L g3428 ( 
.A1(n_3263),
.A2(n_3138),
.A3(n_3154),
.B(n_3088),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3172),
.B(n_526),
.Y(n_3429)
);

OAI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3027),
.A2(n_526),
.B(n_527),
.Y(n_3430)
);

O2A1O1Ixp33_ASAP7_75t_SL g3431 ( 
.A1(n_2958),
.A2(n_530),
.B(n_527),
.C(n_529),
.Y(n_3431)
);

A2O1A1Ixp33_ASAP7_75t_L g3432 ( 
.A1(n_2939),
.A2(n_531),
.B(n_529),
.C(n_530),
.Y(n_3432)
);

INVx4_ASAP7_75t_L g3433 ( 
.A(n_3024),
.Y(n_3433)
);

AO32x2_ASAP7_75t_L g3434 ( 
.A1(n_2857),
.A2(n_532),
.A3(n_529),
.B1(n_531),
.B2(n_533),
.Y(n_3434)
);

OAI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_3149),
.A2(n_531),
.B(n_532),
.Y(n_3435)
);

OAI21xp5_ASAP7_75t_SL g3436 ( 
.A1(n_3013),
.A2(n_540),
.B(n_532),
.Y(n_3436)
);

OAI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3160),
.A2(n_533),
.B(n_535),
.Y(n_3437)
);

AOI21xp5_ASAP7_75t_L g3438 ( 
.A1(n_3175),
.A2(n_3186),
.B(n_3184),
.Y(n_3438)
);

BUFx6f_ASAP7_75t_L g3439 ( 
.A(n_2932),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2983),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_2987),
.Y(n_3441)
);

AO31x2_ASAP7_75t_L g3442 ( 
.A1(n_3279),
.A2(n_537),
.A3(n_535),
.B(n_536),
.Y(n_3442)
);

AOI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3213),
.A2(n_536),
.B(n_537),
.Y(n_3443)
);

AO31x2_ASAP7_75t_L g3444 ( 
.A1(n_3182),
.A2(n_538),
.A3(n_536),
.B(n_537),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3215),
.Y(n_3445)
);

OR2x2_ASAP7_75t_L g3446 ( 
.A(n_2920),
.B(n_539),
.Y(n_3446)
);

OAI21x1_ASAP7_75t_L g3447 ( 
.A1(n_3167),
.A2(n_541),
.B(n_540),
.Y(n_3447)
);

AOI221xp5_ASAP7_75t_L g3448 ( 
.A1(n_2895),
.A2(n_542),
.B1(n_539),
.B2(n_541),
.C(n_543),
.Y(n_3448)
);

INVx2_ASAP7_75t_L g3449 ( 
.A(n_2993),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_2990),
.Y(n_3450)
);

INVx4_ASAP7_75t_L g3451 ( 
.A(n_2890),
.Y(n_3451)
);

CKINVDCx20_ASAP7_75t_R g3452 ( 
.A(n_2974),
.Y(n_3452)
);

AO31x2_ASAP7_75t_L g3453 ( 
.A1(n_3182),
.A2(n_543),
.A3(n_541),
.B(n_542),
.Y(n_3453)
);

OAI21x1_ASAP7_75t_L g3454 ( 
.A1(n_2846),
.A2(n_543),
.B(n_544),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_3217),
.B(n_544),
.Y(n_3455)
);

OAI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_2952),
.A2(n_544),
.B(n_545),
.Y(n_3456)
);

OAI21xp5_ASAP7_75t_L g3457 ( 
.A1(n_3231),
.A2(n_545),
.B(n_546),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_2855),
.Y(n_3458)
);

NAND3xp33_ASAP7_75t_SL g3459 ( 
.A(n_2875),
.B(n_546),
.C(n_547),
.Y(n_3459)
);

OR2x6_ASAP7_75t_L g3460 ( 
.A(n_3086),
.B(n_546),
.Y(n_3460)
);

CKINVDCx11_ASAP7_75t_R g3461 ( 
.A(n_3061),
.Y(n_3461)
);

CKINVDCx5p33_ASAP7_75t_R g3462 ( 
.A(n_2845),
.Y(n_3462)
);

AOI21xp5_ASAP7_75t_L g3463 ( 
.A1(n_3242),
.A2(n_547),
.B(n_548),
.Y(n_3463)
);

AOI21xp5_ASAP7_75t_L g3464 ( 
.A1(n_3244),
.A2(n_547),
.B(n_548),
.Y(n_3464)
);

BUFx2_ASAP7_75t_R g3465 ( 
.A(n_3029),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_3280),
.B(n_549),
.Y(n_3466)
);

OAI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_2996),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3032),
.Y(n_3468)
);

INVx2_ASAP7_75t_L g3469 ( 
.A(n_3036),
.Y(n_3469)
);

A2O1A1Ixp33_ASAP7_75t_L g3470 ( 
.A1(n_3122),
.A2(n_553),
.B(n_550),
.C(n_551),
.Y(n_3470)
);

AOI21xp5_ASAP7_75t_L g3471 ( 
.A1(n_2862),
.A2(n_553),
.B(n_554),
.Y(n_3471)
);

OA21x2_ASAP7_75t_L g3472 ( 
.A1(n_2957),
.A2(n_554),
.B(n_555),
.Y(n_3472)
);

AND2x4_ASAP7_75t_L g3473 ( 
.A(n_2883),
.B(n_2948),
.Y(n_3473)
);

A2O1A1Ixp33_ASAP7_75t_L g3474 ( 
.A1(n_3188),
.A2(n_557),
.B(n_555),
.C(n_556),
.Y(n_3474)
);

HB1xp67_ASAP7_75t_L g3475 ( 
.A(n_2971),
.Y(n_3475)
);

NOR2xp67_ASAP7_75t_L g3476 ( 
.A(n_2883),
.B(n_556),
.Y(n_3476)
);

AOI21x1_ASAP7_75t_L g3477 ( 
.A1(n_3078),
.A2(n_656),
.B(n_655),
.Y(n_3477)
);

OAI21x1_ASAP7_75t_L g3478 ( 
.A1(n_2846),
.A2(n_556),
.B(n_558),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_2991),
.B(n_558),
.Y(n_3479)
);

NOR2xp33_ASAP7_75t_SL g3480 ( 
.A(n_3046),
.B(n_559),
.Y(n_3480)
);

A2O1A1Ixp33_ASAP7_75t_L g3481 ( 
.A1(n_3000),
.A2(n_2959),
.B(n_3292),
.C(n_3205),
.Y(n_3481)
);

CKINVDCx11_ASAP7_75t_R g3482 ( 
.A(n_3127),
.Y(n_3482)
);

AO31x2_ASAP7_75t_L g3483 ( 
.A1(n_2865),
.A2(n_561),
.A3(n_559),
.B(n_560),
.Y(n_3483)
);

AOI221x1_ASAP7_75t_L g3484 ( 
.A1(n_2852),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.C(n_562),
.Y(n_3484)
);

INVx6_ASAP7_75t_L g3485 ( 
.A(n_3131),
.Y(n_3485)
);

O2A1O1Ixp33_ASAP7_75t_L g3486 ( 
.A1(n_2853),
.A2(n_565),
.B(n_563),
.C(n_564),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_2876),
.Y(n_3487)
);

AO31x2_ASAP7_75t_L g3488 ( 
.A1(n_2864),
.A2(n_565),
.A3(n_563),
.B(n_564),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3019),
.B(n_564),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_2891),
.Y(n_3490)
);

A2O1A1Ixp33_ASAP7_75t_L g3491 ( 
.A1(n_3119),
.A2(n_567),
.B(n_565),
.C(n_566),
.Y(n_3491)
);

O2A1O1Ixp33_ASAP7_75t_L g3492 ( 
.A1(n_3041),
.A2(n_568),
.B(n_566),
.C(n_567),
.Y(n_3492)
);

OAI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_3103),
.A2(n_570),
.B1(n_567),
.B2(n_569),
.Y(n_3493)
);

OR2x2_ASAP7_75t_L g3494 ( 
.A(n_2965),
.B(n_569),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2893),
.Y(n_3495)
);

AO32x2_ASAP7_75t_L g3496 ( 
.A1(n_2910),
.A2(n_573),
.A3(n_570),
.B1(n_571),
.B2(n_574),
.Y(n_3496)
);

AOI21xp5_ASAP7_75t_L g3497 ( 
.A1(n_3273),
.A2(n_571),
.B(n_573),
.Y(n_3497)
);

AOI21xp5_ASAP7_75t_L g3498 ( 
.A1(n_3273),
.A2(n_571),
.B(n_573),
.Y(n_3498)
);

INVx6_ASAP7_75t_L g3499 ( 
.A(n_3131),
.Y(n_3499)
);

OAI21x1_ASAP7_75t_L g3500 ( 
.A1(n_3056),
.A2(n_574),
.B(n_575),
.Y(n_3500)
);

INVx5_ASAP7_75t_L g3501 ( 
.A(n_2889),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3018),
.B(n_574),
.Y(n_3502)
);

INVxp67_ASAP7_75t_SL g3503 ( 
.A(n_3026),
.Y(n_3503)
);

O2A1O1Ixp33_ASAP7_75t_L g3504 ( 
.A1(n_3067),
.A2(n_577),
.B(n_575),
.C(n_576),
.Y(n_3504)
);

O2A1O1Ixp33_ASAP7_75t_L g3505 ( 
.A1(n_2847),
.A2(n_579),
.B(n_577),
.C(n_578),
.Y(n_3505)
);

A2O1A1Ixp33_ASAP7_75t_L g3506 ( 
.A1(n_3147),
.A2(n_580),
.B(n_578),
.C(n_579),
.Y(n_3506)
);

AOI21xp5_ASAP7_75t_L g3507 ( 
.A1(n_3273),
.A2(n_580),
.B(n_581),
.Y(n_3507)
);

O2A1O1Ixp5_ASAP7_75t_SL g3508 ( 
.A1(n_3220),
.A2(n_2976),
.B(n_3039),
.C(n_3025),
.Y(n_3508)
);

NAND2x1p5_ASAP7_75t_L g3509 ( 
.A(n_2848),
.B(n_581),
.Y(n_3509)
);

AO32x2_ASAP7_75t_L g3510 ( 
.A1(n_2911),
.A2(n_584),
.A3(n_582),
.B1(n_583),
.B2(n_585),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_3285),
.A2(n_582),
.B(n_583),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3285),
.A2(n_583),
.B(n_584),
.Y(n_3512)
);

AND2x4_ASAP7_75t_L g3513 ( 
.A(n_2948),
.B(n_584),
.Y(n_3513)
);

AOI211x1_ASAP7_75t_L g3514 ( 
.A1(n_2945),
.A2(n_587),
.B(n_585),
.C(n_586),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3204),
.B(n_585),
.Y(n_3515)
);

O2A1O1Ixp33_ASAP7_75t_L g3516 ( 
.A1(n_2863),
.A2(n_588),
.B(n_586),
.C(n_587),
.Y(n_3516)
);

INVxp67_ASAP7_75t_SL g3517 ( 
.A(n_3255),
.Y(n_3517)
);

OAI21x1_ASAP7_75t_L g3518 ( 
.A1(n_3056),
.A2(n_587),
.B(n_588),
.Y(n_3518)
);

OAI21xp5_ASAP7_75t_SL g3519 ( 
.A1(n_2975),
.A2(n_589),
.B(n_590),
.Y(n_3519)
);

BUFx3_ASAP7_75t_L g3520 ( 
.A(n_3114),
.Y(n_3520)
);

BUFx3_ASAP7_75t_L g3521 ( 
.A(n_3195),
.Y(n_3521)
);

NOR2xp33_ASAP7_75t_L g3522 ( 
.A(n_3267),
.B(n_590),
.Y(n_3522)
);

OR2x6_ASAP7_75t_L g3523 ( 
.A(n_3068),
.B(n_591),
.Y(n_3523)
);

INVx4_ASAP7_75t_L g3524 ( 
.A(n_2988),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3251),
.A2(n_594),
.B1(n_592),
.B2(n_593),
.Y(n_3525)
);

AOI21xp5_ASAP7_75t_L g3526 ( 
.A1(n_3100),
.A2(n_3211),
.B(n_2901),
.Y(n_3526)
);

AOI21xp5_ASAP7_75t_L g3527 ( 
.A1(n_3211),
.A2(n_594),
.B(n_595),
.Y(n_3527)
);

AND2x2_ASAP7_75t_L g3528 ( 
.A(n_3103),
.B(n_595),
.Y(n_3528)
);

BUFx6f_ASAP7_75t_L g3529 ( 
.A(n_3206),
.Y(n_3529)
);

AOI221xp5_ASAP7_75t_SL g3530 ( 
.A1(n_3189),
.A2(n_598),
.B1(n_596),
.B2(n_597),
.C(n_599),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2898),
.B(n_596),
.Y(n_3531)
);

AO31x2_ASAP7_75t_L g3532 ( 
.A1(n_2888),
.A2(n_599),
.A3(n_597),
.B(n_598),
.Y(n_3532)
);

CKINVDCx6p67_ASAP7_75t_R g3533 ( 
.A(n_3142),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_2872),
.Y(n_3534)
);

OAI21xp5_ASAP7_75t_L g3535 ( 
.A1(n_3193),
.A2(n_600),
.B(n_601),
.Y(n_3535)
);

AO21x1_ASAP7_75t_L g3536 ( 
.A1(n_3108),
.A2(n_601),
.B(n_602),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_2881),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_3048),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_2887),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3079),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3128),
.B(n_603),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3054),
.B(n_604),
.Y(n_3542)
);

AO31x2_ASAP7_75t_L g3543 ( 
.A1(n_2894),
.A2(n_606),
.A3(n_604),
.B(n_605),
.Y(n_3543)
);

AND2x4_ASAP7_75t_L g3544 ( 
.A(n_2988),
.B(n_605),
.Y(n_3544)
);

AO21x1_ASAP7_75t_L g3545 ( 
.A1(n_3108),
.A2(n_607),
.B(n_608),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_SL g3546 ( 
.A(n_3075),
.B(n_607),
.Y(n_3546)
);

O2A1O1Ixp33_ASAP7_75t_SL g3547 ( 
.A1(n_3269),
.A2(n_612),
.B(n_609),
.C(n_611),
.Y(n_3547)
);

AOI21xp5_ASAP7_75t_SL g3548 ( 
.A1(n_3153),
.A2(n_609),
.B(n_611),
.Y(n_3548)
);

O2A1O1Ixp33_ASAP7_75t_L g3549 ( 
.A1(n_2878),
.A2(n_613),
.B(n_611),
.C(n_612),
.Y(n_3549)
);

AOI21xp5_ASAP7_75t_L g3550 ( 
.A1(n_3250),
.A2(n_614),
.B(n_615),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_2995),
.B(n_616),
.Y(n_3551)
);

INVx3_ASAP7_75t_L g3552 ( 
.A(n_3106),
.Y(n_3552)
);

INVxp67_ASAP7_75t_L g3553 ( 
.A(n_3060),
.Y(n_3553)
);

AO31x2_ASAP7_75t_L g3554 ( 
.A1(n_2930),
.A2(n_618),
.A3(n_616),
.B(n_617),
.Y(n_3554)
);

OR2x2_ASAP7_75t_L g3555 ( 
.A(n_2858),
.B(n_617),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3101),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3317),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3321),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_SL g3559 ( 
.A(n_3501),
.B(n_3075),
.Y(n_3559)
);

OAI21xp5_ASAP7_75t_SL g3560 ( 
.A1(n_3436),
.A2(n_3117),
.B(n_3005),
.Y(n_3560)
);

OAI22xp5_ASAP7_75t_L g3561 ( 
.A1(n_3345),
.A2(n_3194),
.B1(n_2938),
.B2(n_3277),
.Y(n_3561)
);

CKINVDCx5p33_ASAP7_75t_R g3562 ( 
.A(n_3389),
.Y(n_3562)
);

BUFx6f_ASAP7_75t_L g3563 ( 
.A(n_3485),
.Y(n_3563)
);

BUFx2_ASAP7_75t_L g3564 ( 
.A(n_3422),
.Y(n_3564)
);

INVx6_ASAP7_75t_L g3565 ( 
.A(n_3433),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3390),
.B(n_3152),
.Y(n_3566)
);

BUFx10_ASAP7_75t_L g3567 ( 
.A(n_3445),
.Y(n_3567)
);

INVx1_ASAP7_75t_SL g3568 ( 
.A(n_3482),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3344),
.Y(n_3569)
);

OAI22xp33_ASAP7_75t_L g3570 ( 
.A1(n_3409),
.A2(n_3001),
.B1(n_3121),
.B2(n_3058),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3355),
.Y(n_3571)
);

INVx3_ASAP7_75t_L g3572 ( 
.A(n_3451),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3383),
.Y(n_3573)
);

INVx4_ASAP7_75t_L g3574 ( 
.A(n_3378),
.Y(n_3574)
);

CKINVDCx11_ASAP7_75t_R g3575 ( 
.A(n_3425),
.Y(n_3575)
);

AOI22xp33_ASAP7_75t_SL g3576 ( 
.A1(n_3378),
.A2(n_2889),
.B1(n_3153),
.B2(n_3267),
.Y(n_3576)
);

OAI21xp33_ASAP7_75t_L g3577 ( 
.A1(n_3480),
.A2(n_2856),
.B(n_3225),
.Y(n_3577)
);

AOI22xp33_ASAP7_75t_L g3578 ( 
.A1(n_3363),
.A2(n_3218),
.B1(n_3291),
.B2(n_3290),
.Y(n_3578)
);

OAI22xp33_ASAP7_75t_SL g3579 ( 
.A1(n_3460),
.A2(n_3523),
.B1(n_3410),
.B2(n_3318),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3449),
.Y(n_3580)
);

OAI22xp5_ASAP7_75t_L g3581 ( 
.A1(n_3476),
.A2(n_2933),
.B1(n_2984),
.B2(n_3156),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_SL g3582 ( 
.A1(n_3473),
.A2(n_2889),
.B1(n_3168),
.B2(n_3180),
.Y(n_3582)
);

AOI22xp33_ASAP7_75t_L g3583 ( 
.A1(n_3318),
.A2(n_3307),
.B1(n_3459),
.B2(n_3310),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3469),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3296),
.Y(n_3585)
);

AND2x4_ASAP7_75t_L g3586 ( 
.A(n_3501),
.B(n_2889),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3387),
.Y(n_3587)
);

OAI22xp33_ASAP7_75t_L g3588 ( 
.A1(n_3460),
.A2(n_3145),
.B1(n_3107),
.B2(n_3116),
.Y(n_3588)
);

AOI22xp33_ASAP7_75t_SL g3589 ( 
.A1(n_3365),
.A2(n_2854),
.B1(n_3286),
.B2(n_2914),
.Y(n_3589)
);

INVx4_ASAP7_75t_SL g3590 ( 
.A(n_3523),
.Y(n_3590)
);

INVx2_ASAP7_75t_SL g3591 ( 
.A(n_3529),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_3458),
.Y(n_3592)
);

OAI22xp33_ASAP7_75t_L g3593 ( 
.A1(n_3519),
.A2(n_3271),
.B1(n_3091),
.B2(n_3161),
.Y(n_3593)
);

AOI22xp33_ASAP7_75t_L g3594 ( 
.A1(n_3448),
.A2(n_3287),
.B1(n_3247),
.B2(n_3260),
.Y(n_3594)
);

AOI22xp5_ASAP7_75t_L g3595 ( 
.A1(n_3553),
.A2(n_3513),
.B1(n_3400),
.B2(n_3382),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3394),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3461),
.A2(n_3178),
.B1(n_3126),
.B2(n_3155),
.Y(n_3597)
);

OAI22xp33_ASAP7_75t_L g3598 ( 
.A1(n_3377),
.A2(n_3098),
.B1(n_3223),
.B2(n_3210),
.Y(n_3598)
);

CKINVDCx20_ASAP7_75t_R g3599 ( 
.A(n_3452),
.Y(n_3599)
);

BUFx2_ASAP7_75t_L g3600 ( 
.A(n_3520),
.Y(n_3600)
);

BUFx3_ASAP7_75t_L g3601 ( 
.A(n_3322),
.Y(n_3601)
);

BUFx8_ASAP7_75t_SL g3602 ( 
.A(n_3462),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_SL g3603 ( 
.A1(n_3517),
.A2(n_3286),
.B1(n_3219),
.B2(n_3221),
.Y(n_3603)
);

OAI22xp5_ASAP7_75t_L g3604 ( 
.A1(n_3404),
.A2(n_3003),
.B1(n_3123),
.B2(n_3034),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3438),
.B(n_2980),
.Y(n_3605)
);

INVx1_ASAP7_75t_L g3606 ( 
.A(n_3398),
.Y(n_3606)
);

BUFx2_ASAP7_75t_L g3607 ( 
.A(n_3521),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_3340),
.A2(n_3266),
.B1(n_3202),
.B2(n_3144),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3412),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3413),
.Y(n_3610)
);

INVx2_ASAP7_75t_L g3611 ( 
.A(n_3538),
.Y(n_3611)
);

BUFx2_ASAP7_75t_L g3612 ( 
.A(n_3485),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3328),
.B(n_3110),
.Y(n_3613)
);

AOI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3361),
.A2(n_2899),
.B1(n_3139),
.B2(n_2922),
.Y(n_3614)
);

INVx3_ASAP7_75t_L g3615 ( 
.A(n_3499),
.Y(n_3615)
);

OAI21xp33_ASAP7_75t_L g3616 ( 
.A1(n_3548),
.A2(n_2967),
.B(n_2942),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3440),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_SL g3618 ( 
.A1(n_3528),
.A2(n_3286),
.B1(n_3157),
.B2(n_3235),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3540),
.Y(n_3619)
);

AOI22xp33_ASAP7_75t_L g3620 ( 
.A1(n_3354),
.A2(n_3207),
.B1(n_2921),
.B2(n_2986),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3522),
.A2(n_3137),
.B1(n_3181),
.B2(n_3174),
.Y(n_3621)
);

OAI22xp5_ASAP7_75t_L g3622 ( 
.A1(n_3364),
.A2(n_3042),
.B1(n_3070),
.B2(n_3028),
.Y(n_3622)
);

AOI22xp33_ASAP7_75t_L g3623 ( 
.A1(n_3313),
.A2(n_2977),
.B1(n_3077),
.B2(n_3057),
.Y(n_3623)
);

CKINVDCx6p67_ASAP7_75t_R g3624 ( 
.A(n_3332),
.Y(n_3624)
);

HB1xp67_ASAP7_75t_L g3625 ( 
.A(n_3373),
.Y(n_3625)
);

OAI22xp33_ASAP7_75t_L g3626 ( 
.A1(n_3414),
.A2(n_2962),
.B1(n_3136),
.B2(n_3129),
.Y(n_3626)
);

AOI22xp33_ASAP7_75t_L g3627 ( 
.A1(n_3457),
.A2(n_3173),
.B1(n_3082),
.B2(n_3099),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3556),
.Y(n_3628)
);

CKINVDCx11_ASAP7_75t_R g3629 ( 
.A(n_3393),
.Y(n_3629)
);

INVx1_ASAP7_75t_L g3630 ( 
.A(n_3441),
.Y(n_3630)
);

AOI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3466),
.A2(n_3199),
.B1(n_3201),
.B2(n_3190),
.Y(n_3631)
);

OAI21xp5_ASAP7_75t_SL g3632 ( 
.A1(n_3509),
.A2(n_3222),
.B(n_3165),
.Y(n_3632)
);

BUFx12f_ASAP7_75t_L g3633 ( 
.A(n_3439),
.Y(n_3633)
);

AOI22xp33_ASAP7_75t_L g3634 ( 
.A1(n_3324),
.A2(n_3105),
.B1(n_3109),
.B2(n_3044),
.Y(n_3634)
);

CKINVDCx20_ASAP7_75t_R g3635 ( 
.A(n_3533),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3370),
.Y(n_3636)
);

OAI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3396),
.A2(n_3113),
.B1(n_2999),
.B2(n_3031),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3450),
.Y(n_3638)
);

INVx1_ASAP7_75t_L g3639 ( 
.A(n_3468),
.Y(n_3639)
);

CKINVDCx20_ASAP7_75t_R g3640 ( 
.A(n_3439),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3385),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_L g3642 ( 
.A1(n_3314),
.A2(n_3115),
.B1(n_3293),
.B2(n_3281),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3487),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3467),
.A2(n_3033),
.B1(n_2964),
.B2(n_3212),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3490),
.Y(n_3645)
);

AOI22xp33_ASAP7_75t_L g3646 ( 
.A1(n_3391),
.A2(n_3545),
.B1(n_3536),
.B2(n_3423),
.Y(n_3646)
);

AOI22xp33_ASAP7_75t_L g3647 ( 
.A1(n_3435),
.A2(n_3237),
.B1(n_3262),
.B2(n_3233),
.Y(n_3647)
);

OAI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_3481),
.A2(n_3118),
.B1(n_3170),
.B2(n_3246),
.Y(n_3648)
);

BUFx12f_ASAP7_75t_L g3649 ( 
.A(n_3348),
.Y(n_3649)
);

BUFx2_ASAP7_75t_L g3650 ( 
.A(n_3475),
.Y(n_3650)
);

BUFx3_ASAP7_75t_L g3651 ( 
.A(n_3552),
.Y(n_3651)
);

OAI22xp5_ASAP7_75t_SL g3652 ( 
.A1(n_3524),
.A2(n_3006),
.B1(n_3085),
.B2(n_3011),
.Y(n_3652)
);

INVx1_ASAP7_75t_L g3653 ( 
.A(n_3495),
.Y(n_3653)
);

BUFx10_ASAP7_75t_L g3654 ( 
.A(n_3388),
.Y(n_3654)
);

INVxp67_ASAP7_75t_SL g3655 ( 
.A(n_3503),
.Y(n_3655)
);

OAI22xp5_ASAP7_75t_L g3656 ( 
.A1(n_3299),
.A2(n_3283),
.B1(n_2997),
.B2(n_2849),
.Y(n_3656)
);

INVxp67_ASAP7_75t_L g3657 ( 
.A(n_3406),
.Y(n_3657)
);

AOI22xp33_ASAP7_75t_SL g3658 ( 
.A1(n_3493),
.A2(n_3274),
.B1(n_3240),
.B2(n_3258),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3534),
.B(n_2905),
.Y(n_3659)
);

OAI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3470),
.A2(n_3514),
.B1(n_3525),
.B2(n_3491),
.Y(n_3660)
);

CKINVDCx16_ASAP7_75t_R g3661 ( 
.A(n_3343),
.Y(n_3661)
);

AOI22xp33_ASAP7_75t_SL g3662 ( 
.A1(n_3353),
.A2(n_3274),
.B1(n_3258),
.B2(n_3254),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3408),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_SL g3664 ( 
.A1(n_3353),
.A2(n_3241),
.B1(n_3214),
.B2(n_3047),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3408),
.Y(n_3665)
);

NAND2xp5_ASAP7_75t_L g3666 ( 
.A(n_3537),
.B(n_2908),
.Y(n_3666)
);

INVx8_ASAP7_75t_L g3667 ( 
.A(n_3544),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3483),
.Y(n_3668)
);

INVx1_ASAP7_75t_L g3669 ( 
.A(n_3483),
.Y(n_3669)
);

INVx1_ASAP7_75t_SL g3670 ( 
.A(n_3359),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3374),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3323),
.A2(n_2882),
.B(n_2866),
.Y(n_3672)
);

BUFx3_ASAP7_75t_L g3673 ( 
.A(n_3399),
.Y(n_3673)
);

INVx2_ASAP7_75t_SL g3674 ( 
.A(n_3446),
.Y(n_3674)
);

HB1xp67_ASAP7_75t_L g3675 ( 
.A(n_3337),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3454),
.Y(n_3676)
);

BUFx4f_ASAP7_75t_SL g3677 ( 
.A(n_3465),
.Y(n_3677)
);

INVx4_ASAP7_75t_L g3678 ( 
.A(n_3315),
.Y(n_3678)
);

INVx4_ASAP7_75t_L g3679 ( 
.A(n_3326),
.Y(n_3679)
);

INVxp67_ASAP7_75t_L g3680 ( 
.A(n_3494),
.Y(n_3680)
);

OAI22x1_ASAP7_75t_L g3681 ( 
.A1(n_3381),
.A2(n_3023),
.B1(n_3245),
.B2(n_3243),
.Y(n_3681)
);

BUFx10_ASAP7_75t_L g3682 ( 
.A(n_3424),
.Y(n_3682)
);

INVx2_ASAP7_75t_L g3683 ( 
.A(n_3478),
.Y(n_3683)
);

BUFx10_ASAP7_75t_L g3684 ( 
.A(n_3325),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_3444),
.Y(n_3685)
);

AOI22xp5_ASAP7_75t_L g3686 ( 
.A1(n_3539),
.A2(n_2840),
.B1(n_3158),
.B2(n_3227),
.Y(n_3686)
);

NAND2x1p5_ASAP7_75t_L g3687 ( 
.A(n_3546),
.B(n_3200),
.Y(n_3687)
);

OAI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3506),
.A2(n_3183),
.B1(n_3169),
.B2(n_2919),
.Y(n_3688)
);

INVx3_ASAP7_75t_L g3689 ( 
.A(n_3306),
.Y(n_3689)
);

CKINVDCx6p67_ASAP7_75t_R g3690 ( 
.A(n_3555),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3335),
.B(n_2923),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3453),
.Y(n_3692)
);

AOI22xp33_ASAP7_75t_L g3693 ( 
.A1(n_3386),
.A2(n_3176),
.B1(n_3208),
.B2(n_3264),
.Y(n_3693)
);

BUFx12f_ASAP7_75t_L g3694 ( 
.A(n_3304),
.Y(n_3694)
);

AOI22xp33_ASAP7_75t_L g3695 ( 
.A1(n_3456),
.A2(n_3134),
.B1(n_2927),
.B2(n_2968),
.Y(n_3695)
);

BUFx10_ASAP7_75t_L g3696 ( 
.A(n_3380),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3415),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3311),
.A2(n_2972),
.B1(n_2925),
.B2(n_2940),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3437),
.A2(n_2941),
.B1(n_2950),
.B2(n_2937),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3392),
.B(n_3112),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3419),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3542),
.B(n_3141),
.Y(n_3702)
);

BUFx8_ASAP7_75t_L g3703 ( 
.A(n_3434),
.Y(n_3703)
);

AOI22xp5_ASAP7_75t_L g3704 ( 
.A1(n_3515),
.A2(n_2918),
.B1(n_3171),
.B2(n_3252),
.Y(n_3704)
);

BUFx3_ASAP7_75t_L g3705 ( 
.A(n_3395),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3352),
.B(n_3143),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3429),
.Y(n_3707)
);

INVx2_ASAP7_75t_SL g3708 ( 
.A(n_3346),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_SL g3709 ( 
.A1(n_3417),
.A2(n_3198),
.B1(n_3185),
.B2(n_2882),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3421),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3455),
.Y(n_3711)
);

CKINVDCx5p33_ASAP7_75t_R g3712 ( 
.A(n_3479),
.Y(n_3712)
);

INVx2_ASAP7_75t_L g3713 ( 
.A(n_3447),
.Y(n_3713)
);

NAND2x1p5_ASAP7_75t_L g3714 ( 
.A(n_3368),
.B(n_2866),
.Y(n_3714)
);

CKINVDCx20_ASAP7_75t_R g3715 ( 
.A(n_3489),
.Y(n_3715)
);

AND2x2_ASAP7_75t_L g3716 ( 
.A(n_3541),
.B(n_3531),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3535),
.A2(n_3275),
.B1(n_3203),
.B2(n_2882),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3384),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_L g3719 ( 
.A1(n_3502),
.A2(n_3275),
.B1(n_3203),
.B2(n_2892),
.Y(n_3719)
);

INVx4_ASAP7_75t_L g3720 ( 
.A(n_3472),
.Y(n_3720)
);

INVxp67_ASAP7_75t_SL g3721 ( 
.A(n_3500),
.Y(n_3721)
);

CKINVDCx11_ASAP7_75t_R g3722 ( 
.A(n_3431),
.Y(n_3722)
);

BUFx12f_ASAP7_75t_L g3723 ( 
.A(n_3434),
.Y(n_3723)
);

BUFx3_ASAP7_75t_L g3724 ( 
.A(n_3401),
.Y(n_3724)
);

INVx6_ASAP7_75t_L g3725 ( 
.A(n_3376),
.Y(n_3725)
);

CKINVDCx11_ASAP7_75t_R g3726 ( 
.A(n_3527),
.Y(n_3726)
);

CKINVDCx5p33_ASAP7_75t_R g3727 ( 
.A(n_3551),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3360),
.B(n_619),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3488),
.Y(n_3729)
);

INVx2_ASAP7_75t_SL g3730 ( 
.A(n_3572),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3579),
.B(n_3356),
.Y(n_3731)
);

OAI21x1_ASAP7_75t_L g3732 ( 
.A1(n_3672),
.A2(n_3372),
.B(n_3301),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3557),
.Y(n_3733)
);

INVx2_ASAP7_75t_SL g3734 ( 
.A(n_3567),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3558),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_3681),
.A2(n_3371),
.B(n_3319),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3729),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3585),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3663),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3569),
.Y(n_3740)
);

OAI21x1_ASAP7_75t_L g3741 ( 
.A1(n_3713),
.A2(n_3312),
.B(n_3418),
.Y(n_3741)
);

OAI21x1_ASAP7_75t_L g3742 ( 
.A1(n_3718),
.A2(n_3303),
.B(n_3298),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3571),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3573),
.Y(n_3744)
);

INVx1_ASAP7_75t_L g3745 ( 
.A(n_3587),
.Y(n_3745)
);

AOI22xp33_ASAP7_75t_L g3746 ( 
.A1(n_3723),
.A2(n_3341),
.B1(n_3338),
.B2(n_3350),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3592),
.Y(n_3747)
);

BUFx6f_ASAP7_75t_L g3748 ( 
.A(n_3563),
.Y(n_3748)
);

OR2x2_ASAP7_75t_L g3749 ( 
.A(n_3661),
.B(n_3442),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3611),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3596),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_3619),
.Y(n_3752)
);

BUFx2_ASAP7_75t_L g3753 ( 
.A(n_3600),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3606),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3628),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3609),
.Y(n_3756)
);

AO31x2_ASAP7_75t_L g3757 ( 
.A1(n_3720),
.A2(n_3308),
.A3(n_3342),
.B(n_3331),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3610),
.Y(n_3758)
);

HB1xp67_ASAP7_75t_L g3759 ( 
.A(n_3655),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3613),
.B(n_3369),
.Y(n_3760)
);

INVx3_ASAP7_75t_L g3761 ( 
.A(n_3586),
.Y(n_3761)
);

INVx2_ASAP7_75t_L g3762 ( 
.A(n_3580),
.Y(n_3762)
);

BUFx3_ASAP7_75t_L g3763 ( 
.A(n_3640),
.Y(n_3763)
);

BUFx6f_ASAP7_75t_L g3764 ( 
.A(n_3563),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3617),
.Y(n_3765)
);

AND2x4_ASAP7_75t_L g3766 ( 
.A(n_3708),
.B(n_3518),
.Y(n_3766)
);

INVx2_ASAP7_75t_L g3767 ( 
.A(n_3584),
.Y(n_3767)
);

INVx1_ASAP7_75t_L g3768 ( 
.A(n_3630),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3638),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3639),
.Y(n_3770)
);

AND2x2_ASAP7_75t_L g3771 ( 
.A(n_3657),
.B(n_3369),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3643),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3645),
.Y(n_3773)
);

INVx3_ASAP7_75t_L g3774 ( 
.A(n_3586),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3653),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3636),
.Y(n_3776)
);

INVx3_ASAP7_75t_L g3777 ( 
.A(n_3684),
.Y(n_3777)
);

AND2x4_ASAP7_75t_L g3778 ( 
.A(n_3590),
.B(n_3362),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3625),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3641),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3706),
.Y(n_3781)
);

OR2x2_ASAP7_75t_L g3782 ( 
.A(n_3650),
.B(n_3362),
.Y(n_3782)
);

CKINVDCx5p33_ASAP7_75t_R g3783 ( 
.A(n_3575),
.Y(n_3783)
);

INVx1_ASAP7_75t_L g3784 ( 
.A(n_3675),
.Y(n_3784)
);

INVx3_ASAP7_75t_L g3785 ( 
.A(n_3684),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3700),
.B(n_3496),
.Y(n_3786)
);

INVx1_ASAP7_75t_L g3787 ( 
.A(n_3605),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3566),
.Y(n_3788)
);

HB1xp67_ASAP7_75t_L g3789 ( 
.A(n_3612),
.Y(n_3789)
);

CKINVDCx12_ASAP7_75t_R g3790 ( 
.A(n_3677),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3674),
.B(n_3496),
.Y(n_3791)
);

BUFx3_ASAP7_75t_L g3792 ( 
.A(n_3633),
.Y(n_3792)
);

BUFx6f_ASAP7_75t_L g3793 ( 
.A(n_3563),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_3697),
.B(n_3530),
.Y(n_3794)
);

AND2x4_ASAP7_75t_L g3795 ( 
.A(n_3590),
.B(n_3679),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3701),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3707),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3711),
.Y(n_3798)
);

INVx2_ASAP7_75t_SL g3799 ( 
.A(n_3567),
.Y(n_3799)
);

OR2x2_ASAP7_75t_L g3800 ( 
.A(n_3680),
.B(n_3366),
.Y(n_3800)
);

OAI21x1_ASAP7_75t_L g3801 ( 
.A1(n_3710),
.A2(n_3327),
.B(n_3316),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3685),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3671),
.B(n_3300),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3692),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3668),
.Y(n_3805)
);

BUFx3_ASAP7_75t_L g3806 ( 
.A(n_3635),
.Y(n_3806)
);

AOI22xp33_ASAP7_75t_L g3807 ( 
.A1(n_3604),
.A2(n_3427),
.B1(n_3295),
.B2(n_3497),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3676),
.A2(n_3351),
.B(n_3302),
.Y(n_3808)
);

HB1xp67_ASAP7_75t_L g3809 ( 
.A(n_3607),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3669),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3665),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3702),
.Y(n_3812)
);

INVx3_ASAP7_75t_L g3813 ( 
.A(n_3678),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3683),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3721),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3728),
.Y(n_3816)
);

BUFx6f_ASAP7_75t_L g3817 ( 
.A(n_3673),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3659),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3666),
.Y(n_3819)
);

BUFx3_ASAP7_75t_L g3820 ( 
.A(n_3649),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3716),
.B(n_3510),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3724),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3691),
.Y(n_3823)
);

AND2x2_ASAP7_75t_L g3824 ( 
.A(n_3705),
.B(n_3333),
.Y(n_3824)
);

INVx2_ASAP7_75t_SL g3825 ( 
.A(n_3601),
.Y(n_3825)
);

OAI21x1_ASAP7_75t_L g3826 ( 
.A1(n_3689),
.A2(n_3334),
.B(n_3358),
.Y(n_3826)
);

OA21x2_ASAP7_75t_L g3827 ( 
.A1(n_3583),
.A2(n_3560),
.B(n_3717),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3564),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3703),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3703),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3690),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3654),
.Y(n_3832)
);

BUFx6f_ASAP7_75t_L g3833 ( 
.A(n_3651),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3654),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3670),
.Y(n_3835)
);

HB1xp67_ASAP7_75t_L g3836 ( 
.A(n_3615),
.Y(n_3836)
);

AO21x2_ASAP7_75t_L g3837 ( 
.A1(n_3561),
.A2(n_3379),
.B(n_3367),
.Y(n_3837)
);

BUFx3_ASAP7_75t_L g3838 ( 
.A(n_3565),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_L g3839 ( 
.A(n_3595),
.B(n_3347),
.Y(n_3839)
);

INVx3_ASAP7_75t_L g3840 ( 
.A(n_3574),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3662),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3725),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3696),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3597),
.B(n_3333),
.Y(n_3844)
);

INVx3_ASAP7_75t_L g3845 ( 
.A(n_3694),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3725),
.Y(n_3846)
);

OR2x2_ASAP7_75t_L g3847 ( 
.A(n_3759),
.B(n_3568),
.Y(n_3847)
);

OAI22xp33_ASAP7_75t_L g3848 ( 
.A1(n_3813),
.A2(n_3614),
.B1(n_3667),
.B2(n_3686),
.Y(n_3848)
);

OR2x6_ASAP7_75t_L g3849 ( 
.A(n_3795),
.B(n_3667),
.Y(n_3849)
);

O2A1O1Ixp33_ASAP7_75t_L g3850 ( 
.A1(n_3731),
.A2(n_3588),
.B(n_3577),
.C(n_3616),
.Y(n_3850)
);

AND2x2_ASAP7_75t_L g3851 ( 
.A(n_3753),
.B(n_3682),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3733),
.Y(n_3852)
);

OA21x2_ASAP7_75t_L g3853 ( 
.A1(n_3736),
.A2(n_3719),
.B(n_3646),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3779),
.B(n_3727),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3809),
.B(n_3664),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3735),
.Y(n_3856)
);

A2O1A1Ixp33_ASAP7_75t_L g3857 ( 
.A1(n_3813),
.A2(n_3576),
.B(n_3582),
.C(n_3589),
.Y(n_3857)
);

NAND4xp25_ASAP7_75t_L g3858 ( 
.A(n_3844),
.B(n_3618),
.C(n_3608),
.D(n_3620),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3784),
.B(n_3712),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3821),
.B(n_3631),
.Y(n_3860)
);

OR2x2_ASAP7_75t_L g3861 ( 
.A(n_3787),
.B(n_3591),
.Y(n_3861)
);

AND2x4_ASAP7_75t_L g3862 ( 
.A(n_3795),
.B(n_3559),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3829),
.B(n_3624),
.Y(n_3863)
);

AOI221x1_ASAP7_75t_L g3864 ( 
.A1(n_3840),
.A2(n_3526),
.B1(n_3656),
.B2(n_3320),
.C(n_3309),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3740),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3789),
.B(n_3603),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3824),
.B(n_3621),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_3786),
.B(n_3647),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3828),
.B(n_3658),
.Y(n_3869)
);

OAI21xp5_ASAP7_75t_L g3870 ( 
.A1(n_3746),
.A2(n_3715),
.B(n_3632),
.Y(n_3870)
);

OAI21x1_ASAP7_75t_SL g3871 ( 
.A1(n_3830),
.A2(n_3477),
.B(n_3403),
.Y(n_3871)
);

OA21x2_ASAP7_75t_L g3872 ( 
.A1(n_3841),
.A2(n_3484),
.B(n_3416),
.Y(n_3872)
);

AOI221xp5_ASAP7_75t_L g3873 ( 
.A1(n_3839),
.A2(n_3570),
.B1(n_3598),
.B2(n_3593),
.C(n_3637),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3788),
.B(n_3709),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3743),
.Y(n_3875)
);

OAI22xp5_ASAP7_75t_L g3876 ( 
.A1(n_3749),
.A2(n_3578),
.B1(n_3704),
.B2(n_3687),
.Y(n_3876)
);

AOI21xp5_ASAP7_75t_L g3877 ( 
.A1(n_3841),
.A2(n_3397),
.B(n_3547),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3744),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3781),
.B(n_3488),
.Y(n_3879)
);

OA21x2_ASAP7_75t_L g3880 ( 
.A1(n_3808),
.A2(n_3402),
.B(n_3642),
.Y(n_3880)
);

INVxp67_ASAP7_75t_L g3881 ( 
.A(n_3836),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_L g3882 ( 
.A(n_3771),
.B(n_3623),
.Y(n_3882)
);

AOI221xp5_ASAP7_75t_L g3883 ( 
.A1(n_3816),
.A2(n_3486),
.B1(n_3581),
.B2(n_3626),
.C(n_3660),
.Y(n_3883)
);

BUFx2_ASAP7_75t_L g3884 ( 
.A(n_3833),
.Y(n_3884)
);

INVxp67_ASAP7_75t_L g3885 ( 
.A(n_3730),
.Y(n_3885)
);

AND2x4_ASAP7_75t_L g3886 ( 
.A(n_3777),
.B(n_3599),
.Y(n_3886)
);

BUFx3_ASAP7_75t_L g3887 ( 
.A(n_3792),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3823),
.B(n_3696),
.Y(n_3888)
);

INVx1_ASAP7_75t_SL g3889 ( 
.A(n_3838),
.Y(n_3889)
);

AND2x2_ASAP7_75t_L g3890 ( 
.A(n_3835),
.B(n_3812),
.Y(n_3890)
);

NOR2xp33_ASAP7_75t_L g3891 ( 
.A(n_3817),
.B(n_3833),
.Y(n_3891)
);

AND2x2_ASAP7_75t_L g3892 ( 
.A(n_3818),
.B(n_3726),
.Y(n_3892)
);

A2O1A1Ixp33_ASAP7_75t_L g3893 ( 
.A1(n_3777),
.A2(n_3492),
.B(n_3504),
.C(n_3297),
.Y(n_3893)
);

NAND2xp33_ASAP7_75t_L g3894 ( 
.A(n_3845),
.B(n_3562),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3819),
.B(n_3714),
.Y(n_3895)
);

AO32x1_ASAP7_75t_L g3896 ( 
.A1(n_3843),
.A2(n_3648),
.A3(n_3622),
.B1(n_3688),
.B2(n_3722),
.Y(n_3896)
);

O2A1O1Ixp33_ASAP7_75t_L g3897 ( 
.A1(n_3794),
.A2(n_3405),
.B(n_3432),
.C(n_3375),
.Y(n_3897)
);

OAI22xp5_ASAP7_75t_L g3898 ( 
.A1(n_3785),
.A2(n_3594),
.B1(n_3627),
.B2(n_3634),
.Y(n_3898)
);

AND2x4_ASAP7_75t_L g3899 ( 
.A(n_3761),
.B(n_3336),
.Y(n_3899)
);

OAI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_3778),
.A2(n_3508),
.B(n_3474),
.Y(n_3900)
);

BUFx8_ASAP7_75t_SL g3901 ( 
.A(n_3783),
.Y(n_3901)
);

A2O1A1Ixp33_ASAP7_75t_L g3902 ( 
.A1(n_3778),
.A2(n_3516),
.B(n_3549),
.C(n_3505),
.Y(n_3902)
);

OR2x2_ASAP7_75t_L g3903 ( 
.A(n_3745),
.B(n_3532),
.Y(n_3903)
);

OAI22xp5_ASAP7_75t_L g3904 ( 
.A1(n_3807),
.A2(n_3695),
.B1(n_3652),
.B2(n_3698),
.Y(n_3904)
);

INVx1_ASAP7_75t_L g3905 ( 
.A(n_3747),
.Y(n_3905)
);

INVxp67_ASAP7_75t_L g3906 ( 
.A(n_3833),
.Y(n_3906)
);

NOR2xp33_ASAP7_75t_L g3907 ( 
.A(n_3817),
.B(n_3565),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3738),
.Y(n_3908)
);

OAI21x1_ASAP7_75t_L g3909 ( 
.A1(n_3732),
.A2(n_3407),
.B(n_3498),
.Y(n_3909)
);

NOR2x1_ASAP7_75t_SL g3910 ( 
.A(n_3734),
.B(n_3799),
.Y(n_3910)
);

A2O1A1Ixp33_ASAP7_75t_L g3911 ( 
.A1(n_3840),
.A2(n_3420),
.B(n_3443),
.C(n_3426),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3827),
.A2(n_3644),
.B1(n_3699),
.B2(n_3693),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3796),
.B(n_2916),
.Y(n_3913)
);

INVx3_ASAP7_75t_SL g3914 ( 
.A(n_3820),
.Y(n_3914)
);

BUFx2_ASAP7_75t_SL g3915 ( 
.A(n_3817),
.Y(n_3915)
);

OAI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3827),
.A2(n_3511),
.B(n_3507),
.Y(n_3916)
);

A2O1A1Ixp33_ASAP7_75t_L g3917 ( 
.A1(n_3825),
.A2(n_3463),
.B(n_3464),
.C(n_3512),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3852),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3856),
.Y(n_3919)
);

OR2x2_ASAP7_75t_L g3920 ( 
.A(n_3867),
.B(n_3782),
.Y(n_3920)
);

INVxp67_ASAP7_75t_L g3921 ( 
.A(n_3910),
.Y(n_3921)
);

AOI22xp5_ASAP7_75t_L g3922 ( 
.A1(n_3873),
.A2(n_3842),
.B1(n_3846),
.B2(n_3760),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3865),
.Y(n_3923)
);

BUFx2_ASAP7_75t_L g3924 ( 
.A(n_3884),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3882),
.B(n_3800),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3851),
.B(n_3831),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3875),
.Y(n_3927)
);

OAI22xp5_ASAP7_75t_L g3928 ( 
.A1(n_3857),
.A2(n_3834),
.B1(n_3832),
.B2(n_3774),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3908),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3868),
.B(n_3791),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3890),
.B(n_3774),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3878),
.Y(n_3932)
);

OR2x2_ASAP7_75t_L g3933 ( 
.A(n_3860),
.B(n_3797),
.Y(n_3933)
);

OR2x2_ASAP7_75t_L g3934 ( 
.A(n_3905),
.B(n_3847),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3861),
.Y(n_3935)
);

OR2x2_ASAP7_75t_L g3936 ( 
.A(n_3879),
.B(n_3798),
.Y(n_3936)
);

INVx1_ASAP7_75t_L g3937 ( 
.A(n_3903),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3881),
.B(n_3822),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3899),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3874),
.B(n_3751),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3899),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3892),
.B(n_3754),
.Y(n_3942)
);

OR2x2_ASAP7_75t_L g3943 ( 
.A(n_3855),
.B(n_3756),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3913),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3895),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3866),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3869),
.B(n_3758),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3888),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3858),
.A2(n_3766),
.B1(n_3837),
.B2(n_3737),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3854),
.B(n_3859),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3906),
.Y(n_3951)
);

INVx3_ASAP7_75t_L g3952 ( 
.A(n_3849),
.Y(n_3952)
);

INVx1_ASAP7_75t_SL g3953 ( 
.A(n_3914),
.Y(n_3953)
);

INVx3_ASAP7_75t_L g3954 ( 
.A(n_3849),
.Y(n_3954)
);

HB1xp67_ASAP7_75t_L g3955 ( 
.A(n_3885),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3891),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3889),
.B(n_3765),
.Y(n_3957)
);

INVx2_ASAP7_75t_SL g3958 ( 
.A(n_3887),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3886),
.B(n_3768),
.Y(n_3959)
);

INVxp33_ASAP7_75t_L g3960 ( 
.A(n_3901),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3870),
.A2(n_3766),
.B1(n_3737),
.B2(n_3815),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3862),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3880),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3863),
.B(n_3769),
.Y(n_3964)
);

BUFx5_ASAP7_75t_L g3965 ( 
.A(n_3909),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3915),
.B(n_3770),
.Y(n_3966)
);

INVx3_ASAP7_75t_L g3967 ( 
.A(n_3853),
.Y(n_3967)
);

INVx2_ASAP7_75t_L g3968 ( 
.A(n_3880),
.Y(n_3968)
);

OR2x2_ASAP7_75t_L g3969 ( 
.A(n_3898),
.B(n_3772),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3872),
.Y(n_3970)
);

AND2x2_ASAP7_75t_L g3971 ( 
.A(n_3907),
.B(n_3773),
.Y(n_3971)
);

HB1xp67_ASAP7_75t_L g3972 ( 
.A(n_3912),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3883),
.B(n_3775),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3853),
.B(n_3780),
.Y(n_3974)
);

AOI221xp5_ASAP7_75t_L g3975 ( 
.A1(n_3972),
.A2(n_3850),
.B1(n_3848),
.B2(n_3904),
.C(n_3876),
.Y(n_3975)
);

NOR2xp33_ASAP7_75t_L g3976 ( 
.A(n_3953),
.B(n_3806),
.Y(n_3976)
);

AND2x2_ASAP7_75t_L g3977 ( 
.A(n_3962),
.B(n_3815),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3970),
.Y(n_3978)
);

INVx4_ASAP7_75t_L g3979 ( 
.A(n_3952),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3937),
.Y(n_3980)
);

INVx1_ASAP7_75t_L g3981 ( 
.A(n_3918),
.Y(n_3981)
);

AO21x2_ASAP7_75t_L g3982 ( 
.A1(n_3963),
.A2(n_3900),
.B(n_3871),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3918),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3924),
.B(n_3750),
.Y(n_3984)
);

OAI33xp33_ASAP7_75t_L g3985 ( 
.A1(n_3928),
.A2(n_3803),
.A3(n_3897),
.B1(n_3810),
.B2(n_3805),
.B3(n_3811),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3931),
.B(n_3752),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3919),
.Y(n_3987)
);

BUFx2_ASAP7_75t_L g3988 ( 
.A(n_3921),
.Y(n_3988)
);

INVx2_ASAP7_75t_L g3989 ( 
.A(n_3929),
.Y(n_3989)
);

OR2x2_ASAP7_75t_L g3990 ( 
.A(n_3925),
.B(n_3920),
.Y(n_3990)
);

NAND3xp33_ASAP7_75t_L g3991 ( 
.A(n_3949),
.B(n_3864),
.C(n_3916),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3933),
.B(n_3802),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3923),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3946),
.B(n_3755),
.Y(n_3994)
);

NOR2x1_ASAP7_75t_SL g3995 ( 
.A(n_3958),
.B(n_3763),
.Y(n_3995)
);

OR2x6_ASAP7_75t_L g3996 ( 
.A(n_3952),
.B(n_3877),
.Y(n_3996)
);

AND2x2_ASAP7_75t_L g3997 ( 
.A(n_3946),
.B(n_3762),
.Y(n_3997)
);

INVx1_ASAP7_75t_L g3998 ( 
.A(n_3927),
.Y(n_3998)
);

HB1xp67_ASAP7_75t_L g3999 ( 
.A(n_3955),
.Y(n_3999)
);

INVx1_ASAP7_75t_L g4000 ( 
.A(n_3932),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3959),
.B(n_3767),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3969),
.B(n_3872),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3948),
.B(n_3776),
.Y(n_4003)
);

HB1xp67_ASAP7_75t_L g4004 ( 
.A(n_3934),
.Y(n_4004)
);

AND2x2_ASAP7_75t_L g4005 ( 
.A(n_3935),
.B(n_3804),
.Y(n_4005)
);

INVxp67_ASAP7_75t_L g4006 ( 
.A(n_3938),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3936),
.Y(n_4007)
);

AND2x2_ASAP7_75t_L g4008 ( 
.A(n_3945),
.B(n_3739),
.Y(n_4008)
);

INVx3_ASAP7_75t_L g4009 ( 
.A(n_3954),
.Y(n_4009)
);

INVx5_ASAP7_75t_L g4010 ( 
.A(n_3967),
.Y(n_4010)
);

INVx1_ASAP7_75t_SL g4011 ( 
.A(n_3957),
.Y(n_4011)
);

INVx4_ASAP7_75t_L g4012 ( 
.A(n_3966),
.Y(n_4012)
);

INVx1_ASAP7_75t_L g4013 ( 
.A(n_3944),
.Y(n_4013)
);

OAI22xp5_ASAP7_75t_SL g4014 ( 
.A1(n_3960),
.A2(n_3790),
.B1(n_3894),
.B2(n_3629),
.Y(n_4014)
);

OAI31xp33_ASAP7_75t_SL g4015 ( 
.A1(n_3950),
.A2(n_3896),
.A3(n_3826),
.B(n_3430),
.Y(n_4015)
);

INVx3_ASAP7_75t_L g4016 ( 
.A(n_3941),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3974),
.Y(n_4017)
);

AND2x4_ASAP7_75t_L g4018 ( 
.A(n_3939),
.B(n_3757),
.Y(n_4018)
);

NOR2xp33_ASAP7_75t_L g4019 ( 
.A(n_3947),
.B(n_3602),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3978),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3979),
.B(n_3956),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3979),
.B(n_3939),
.Y(n_4022)
);

AND2x2_ASAP7_75t_L g4023 ( 
.A(n_3988),
.B(n_3942),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3978),
.B(n_3930),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3998),
.Y(n_4025)
);

OR2x2_ASAP7_75t_L g4026 ( 
.A(n_3990),
.B(n_3943),
.Y(n_4026)
);

INVx2_ASAP7_75t_L g4027 ( 
.A(n_3999),
.Y(n_4027)
);

AND2x2_ASAP7_75t_L g4028 ( 
.A(n_4009),
.B(n_3971),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_4009),
.B(n_3964),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_4002),
.B(n_3967),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_4012),
.B(n_3926),
.Y(n_4031)
);

INVx2_ASAP7_75t_L g4032 ( 
.A(n_3993),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3998),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_SL g4034 ( 
.A(n_4010),
.B(n_3965),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_4000),
.Y(n_4035)
);

OR2x2_ASAP7_75t_L g4036 ( 
.A(n_4004),
.B(n_3940),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3981),
.Y(n_4037)
);

NOR3xp33_ASAP7_75t_SL g4038 ( 
.A(n_4014),
.B(n_3902),
.C(n_3893),
.Y(n_4038)
);

BUFx2_ASAP7_75t_L g4039 ( 
.A(n_3996),
.Y(n_4039)
);

OR2x6_ASAP7_75t_L g4040 ( 
.A(n_3996),
.B(n_3968),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_4017),
.B(n_3951),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_4011),
.B(n_3961),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3980),
.B(n_3973),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3983),
.Y(n_4044)
);

AOI22xp5_ASAP7_75t_L g4045 ( 
.A1(n_3975),
.A2(n_3922),
.B1(n_3917),
.B2(n_3911),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3987),
.Y(n_4046)
);

NOR2x1_ASAP7_75t_L g4047 ( 
.A(n_3995),
.B(n_3748),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_4045),
.B(n_3980),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_4043),
.B(n_3991),
.Y(n_4049)
);

NOR3xp33_ASAP7_75t_L g4050 ( 
.A(n_4039),
.B(n_3985),
.C(n_3976),
.Y(n_4050)
);

INVx1_ASAP7_75t_L g4051 ( 
.A(n_4027),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_4037),
.Y(n_4052)
);

OR2x2_ASAP7_75t_L g4053 ( 
.A(n_4024),
.B(n_3992),
.Y(n_4053)
);

NAND3xp33_ASAP7_75t_L g4054 ( 
.A(n_4038),
.B(n_4015),
.C(n_4010),
.Y(n_4054)
);

INVx2_ASAP7_75t_L g4055 ( 
.A(n_4031),
.Y(n_4055)
);

OR2x6_ASAP7_75t_L g4056 ( 
.A(n_4047),
.B(n_4019),
.Y(n_4056)
);

INVx1_ASAP7_75t_SL g4057 ( 
.A(n_4021),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_4044),
.Y(n_4058)
);

HB1xp67_ASAP7_75t_L g4059 ( 
.A(n_4020),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_4046),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_4032),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_4042),
.B(n_3984),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_4025),
.Y(n_4063)
);

OR2x2_ASAP7_75t_L g4064 ( 
.A(n_4030),
.B(n_4013),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_4033),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_4035),
.Y(n_4066)
);

HB1xp67_ASAP7_75t_L g4067 ( 
.A(n_4040),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_L g4068 ( 
.A(n_4036),
.B(n_4018),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_4026),
.B(n_4023),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_4022),
.B(n_4007),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_4040),
.B(n_4016),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_4040),
.B(n_4016),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_4041),
.B(n_4013),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_4029),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_4028),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4034),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_4034),
.B(n_3994),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_4020),
.Y(n_4078)
);

INVx1_ASAP7_75t_L g4079 ( 
.A(n_4027),
.Y(n_4079)
);

AND2x2_ASAP7_75t_L g4080 ( 
.A(n_4056),
.B(n_3982),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_4055),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_4056),
.B(n_3982),
.Y(n_4082)
);

INVxp33_ASAP7_75t_L g4083 ( 
.A(n_4067),
.Y(n_4083)
);

INVx2_ASAP7_75t_L g4084 ( 
.A(n_4061),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_4062),
.B(n_4057),
.Y(n_4085)
);

NOR2x1_ASAP7_75t_L g4086 ( 
.A(n_4054),
.B(n_3471),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_4071),
.B(n_4006),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_4053),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_L g4089 ( 
.A(n_4050),
.B(n_3977),
.Y(n_4089)
);

AOI33xp33_ASAP7_75t_L g4090 ( 
.A1(n_4076),
.A2(n_4008),
.A3(n_4005),
.B1(n_4001),
.B2(n_4003),
.B3(n_3997),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4059),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_4049),
.A2(n_3896),
.B(n_3989),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_4072),
.B(n_3986),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_4052),
.B(n_3965),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4058),
.B(n_3965),
.Y(n_4095)
);

O2A1O1Ixp33_ASAP7_75t_L g4096 ( 
.A1(n_4048),
.A2(n_3305),
.B(n_3234),
.C(n_3261),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_4077),
.B(n_3965),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_4051),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_4075),
.B(n_3965),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_L g4100 ( 
.A(n_4069),
.B(n_619),
.Y(n_4100)
);

NOR2xp33_ASAP7_75t_L g4101 ( 
.A(n_4074),
.B(n_4068),
.Y(n_4101)
);

INVx1_ASAP7_75t_SL g4102 ( 
.A(n_4079),
.Y(n_4102)
);

INVxp67_ASAP7_75t_SL g4103 ( 
.A(n_4060),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_4064),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4070),
.B(n_3764),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_4073),
.B(n_3757),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4065),
.Y(n_4107)
);

NAND2x1p5_ASAP7_75t_L g4108 ( 
.A(n_4065),
.B(n_3764),
.Y(n_4108)
);

CKINVDCx5p33_ASAP7_75t_R g4109 ( 
.A(n_4063),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4066),
.B(n_3366),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_4066),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_L g4112 ( 
.A(n_4078),
.B(n_3543),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_4078),
.B(n_3793),
.Y(n_4113)
);

OR2x2_ASAP7_75t_L g4114 ( 
.A(n_4088),
.B(n_620),
.Y(n_4114)
);

INVx2_ASAP7_75t_L g4115 ( 
.A(n_4084),
.Y(n_4115)
);

XNOR2x1_ASAP7_75t_L g4116 ( 
.A(n_4109),
.B(n_621),
.Y(n_4116)
);

INVx2_ASAP7_75t_L g4117 ( 
.A(n_4081),
.Y(n_4117)
);

AOI22xp5_ASAP7_75t_L g4118 ( 
.A1(n_4083),
.A2(n_3329),
.B1(n_3411),
.B2(n_3550),
.Y(n_4118)
);

OAI22xp5_ASAP7_75t_L g4119 ( 
.A1(n_4089),
.A2(n_3814),
.B1(n_3357),
.B2(n_3294),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4085),
.Y(n_4120)
);

INVx1_ASAP7_75t_SL g4121 ( 
.A(n_4102),
.Y(n_4121)
);

AOI32xp33_ASAP7_75t_L g4122 ( 
.A1(n_4080),
.A2(n_4082),
.A3(n_4086),
.B1(n_4087),
.B2(n_4091),
.Y(n_4122)
);

OAI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_4092),
.A2(n_3021),
.B(n_3248),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_4104),
.B(n_3554),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4103),
.Y(n_4125)
);

NOR2xp33_ASAP7_75t_L g4126 ( 
.A(n_4101),
.B(n_621),
.Y(n_4126)
);

INVxp67_ASAP7_75t_L g4127 ( 
.A(n_4100),
.Y(n_4127)
);

INVx1_ASAP7_75t_SL g4128 ( 
.A(n_4102),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_4093),
.B(n_3336),
.Y(n_4129)
);

OAI221xp5_ASAP7_75t_SL g4130 ( 
.A1(n_4090),
.A2(n_3288),
.B1(n_3289),
.B2(n_3270),
.C(n_3330),
.Y(n_4130)
);

OR2x6_ASAP7_75t_L g4131 ( 
.A(n_4125),
.B(n_4098),
.Y(n_4131)
);

AOI22xp33_ASAP7_75t_L g4132 ( 
.A1(n_4121),
.A2(n_4097),
.B1(n_4099),
.B2(n_4106),
.Y(n_4132)
);

NAND2xp5_ASAP7_75t_L g4133 ( 
.A(n_4128),
.B(n_4107),
.Y(n_4133)
);

NOR2xp33_ASAP7_75t_R g4134 ( 
.A(n_4114),
.B(n_621),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4127),
.B(n_4111),
.Y(n_4135)
);

A2O1A1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_4122),
.A2(n_4096),
.B(n_4094),
.C(n_4095),
.Y(n_4136)
);

INVxp67_ASAP7_75t_L g4137 ( 
.A(n_4126),
.Y(n_4137)
);

A2O1A1Ixp33_ASAP7_75t_SL g4138 ( 
.A1(n_4115),
.A2(n_4112),
.B(n_4110),
.C(n_4113),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_4124),
.A2(n_4108),
.B(n_4105),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_4129),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_4123),
.B(n_4119),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_4118),
.Y(n_4142)
);

OAI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_4130),
.A2(n_3339),
.B(n_3428),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4120),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_4121),
.B(n_622),
.Y(n_4145)
);

AOI21xp5_ASAP7_75t_L g4146 ( 
.A1(n_4116),
.A2(n_3087),
.B(n_3742),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_4117),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_4121),
.B(n_657),
.Y(n_4148)
);

AOI22xp5_ASAP7_75t_L g4149 ( 
.A1(n_4120),
.A2(n_3349),
.B1(n_3801),
.B2(n_3741),
.Y(n_4149)
);

OAI221xp5_ASAP7_75t_L g4150 ( 
.A1(n_4136),
.A2(n_3203),
.B1(n_662),
.B2(n_659),
.C(n_661),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4145),
.Y(n_4151)
);

AOI22xp5_ASAP7_75t_L g4152 ( 
.A1(n_4141),
.A2(n_2928),
.B1(n_2951),
.B2(n_2912),
.Y(n_4152)
);

A2O1A1Ixp33_ASAP7_75t_L g4153 ( 
.A1(n_4137),
.A2(n_664),
.B(n_661),
.C(n_662),
.Y(n_4153)
);

AND2x4_ASAP7_75t_L g4154 ( 
.A(n_4147),
.B(n_664),
.Y(n_4154)
);

OAI22xp33_ASAP7_75t_SL g4155 ( 
.A1(n_4133),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4148),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_4131),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4131),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_L g4159 ( 
.A(n_4142),
.B(n_667),
.Y(n_4159)
);

OAI221xp5_ASAP7_75t_L g4160 ( 
.A1(n_4138),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.C(n_672),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4144),
.Y(n_4161)
);

INVxp67_ASAP7_75t_SL g4162 ( 
.A(n_4135),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4140),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4134),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4146),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_4149),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_4132),
.B(n_675),
.Y(n_4167)
);

NOR2xp33_ASAP7_75t_SL g4168 ( 
.A(n_4157),
.B(n_4139),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4164),
.Y(n_4169)
);

OAI211xp5_ASAP7_75t_L g4170 ( 
.A1(n_4158),
.A2(n_4143),
.B(n_677),
.C(n_675),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4154),
.Y(n_4171)
);

NAND2xp5_ASAP7_75t_L g4172 ( 
.A(n_4165),
.B(n_4154),
.Y(n_4172)
);

AOI221xp5_ASAP7_75t_L g4173 ( 
.A1(n_4160),
.A2(n_678),
.B1(n_676),
.B2(n_677),
.C(n_679),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4163),
.Y(n_4174)
);

NOR2xp33_ASAP7_75t_L g4175 ( 
.A(n_4167),
.B(n_681),
.Y(n_4175)
);

OAI321xp33_ASAP7_75t_L g4176 ( 
.A1(n_4166),
.A2(n_3014),
.A3(n_2970),
.B1(n_3071),
.B2(n_2992),
.C(n_2954),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4162),
.B(n_682),
.Y(n_4177)
);

OAI221xp5_ASAP7_75t_L g4178 ( 
.A1(n_4150),
.A2(n_685),
.B1(n_683),
.B2(n_684),
.C(n_686),
.Y(n_4178)
);

NAND3xp33_ASAP7_75t_L g4179 ( 
.A(n_4161),
.B(n_683),
.C(n_684),
.Y(n_4179)
);

XOR2xp5_ASAP7_75t_L g4180 ( 
.A(n_4155),
.B(n_686),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4153),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_4151),
.B(n_4156),
.Y(n_4182)
);

AND2x2_ASAP7_75t_L g4183 ( 
.A(n_4152),
.B(n_689),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4157),
.B(n_690),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4165),
.B(n_691),
.Y(n_4185)
);

NOR2x1_ASAP7_75t_L g4186 ( 
.A(n_4159),
.B(n_692),
.Y(n_4186)
);

AOI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_4168),
.A2(n_3275),
.B1(n_3071),
.B2(n_3074),
.Y(n_4187)
);

AOI221xp5_ASAP7_75t_L g4188 ( 
.A1(n_4174),
.A2(n_695),
.B1(n_693),
.B2(n_694),
.C(n_697),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4177),
.B(n_693),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_L g4190 ( 
.A(n_4184),
.B(n_694),
.Y(n_4190)
);

AOI222xp33_ASAP7_75t_L g4191 ( 
.A1(n_4181),
.A2(n_699),
.B1(n_701),
.B2(n_695),
.C1(n_698),
.C2(n_700),
.Y(n_4191)
);

AOI221xp5_ASAP7_75t_L g4192 ( 
.A1(n_4170),
.A2(n_4169),
.B1(n_4171),
.B2(n_4172),
.C(n_4176),
.Y(n_4192)
);

NOR2xp33_ASAP7_75t_L g4193 ( 
.A(n_4185),
.B(n_700),
.Y(n_4193)
);

AOI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_4180),
.A2(n_3071),
.B1(n_3074),
.B2(n_3014),
.Y(n_4194)
);

XNOR2x1_ASAP7_75t_L g4195 ( 
.A(n_4186),
.B(n_703),
.Y(n_4195)
);

INVx2_ASAP7_75t_L g4196 ( 
.A(n_4183),
.Y(n_4196)
);

AOI321xp33_ASAP7_75t_L g4197 ( 
.A1(n_4182),
.A2(n_708),
.A3(n_710),
.B1(n_704),
.B2(n_705),
.C(n_709),
.Y(n_4197)
);

AOI211xp5_ASAP7_75t_L g4198 ( 
.A1(n_4178),
.A2(n_717),
.B(n_714),
.C(n_716),
.Y(n_4198)
);

AND5x1_ASAP7_75t_L g4199 ( 
.A(n_4173),
.B(n_722),
.C(n_720),
.D(n_721),
.E(n_723),
.Y(n_4199)
);

O2A1O1Ixp33_ASAP7_75t_L g4200 ( 
.A1(n_4179),
.A2(n_723),
.B(n_721),
.C(n_722),
.Y(n_4200)
);

AOI22xp5_ASAP7_75t_L g4201 ( 
.A1(n_4175),
.A2(n_3132),
.B1(n_3164),
.B2(n_3074),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_4190),
.B(n_724),
.Y(n_4202)
);

OA22x2_ASAP7_75t_L g4203 ( 
.A1(n_4196),
.A2(n_726),
.B1(n_724),
.B2(n_725),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4189),
.Y(n_4204)
);

OAI221xp5_ASAP7_75t_L g4205 ( 
.A1(n_4197),
.A2(n_730),
.B1(n_727),
.B2(n_728),
.C(n_731),
.Y(n_4205)
);

NOR2xp33_ASAP7_75t_L g4206 ( 
.A(n_4195),
.B(n_728),
.Y(n_4206)
);

AOI32xp33_ASAP7_75t_L g4207 ( 
.A1(n_4198),
.A2(n_735),
.A3(n_733),
.B1(n_734),
.B2(n_736),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4200),
.Y(n_4208)
);

OR2x6_ASAP7_75t_L g4209 ( 
.A(n_4193),
.B(n_3164),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_4191),
.B(n_737),
.Y(n_4210)
);

BUFx12f_ASAP7_75t_L g4211 ( 
.A(n_4199),
.Y(n_4211)
);

OAI221xp5_ASAP7_75t_L g4212 ( 
.A1(n_4188),
.A2(n_4194),
.B1(n_4187),
.B2(n_4201),
.C(n_740),
.Y(n_4212)
);

AOI221xp5_ASAP7_75t_SL g4213 ( 
.A1(n_4192),
.A2(n_742),
.B1(n_738),
.B2(n_739),
.C(n_743),
.Y(n_4213)
);

AOI222xp33_ASAP7_75t_L g4214 ( 
.A1(n_4192),
.A2(n_746),
.B1(n_748),
.B2(n_742),
.C1(n_745),
.C2(n_747),
.Y(n_4214)
);

INVx2_ASAP7_75t_SL g4215 ( 
.A(n_4209),
.Y(n_4215)
);

NOR2x1_ASAP7_75t_L g4216 ( 
.A(n_4208),
.B(n_750),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4203),
.Y(n_4217)
);

NOR2xp33_ASAP7_75t_L g4218 ( 
.A(n_4210),
.B(n_751),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_4202),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_4206),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_4214),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4205),
.Y(n_4222)
);

NOR2x1_ASAP7_75t_L g4223 ( 
.A(n_4204),
.B(n_4212),
.Y(n_4223)
);

NOR2xp67_ASAP7_75t_L g4224 ( 
.A(n_4211),
.B(n_753),
.Y(n_4224)
);

AND2x2_ASAP7_75t_L g4225 ( 
.A(n_4217),
.B(n_4222),
.Y(n_4225)
);

NOR2x1_ASAP7_75t_L g4226 ( 
.A(n_4224),
.B(n_4213),
.Y(n_4226)
);

NAND3xp33_ASAP7_75t_L g4227 ( 
.A(n_4218),
.B(n_4207),
.C(n_755),
.Y(n_4227)
);

NOR3x1_ASAP7_75t_L g4228 ( 
.A(n_4221),
.B(n_756),
.C(n_757),
.Y(n_4228)
);

HB1xp67_ASAP7_75t_L g4229 ( 
.A(n_4216),
.Y(n_4229)
);

OR3x1_ASAP7_75t_L g4230 ( 
.A(n_4219),
.B(n_758),
.C(n_759),
.Y(n_4230)
);

OAI22xp33_ASAP7_75t_L g4231 ( 
.A1(n_4215),
.A2(n_3196),
.B1(n_763),
.B2(n_760),
.Y(n_4231)
);

NOR2xp67_ASAP7_75t_L g4232 ( 
.A(n_4225),
.B(n_4220),
.Y(n_4232)
);

XNOR2xp5_ASAP7_75t_L g4233 ( 
.A(n_4230),
.B(n_4223),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_4228),
.Y(n_4234)
);

AO22x2_ASAP7_75t_L g4235 ( 
.A1(n_4227),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_4235)
);

INVxp67_ASAP7_75t_SL g4236 ( 
.A(n_4232),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4235),
.Y(n_4237)
);

AOI31xp33_ASAP7_75t_L g4238 ( 
.A1(n_4233),
.A2(n_4226),
.A3(n_4229),
.B(n_4231),
.Y(n_4238)
);

INVx1_ASAP7_75t_L g4239 ( 
.A(n_4234),
.Y(n_4239)
);

INVx2_ASAP7_75t_L g4240 ( 
.A(n_4239),
.Y(n_4240)
);

OAI22xp5_ASAP7_75t_L g4241 ( 
.A1(n_4240),
.A2(n_4236),
.B1(n_4237),
.B2(n_4238),
.Y(n_4241)
);

AOI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4241),
.A2(n_768),
.B1(n_766),
.B2(n_767),
.Y(n_4242)
);

AOI22xp5_ASAP7_75t_L g4243 ( 
.A1(n_4242),
.A2(n_772),
.B1(n_769),
.B2(n_770),
.Y(n_4243)
);

NAND3xp33_ASAP7_75t_SL g4244 ( 
.A(n_4243),
.B(n_773),
.C(n_775),
.Y(n_4244)
);

INVx1_ASAP7_75t_L g4245 ( 
.A(n_4244),
.Y(n_4245)
);

OAI221xp5_ASAP7_75t_R g4246 ( 
.A1(n_4245),
.A2(n_779),
.B1(n_777),
.B2(n_778),
.C(n_780),
.Y(n_4246)
);

AOI211xp5_ASAP7_75t_L g4247 ( 
.A1(n_4246),
.A2(n_784),
.B(n_780),
.C(n_783),
.Y(n_4247)
);


endmodule