module fake_jpeg_16980_n_175 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_SL g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_74),
.A2(n_65),
.B1(n_48),
.B2(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_89),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_65),
.B1(n_48),
.B2(n_61),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_51),
.B1(n_62),
.B2(n_67),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_49),
.B1(n_66),
.B2(n_64),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_1),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_49),
.Y(n_106)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_104),
.Y(n_127)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_106),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_2),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_124)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_113),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_56),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_80),
.A2(n_60),
.B1(n_57),
.B2(n_55),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_2),
.B(n_4),
.C(n_5),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_110),
.B(n_98),
.C(n_105),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_20),
.B1(n_46),
.B2(n_45),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_134),
.B1(n_112),
.B2(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_52),
.C(n_19),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_SL g140 ( 
.A(n_132),
.B(n_5),
.C(n_6),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_99),
.A2(n_18),
.B1(n_42),
.B2(n_41),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_97),
.B1(n_101),
.B2(n_102),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_135),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_4),
.Y(n_137)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_24),
.B1(n_43),
.B2(n_40),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_128),
.C(n_134),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_132),
.B(n_122),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_139),
.B(n_130),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_148),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_129),
.C(n_133),
.Y(n_157)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_151),
.B1(n_133),
.B2(n_7),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_144),
.B1(n_125),
.B2(n_123),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_107),
.C(n_131),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_155),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_156),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_16),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_154),
.B(n_149),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_129),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_162),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_160),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_15),
.C(n_35),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_12),
.Y(n_167)
);

NOR3x1_ASAP7_75t_SL g168 ( 
.A(n_167),
.B(n_17),
.C(n_34),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_168),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_169),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_39),
.C(n_33),
.Y(n_172)
);

OAI321xp33_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_31),
.A3(n_27),
.B1(n_25),
.B2(n_9),
.C(n_10),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_6),
.C(n_7),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_174),
.B(n_8),
.Y(n_175)
);


endmodule