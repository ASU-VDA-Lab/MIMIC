module fake_jpeg_11590_n_134 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_10;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_30),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_1),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_1),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_28),
.A2(n_20),
.B1(n_18),
.B2(n_22),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_63),
.B1(n_74),
.B2(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_4),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_22),
.C(n_23),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_68),
.C(n_61),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_31),
.A2(n_32),
.B1(n_48),
.B2(n_50),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_59),
.A2(n_56),
.B1(n_70),
.B2(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_63)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_24),
.B(n_5),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_73),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_28),
.A2(n_25),
.B1(n_16),
.B2(n_24),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_4),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_5),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_90),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_63),
.B(n_64),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_91),
.B(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_88),
.A2(n_66),
.B1(n_75),
.B2(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_56),
.B1(n_70),
.B2(n_55),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_55),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_61),
.C(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_65),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_90),
.B(n_85),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_101),
.C(n_92),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_108),
.B(n_110),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_84),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_86),
.B1(n_91),
.B2(n_93),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_105),
.B1(n_100),
.B2(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_114),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_79),
.Y(n_114)
);

AOI221xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_120),
.B1(n_109),
.B2(n_119),
.C(n_116),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_119),
.C(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_95),
.B1(n_98),
.B2(n_106),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_122),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_110),
.C(n_102),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_103),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_117),
.C(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_97),
.B(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g131 ( 
.A(n_128),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_130),
.A3(n_127),
.B1(n_126),
.B2(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_94),
.Y(n_134)
);


endmodule