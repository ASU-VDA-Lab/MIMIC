module real_jpeg_7231_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_0),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_0),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_0),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_0),
.B(n_82),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_0),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_0),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_0),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_1),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_1),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_1),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_1),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_1),
.B(n_359),
.Y(n_358)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_3),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_3),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_3),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_3),
.B(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_3),
.B(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_3),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B1(n_22),
.B2(n_24),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_5),
.Y(n_93)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_5),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g446 ( 
.A(n_5),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_5),
.Y(n_483)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_5),
.Y(n_510)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_6),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_7),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_7),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_7),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_7),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_7),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_7),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_7),
.B(n_394),
.Y(n_393)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_9),
.Y(n_191)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_9),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_10),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_10),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_10),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_10),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_10),
.B(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_11),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_11),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_11),
.B(n_39),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_11),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_11),
.B(n_270),
.Y(n_315)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_14),
.Y(n_98)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_14),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_14),
.Y(n_303)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_15),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_15),
.Y(n_379)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_15),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_16),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_16),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_16),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_16),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_16),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_16),
.B(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_16),
.B(n_509),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_17),
.B(n_142),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_17),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_17),
.B(n_396),
.Y(n_395)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_521),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_499),
.B(n_520),
.Y(n_25)
);

AOI21x1_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_437),
.B(n_496),
.Y(n_26)
);

AO21x2_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_280),
.B(n_317),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_237),
.B(n_279),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_210),
.B(n_236),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_30),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_166),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_31),
.B(n_166),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_112),
.C(n_150),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_32),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_77),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_33),
.B(n_78),
.C(n_95),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_50),
.C(n_66),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_34),
.B(n_232),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_34),
.Y(n_535)
);

FAx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_42),
.CI(n_46),
.CON(n_34),
.SN(n_34)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_35),
.B(n_42),
.C(n_46),
.Y(n_165)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_37),
.B(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_39),
.Y(n_369)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_40),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_48),
.Y(n_149)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_48),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_49),
.Y(n_139)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_49),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_49),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_50),
.A2(n_66),
.B1(n_67),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_50),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.C(n_63),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_51),
.A2(n_63),
.B1(n_188),
.B2(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_51),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_51),
.A2(n_219),
.B1(n_229),
.B2(n_260),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_51),
.A2(n_114),
.B1(n_115),
.B2(n_219),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_51),
.B(n_229),
.C(n_286),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

OR2x2_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_81),
.Y(n_80)
);

OR2x2_ASAP7_75t_SL g174 ( 
.A(n_52),
.B(n_175),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_52),
.B(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_55),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_56),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_56),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_57),
.B(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_62),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_63),
.A2(n_188),
.B1(n_189),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_63),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_63),
.B(n_189),
.C(n_194),
.Y(n_243)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_72),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_230)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_71),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_71),
.Y(n_388)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g463 ( 
.A(n_76),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_95),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_79),
.A2(n_80),
.B1(n_114),
.B2(n_115),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_79),
.B(n_115),
.C(n_481),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_79),
.A2(n_80),
.B1(n_173),
.B2(n_174),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_79),
.B(n_174),
.C(n_300),
.Y(n_527)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_80),
.B(n_87),
.C(n_92),
.Y(n_201)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_83),
.Y(n_228)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_84),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_84),
.Y(n_348)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_87),
.A2(n_94),
.B1(n_135),
.B2(n_136),
.Y(n_353)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_97),
.B(n_99),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_96),
.B(n_105),
.C(n_107),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_98),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_103),
.B(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_108),
.B(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_108),
.B(n_351),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_108),
.B(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_112),
.B(n_150),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_130),
.C(n_132),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_113),
.A2(n_130),
.B1(n_131),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_129),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_119),
.C(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_115),
.B(n_219),
.C(n_460),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_117),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_117),
.Y(n_335)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_117),
.Y(n_352)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_124),
.B1(n_125),
.B2(n_128),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_124),
.A2(n_125),
.B1(n_245),
.B2(n_251),
.Y(n_244)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_125),
.B(n_246),
.C(n_247),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_132),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_140),
.C(n_146),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_133),
.A2(n_134),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_147),
.Y(n_425)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_145),
.Y(n_297)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_165),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_153),
.C(n_165),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_157),
.C(n_160),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_155),
.A2(n_295),
.B1(n_298),
.B2(n_299),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_155),
.Y(n_299)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_164),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_167),
.B(n_169),
.C(n_209),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_196),
.B1(n_208),
.B2(n_209),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_185),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_171),
.B(n_172),
.C(n_185),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_184),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_173),
.A2(n_174),
.B1(n_255),
.B2(n_256),
.Y(n_529)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_174),
.B(n_276),
.C(n_277),
.Y(n_275)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_182),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_193),
.B2(n_194),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_189),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_189),
.A2(n_192),
.B1(n_229),
.B2(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_189),
.B(n_229),
.C(n_256),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_189),
.A2(n_192),
.B1(n_345),
.B2(n_346),
.Y(n_363)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_192),
.B(n_345),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_193),
.A2(n_194),
.B1(n_450),
.B2(n_454),
.Y(n_449)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_194),
.B(n_444),
.C(n_450),
.Y(n_476)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_196),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_197),
.B(n_199),
.C(n_200),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_205),
.C(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_234),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_211),
.B(n_234),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.C(n_231),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_212),
.A2(n_213),
.B1(n_430),
.B2(n_431),
.Y(n_429)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_216),
.B(n_231),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_230),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_217),
.B(n_417),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_220),
.B(n_230),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.C(n_229),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_221),
.A2(n_222),
.B1(n_226),
.B2(n_227),
.Y(n_342)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_229),
.A2(n_260),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_238),
.B(n_280),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g279 ( 
.A(n_239),
.B(n_240),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_240),
.B(n_281),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_240),
.B(n_281),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_262),
.CI(n_278),
.CON(n_240),
.SN(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_254),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_252),
.B2(n_253),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_243),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_243),
.B(n_253),
.C(n_254),
.Y(n_307)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_250),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_261),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_259),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_265),
.C(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_275),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_273),
.C(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_274),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_271),
.A2(n_274),
.B1(n_471),
.B2(n_472),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_271),
.B(n_471),
.C(n_476),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_274),
.B(n_312),
.C(n_315),
.Y(n_456)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_282),
.B(n_284),
.C(n_305),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_305),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_285),
.B(n_291),
.C(n_292),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

INVx6_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_300),
.B2(n_304),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_295),
.B(n_299),
.C(n_300),
.Y(n_465)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_300),
.A2(n_304),
.B1(n_516),
.B2(n_517),
.Y(n_515)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_303),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_316),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_306),
.B(n_309),
.C(n_311),
.Y(n_492)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_308),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

OAI31xp33_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_433),
.A3(n_434),
.B(n_436),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_427),
.B(n_432),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_412),
.B(n_426),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_364),
.B(n_411),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_354),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_322),
.B(n_354),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_343),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_340),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_340),
.C(n_343),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_331),
.C(n_336),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_326),
.B1(n_331),
.B2(n_332),
.Y(n_356)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx8_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_336),
.B(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_421),
.C(n_422),
.Y(n_420)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_353),
.Y(n_349)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.C(n_363),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_357),
.A2(n_363),
.B1(n_403),
.B2(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_361),
.Y(n_402)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_363),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_405),
.B(n_410),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_390),
.B(n_404),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_374),
.B(n_389),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_385),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_385),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_376),
.A2(n_380),
.B(n_384),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_380),
.Y(n_384)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_384),
.A2(n_392),
.B1(n_398),
.B2(n_399),
.Y(n_391)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx8_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_400),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_392),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_395),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_393),
.A2(n_395),
.B(n_398),
.Y(n_406)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_402),
.B(n_403),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_406),
.B(n_407),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_414),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_416),
.B1(n_418),
.B2(n_419),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_420),
.C(n_423),
.Y(n_428)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_423),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_429),
.Y(n_432)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_430),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_493),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_438),
.A2(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_485),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_439),
.B(n_485),
.Y(n_498)
);

BUFx24_ASAP7_75t_SL g537 ( 
.A(n_439),
.Y(n_537)
);

FAx1_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_457),
.CI(n_467),
.CON(n_439),
.SN(n_439)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_440),
.B(n_457),
.C(n_467),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.C(n_456),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_441),
.A2(n_442),
.B1(n_487),
.B2(n_488),
.Y(n_486)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_443),
.B(n_456),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_448),
.B1(n_449),
.B2(n_455),
.Y(n_443)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_444),
.A2(n_455),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

INVx8_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_450),
.Y(n_454)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_465),
.C(n_466),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_459),
.B1(n_490),
.B2(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_464),
.Y(n_459)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx6_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_466),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_469),
.B1(n_477),
.B2(n_484),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_468),
.B(n_478),
.C(n_479),
.Y(n_518)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_476),
.Y(n_469)
);

CKINVDCx14_ASAP7_75t_R g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx8_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_477),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.C(n_492),
.Y(n_485)
);

FAx1_ASAP7_75t_SL g495 ( 
.A(n_486),
.B(n_489),
.CI(n_492),
.CON(n_495),
.SN(n_495)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_487),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_495),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g538 ( 
.A(n_495),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_519),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_500),
.B(n_519),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_518),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_504),
.B2(n_505),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_503),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_504),
.C(n_518),
.Y(n_533)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_514),
.B2(n_515),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_508),
.Y(n_512)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_511),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_512),
.C(n_514),
.Y(n_525)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g516 ( 
.A(n_517),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_534),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_533),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_524),
.B(n_533),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_531),
.B2(n_532),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_527),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_528),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_529),
.Y(n_530)
);


endmodule