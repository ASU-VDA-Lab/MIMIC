module fake_jpeg_3481_n_680 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_12),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_1),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_62),
.Y(n_140)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx11_ASAP7_75t_SL g180 ( 
.A(n_64),
.Y(n_180)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_65),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_67),
.B(n_79),
.Y(n_151)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_68),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_70),
.B(n_75),
.Y(n_184)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_71),
.Y(n_197)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g189 ( 
.A(n_74),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_16),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_26),
.B(n_0),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_81),
.B(n_110),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_82),
.B(n_90),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_85),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_87),
.Y(n_148)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_91),
.Y(n_191)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_94),
.B(n_95),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_21),
.Y(n_97)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_98),
.Y(n_219)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_99),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_24),
.Y(n_101)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_103),
.B(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_106),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_48),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_48),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_109),
.B(n_111),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_15),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_23),
.B(n_2),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_53),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_112),
.B(n_115),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_53),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_38),
.Y(n_117)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

INVx11_ASAP7_75t_SL g118 ( 
.A(n_47),
.Y(n_118)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_22),
.Y(n_119)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_28),
.B(n_2),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_121),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g220 ( 
.A(n_122),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_36),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_124),
.B(n_33),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_38),
.Y(n_126)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_126),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_127),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_36),
.Y(n_128)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_22),
.Y(n_130)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g131 ( 
.A(n_38),
.Y(n_131)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_98),
.A2(n_27),
.B1(n_58),
.B2(n_54),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_134),
.A2(n_102),
.B1(n_78),
.B2(n_80),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_136),
.B(n_167),
.Y(n_238)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_22),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_142),
.B(n_154),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_58),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_144),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_66),
.A2(n_27),
.B1(n_22),
.B2(n_45),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_157),
.B1(n_177),
.B2(n_54),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_68),
.B(n_59),
.C(n_30),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_27),
.B1(n_58),
.B2(n_54),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_158),
.Y(n_293)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_69),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_159),
.Y(n_237)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_161),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_65),
.Y(n_167)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_172),
.Y(n_273)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_175),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_86),
.A2(n_37),
.B1(n_59),
.B2(n_52),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_101),
.B(n_52),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_178),
.B(n_39),
.Y(n_254)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_89),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_91),
.Y(n_196)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_88),
.Y(n_198)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_92),
.Y(n_207)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_208),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_64),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_108),
.Y(n_214)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_214),
.Y(n_282)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_126),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_218),
.Y(n_234)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_85),
.Y(n_221)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_87),
.B(n_45),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_84),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_226),
.A2(n_240),
.B1(n_244),
.B2(n_277),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_228),
.B(n_233),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_37),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_231),
.B(n_247),
.Y(n_352)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_217),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_232),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_35),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_35),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_236),
.B(n_245),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_142),
.A2(n_123),
.B1(n_99),
.B2(n_77),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_239),
.A2(n_243),
.B1(n_265),
.B2(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_185),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_241),
.Y(n_318)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_242),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_206),
.A2(n_30),
.B1(n_34),
.B2(n_33),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_102),
.B1(n_34),
.B2(n_50),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_32),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_151),
.B(n_32),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_248),
.B(n_254),
.Y(n_310)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_148),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_249),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_157),
.A2(n_31),
.B1(n_26),
.B2(n_39),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_250),
.A2(n_286),
.B1(n_179),
.B2(n_199),
.Y(n_351)
);

BUFx12_ASAP7_75t_L g252 ( 
.A(n_195),
.Y(n_252)
);

BUFx8_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_132),
.Y(n_253)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

BUFx12_ASAP7_75t_L g255 ( 
.A(n_216),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_255),
.Y(n_348)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_162),
.Y(n_256)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

OA22x2_ASAP7_75t_SL g257 ( 
.A1(n_144),
.A2(n_62),
.B1(n_93),
.B2(n_122),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g341 ( 
.A1(n_257),
.A2(n_156),
.B1(n_194),
.B2(n_135),
.Y(n_341)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

BUFx12f_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_260),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_151),
.B(n_60),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_262),
.B(n_264),
.Y(n_363)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_60),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_215),
.A2(n_31),
.B1(n_49),
.B2(n_50),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_215),
.B(n_49),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_178),
.B(n_122),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_267),
.Y(n_345)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_173),
.Y(n_268)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_164),
.B(n_2),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_169),
.B(n_3),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_270),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_188),
.A2(n_47),
.B1(n_113),
.B2(n_125),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_170),
.B(n_3),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_182),
.B(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_6),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_139),
.A2(n_47),
.B1(n_129),
.B2(n_125),
.Y(n_277)
);

INVx11_ASAP7_75t_L g279 ( 
.A(n_139),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_279),
.Y(n_355)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_197),
.Y(n_280)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_280),
.Y(n_325)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_202),
.Y(n_281)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_212),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_217),
.Y(n_285)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_285),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_134),
.A2(n_131),
.B1(n_96),
.B2(n_46),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_210),
.A2(n_131),
.B1(n_96),
.B2(n_46),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_288),
.A2(n_298),
.B1(n_189),
.B2(n_183),
.Y(n_316)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_141),
.B(n_5),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_290),
.A2(n_301),
.B1(n_223),
.B2(n_189),
.Y(n_338)
);

BUFx12f_ASAP7_75t_L g291 ( 
.A(n_166),
.Y(n_291)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_160),
.B(n_5),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_295),
.Y(n_342)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_193),
.Y(n_296)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_174),
.Y(n_297)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_145),
.A2(n_46),
.B1(n_6),
.B2(n_7),
.Y(n_298)
);

INVx11_ASAP7_75t_L g299 ( 
.A(n_174),
.Y(n_299)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_212),
.Y(n_300)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_146),
.B(n_5),
.Y(n_301)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_204),
.B(n_46),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_183),
.C(n_143),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_205),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_305),
.Y(n_373)
);

AOI22x1_ASAP7_75t_SL g307 ( 
.A1(n_278),
.A2(n_153),
.B1(n_140),
.B2(n_176),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_307),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_312),
.B(n_7),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_143),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_314),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_316),
.A2(n_321),
.B1(n_328),
.B2(n_350),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_239),
.A2(n_194),
.B1(n_135),
.B2(n_156),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_240),
.A2(n_155),
.B1(n_201),
.B2(n_200),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_250),
.A2(n_163),
.B1(n_201),
.B2(n_200),
.Y(n_333)
);

OA22x2_ASAP7_75t_L g375 ( 
.A1(n_333),
.A2(n_351),
.B1(n_362),
.B2(n_242),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_292),
.B(n_302),
.C(n_229),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_249),
.C(n_280),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_338),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_292),
.A2(n_133),
.B(n_220),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_339),
.A2(n_341),
.B(n_234),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_238),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_349),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_224),
.B(n_163),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_346),
.B(n_272),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_225),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_244),
.A2(n_191),
.B1(n_199),
.B2(n_152),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_235),
.Y(n_353)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_227),
.Y(n_354)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_257),
.A2(n_191),
.B1(n_152),
.B2(n_150),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_237),
.B1(n_275),
.B2(n_282),
.Y(n_386)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_251),
.Y(n_358)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_261),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_294),
.Y(n_395)
);

NAND2xp67_ASAP7_75t_SL g361 ( 
.A(n_257),
.B(n_133),
.Y(n_361)
);

NOR3xp33_ASAP7_75t_SL g403 ( 
.A(n_361),
.B(n_252),
.C(n_133),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_286),
.A2(n_237),
.B1(n_261),
.B2(n_275),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_335),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_365),
.B(n_372),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_351),
.A2(n_277),
.B1(n_150),
.B2(n_147),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_366),
.A2(n_392),
.B1(n_314),
.B2(n_355),
.Y(n_416)
);

INVx6_ASAP7_75t_L g367 ( 
.A(n_360),
.Y(n_367)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_367),
.Y(n_431)
);

BUFx12_ASAP7_75t_L g370 ( 
.A(n_335),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_335),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_390),
.C(n_396),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_375),
.B(n_403),
.Y(n_424)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_348),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_379),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_315),
.B(n_318),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_388),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_336),
.B(n_281),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_381),
.B(n_337),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_383),
.B(n_393),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_330),
.Y(n_384)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_386),
.A2(n_387),
.B1(n_409),
.B2(n_412),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_303),
.A2(n_345),
.B1(n_341),
.B2(n_305),
.Y(n_387)
);

OA22x2_ASAP7_75t_SL g389 ( 
.A1(n_341),
.A2(n_282),
.B1(n_285),
.B2(n_232),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_389),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_268),
.C(n_234),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_306),
.A2(n_293),
.B(n_246),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_391),
.A2(n_394),
.B(n_410),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_361),
.A2(n_138),
.B1(n_147),
.B2(n_230),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_346),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_314),
.A2(n_293),
.B(n_246),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_395),
.B(n_398),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_332),
.B(n_294),
.C(n_259),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_315),
.B(n_259),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_401),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_400),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_318),
.B(n_319),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_317),
.B(n_323),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_402),
.B(n_404),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_311),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_317),
.B(n_273),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_405),
.B(n_406),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_320),
.B(n_230),
.Y(n_406)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_309),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_407),
.B(n_408),
.Y(n_446)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_309),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_356),
.Y(n_409)
);

INVx13_ASAP7_75t_L g410 ( 
.A(n_348),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_319),
.B(n_273),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_411),
.A2(n_365),
.B1(n_372),
.B2(n_385),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_334),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_310),
.B(n_272),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_413),
.A2(n_352),
.B1(n_363),
.B2(n_347),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_305),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_414),
.B(n_419),
.C(n_421),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_416),
.A2(n_418),
.B1(n_439),
.B2(n_440),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_385),
.A2(n_338),
.B(n_323),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g476 ( 
.A1(n_417),
.A2(n_441),
.B(n_452),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_387),
.A2(n_341),
.B1(n_326),
.B2(n_308),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_378),
.B(n_304),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_304),
.C(n_308),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_393),
.A2(n_326),
.B1(n_342),
.B2(n_312),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_427),
.A2(n_429),
.B1(n_392),
.B2(n_366),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_382),
.A2(n_307),
.B1(n_334),
.B2(n_287),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_432),
.B(n_453),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_354),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_442),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_388),
.A2(n_344),
.B(n_340),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_437),
.A2(n_412),
.B(n_389),
.Y(n_473)
);

AO21x1_ASAP7_75t_L g472 ( 
.A1(n_438),
.A2(n_394),
.B(n_403),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_376),
.A2(n_364),
.B1(n_347),
.B2(n_327),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_376),
.A2(n_364),
.B1(n_325),
.B2(n_327),
.Y(n_440)
);

AND2x2_ASAP7_75t_SL g441 ( 
.A(n_373),
.B(n_311),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_390),
.B(n_337),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_444),
.B(n_447),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_382),
.A2(n_325),
.B1(n_340),
.B2(n_287),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_384),
.B1(n_397),
.B2(n_367),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_373),
.B(n_353),
.Y(n_447)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_358),
.C(n_330),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_451),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_396),
.B(n_313),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_377),
.A2(n_330),
.B(n_344),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_377),
.B(n_313),
.C(n_322),
.Y(n_453)
);

BUFx12_ASAP7_75t_L g455 ( 
.A(n_425),
.Y(n_455)
);

INVx11_ASAP7_75t_L g502 ( 
.A(n_455),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_434),
.B(n_380),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_456),
.B(n_458),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_427),
.B(n_413),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_421),
.B(n_368),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_461),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_430),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_463),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_406),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_324),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_462),
.B(n_469),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_446),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_483),
.B1(n_486),
.B2(n_491),
.Y(n_497)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_465),
.Y(n_499)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_422),
.A2(n_386),
.B1(n_391),
.B2(n_389),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_467),
.A2(n_475),
.B1(n_429),
.B2(n_424),
.Y(n_494)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_468),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_324),
.Y(n_469)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_471),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_472),
.A2(n_473),
.B(n_437),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_474),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_422),
.A2(n_389),
.B1(n_399),
.B2(n_375),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_448),
.B(n_383),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_479),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_454),
.B(n_322),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_439),
.Y(n_480)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_480),
.Y(n_518)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_440),
.Y(n_481)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_420),
.B(n_369),
.Y(n_482)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_418),
.A2(n_375),
.B1(n_371),
.B2(n_369),
.Y(n_483)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_485),
.B(n_487),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_419),
.B(n_371),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_446),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_397),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_492),
.Y(n_514)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_453),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_494),
.A2(n_487),
.B1(n_476),
.B2(n_457),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_473),
.B(n_424),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_495),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_498),
.A2(n_501),
.B(n_526),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_478),
.B(n_415),
.C(n_451),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_500),
.B(n_509),
.Y(n_547)
);

OAI32xp33_ASAP7_75t_L g501 ( 
.A1(n_482),
.A2(n_426),
.A3(n_424),
.B1(n_447),
.B2(n_442),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_456),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_508),
.B(n_528),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_478),
.B(n_433),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_415),
.C(n_444),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_513),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_460),
.A2(n_445),
.B1(n_416),
.B2(n_417),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_512),
.A2(n_515),
.B1(n_367),
.B2(n_331),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_414),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_467),
.A2(n_426),
.B1(n_438),
.B2(n_423),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_464),
.A2(n_423),
.B1(n_441),
.B2(n_452),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_516),
.A2(n_520),
.B1(n_527),
.B2(n_476),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_446),
.Y(n_517)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_517),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_483),
.A2(n_441),
.B1(n_375),
.B2(n_408),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_435),
.C(n_384),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_523),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_488),
.B(n_435),
.C(n_410),
.Y(n_523)
);

AO22x1_ASAP7_75t_L g526 ( 
.A1(n_475),
.A2(n_408),
.B1(n_407),
.B2(n_400),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_480),
.A2(n_490),
.B1(n_481),
.B2(n_463),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_468),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_529),
.A2(n_546),
.B1(n_526),
.B2(n_518),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_503),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_531),
.B(n_539),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g533 ( 
.A(n_525),
.Y(n_533)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_533),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_535),
.B1(n_542),
.B2(n_543),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_497),
.A2(n_470),
.B1(n_488),
.B2(n_465),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_502),
.Y(n_536)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_536),
.Y(n_568)
);

AOI21xp33_ASAP7_75t_L g537 ( 
.A1(n_514),
.A2(n_477),
.B(n_472),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_537),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_494),
.A2(n_466),
.B1(n_485),
.B2(n_471),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_538),
.A2(n_550),
.B1(n_552),
.B2(n_560),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_503),
.A2(n_489),
.B(n_455),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_513),
.B(n_489),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_540),
.B(n_554),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g541 ( 
.A(n_504),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_555),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_516),
.A2(n_400),
.B1(n_455),
.B2(n_407),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_527),
.A2(n_455),
.B1(n_329),
.B2(n_331),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_544),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_SL g548 ( 
.A1(n_520),
.A2(n_279),
.B1(n_329),
.B2(n_291),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_548),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_515),
.A2(n_138),
.B1(n_291),
.B2(n_253),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g551 ( 
.A(n_501),
.B(n_370),
.CI(n_410),
.CON(n_551),
.SN(n_551)
);

OR2x2_ASAP7_75t_L g577 ( 
.A(n_551),
.B(n_523),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_522),
.A2(n_260),
.B1(n_253),
.B2(n_297),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_507),
.Y(n_553)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_553),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_495),
.A2(n_370),
.B1(n_379),
.B2(n_260),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_514),
.B(n_252),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_556),
.B(n_511),
.Y(n_585)
);

CKINVDCx16_ASAP7_75t_R g557 ( 
.A(n_493),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_557),
.B(n_559),
.Y(n_588)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_496),
.B(n_370),
.C(n_379),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_522),
.A2(n_299),
.B1(n_203),
.B2(n_11),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_547),
.B(n_500),
.C(n_521),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_564),
.B(n_556),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_545),
.B(n_505),
.Y(n_566)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_566),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_541),
.B(n_505),
.Y(n_569)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_569),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_530),
.B(n_506),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_570),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_549),
.A2(n_498),
.B(n_495),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_571),
.A2(n_551),
.B(n_550),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_506),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_572),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_519),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_575),
.B(n_578),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g603 ( 
.A(n_577),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_534),
.B(n_519),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_509),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_580),
.B(n_584),
.Y(n_601)
);

INVx13_ASAP7_75t_L g581 ( 
.A(n_536),
.Y(n_581)
);

INVx13_ASAP7_75t_L g607 ( 
.A(n_581),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_582),
.A2(n_542),
.B1(n_532),
.B2(n_554),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_529),
.Y(n_584)
);

MAJx2_ASAP7_75t_L g594 ( 
.A(n_585),
.B(n_587),
.C(n_540),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_524),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_571),
.A2(n_573),
.B(n_577),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_589),
.A2(n_595),
.B(n_602),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_535),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_590),
.B(n_591),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_564),
.B(n_561),
.C(n_558),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_592),
.A2(n_586),
.B1(n_569),
.B2(n_583),
.Y(n_623)
);

XNOR2x1_ASAP7_75t_L g628 ( 
.A(n_594),
.B(n_576),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_588),
.A2(n_532),
.B(n_551),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_563),
.B(n_584),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g614 ( 
.A(n_597),
.B(n_594),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_598),
.B(n_599),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_565),
.B(n_552),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_510),
.C(n_499),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_604),
.B(n_609),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_510),
.Y(n_608)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_608),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_587),
.B(n_499),
.C(n_560),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_585),
.B(n_563),
.C(n_578),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_610),
.Y(n_622)
);

A2O1A1O1Ixp25_ASAP7_75t_L g611 ( 
.A1(n_566),
.A2(n_526),
.B(n_502),
.C(n_255),
.D(n_12),
.Y(n_611)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_611),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_595),
.A2(n_582),
.B1(n_579),
.B2(n_575),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g633 ( 
.A1(n_612),
.A2(n_592),
.B1(n_593),
.B2(n_600),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_603),
.B(n_562),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_613),
.B(n_619),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_614),
.B(n_623),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_603),
.B(n_568),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_589),
.B(n_568),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_620),
.B(n_621),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_601),
.B(n_574),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_596),
.A2(n_579),
.B1(n_572),
.B2(n_586),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_624),
.B(n_625),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_601),
.B(n_570),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_606),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_626),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_593),
.A2(n_576),
.B1(n_581),
.B2(n_11),
.Y(n_627)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_627),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_628),
.B(n_597),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_622),
.B(n_591),
.C(n_604),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_634),
.Y(n_647)
);

MAJx2_ASAP7_75t_L g652 ( 
.A(n_633),
.B(n_637),
.C(n_646),
.Y(n_652)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_616),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_616),
.A2(n_606),
.B(n_605),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_623),
.A2(n_605),
.B(n_602),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_641),
.A2(n_642),
.B1(n_629),
.B2(n_609),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_612),
.A2(n_596),
.B(n_600),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_627),
.Y(n_643)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_643),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_618),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_644),
.B(n_645),
.Y(n_648)
);

CKINVDCx16_ASAP7_75t_R g645 ( 
.A(n_617),
.Y(n_645)
);

AOI21xp33_ASAP7_75t_L g649 ( 
.A1(n_638),
.A2(n_615),
.B(n_630),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_SL g664 ( 
.A1(n_649),
.A2(n_656),
.B(n_636),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_650),
.B(n_639),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_632),
.B(n_625),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_651),
.B(n_653),
.Y(n_660)
);

MAJx2_ASAP7_75t_L g653 ( 
.A(n_633),
.B(n_614),
.C(n_628),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_631),
.B(n_621),
.C(n_610),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_655),
.B(n_657),
.Y(n_661)
);

NOR2x1_ASAP7_75t_L g656 ( 
.A(n_637),
.B(n_607),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_607),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_635),
.B(n_611),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_658),
.B(n_639),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_659),
.B(n_662),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_648),
.A2(n_642),
.B1(n_641),
.B2(n_643),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_663),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_664),
.B(n_666),
.Y(n_668)
);

AO21x1_ASAP7_75t_L g665 ( 
.A1(n_647),
.A2(n_654),
.B(n_656),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_SL g670 ( 
.A1(n_665),
.A2(n_660),
.B(n_661),
.C(n_652),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_652),
.B(n_646),
.C(n_636),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_670),
.A2(n_9),
.B(n_10),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_SL g671 ( 
.A1(n_665),
.A2(n_653),
.B(n_255),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_671),
.B(n_666),
.Y(n_673)
);

XNOR2xp5_ASAP7_75t_L g672 ( 
.A(n_667),
.B(n_659),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_672),
.B(n_673),
.C(n_674),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g676 ( 
.A(n_672),
.B(n_669),
.C(n_668),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_676),
.B(n_46),
.C(n_13),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_677),
.A2(n_675),
.B(n_13),
.Y(n_678)
);

OAI221xp5_ASAP7_75t_SL g679 ( 
.A1(n_678),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_679)
);

AO21x1_ASAP7_75t_L g680 ( 
.A1(n_679),
.A2(n_14),
.B(n_15),
.Y(n_680)
);


endmodule