module fake_netlist_6_934_n_197 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_197);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_197;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_145;
wire n_92;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_66;
wire n_85;
wire n_130;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_196;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVxp33_ASAP7_75t_SL g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

CKINVDCx5p33_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_R g67 ( 
.A(n_52),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_R g68 ( 
.A(n_52),
.B(n_0),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_32),
.B(n_1),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_R g75 ( 
.A(n_41),
.B(n_3),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_44),
.B(n_4),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_44),
.B1(n_49),
.B2(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_47),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_49),
.Y(n_83)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_45),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_42),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_53),
.B1(n_43),
.B2(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_48),
.B1(n_51),
.B2(n_34),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_80),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_59),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_59),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_66),
.B(n_70),
.C(n_69),
.Y(n_97)
);

O2A1O1Ixp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_59),
.B(n_63),
.C(n_70),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AO21x2_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_75),
.B(n_72),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_59),
.B(n_63),
.C(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_79),
.B(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_84),
.B1(n_91),
.B2(n_77),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_83),
.Y(n_111)
);

OAI221xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_84),
.B1(n_69),
.B2(n_73),
.C(n_93),
.Y(n_112)
);

OAI21x1_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_70),
.B(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_77),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_100),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_110),
.A2(n_77),
.B1(n_87),
.B2(n_100),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_77),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_112),
.B1(n_84),
.B2(n_87),
.Y(n_121)
);

AO21x2_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_113),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_116),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_118),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_102),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_116),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_120),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_121),
.B(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_132),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_122),
.Y(n_140)
);

NAND2x1p5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_115),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_143),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_130),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_130),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_129),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_134),
.B1(n_120),
.B2(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_148),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_122),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

AOI211xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_72),
.B(n_75),
.C(n_68),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_151),
.Y(n_165)
);

OAI211xp5_ASAP7_75t_SL g166 ( 
.A1(n_157),
.A2(n_57),
.B(n_64),
.C(n_92),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_68),
.B1(n_87),
.B2(n_73),
.C(n_63),
.Y(n_167)
);

NAND3x1_ASAP7_75t_SL g168 ( 
.A(n_160),
.B(n_5),
.C(n_8),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_87),
.B1(n_126),
.B2(n_115),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_162),
.B(n_126),
.Y(n_170)
);

OAI211xp5_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_159),
.B(n_158),
.C(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_64),
.B1(n_57),
.B2(n_59),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_92),
.C(n_81),
.Y(n_173)
);

AOI222xp33_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_63),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_9),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_63),
.B1(n_11),
.B2(n_12),
.C(n_9),
.Y(n_175)
);

NAND4xp75_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_98),
.C(n_89),
.D(n_95),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.Y(n_177)
);

AOI221xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_113),
.B1(n_90),
.B2(n_89),
.C(n_96),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_107),
.B1(n_90),
.B2(n_96),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_15),
.B(n_17),
.C(n_24),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

AND3x1_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_26),
.C(n_103),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_R g184 ( 
.A(n_177),
.B(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_182),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_99),
.B(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_183),
.B(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_184),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_189),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_191),
.B1(n_186),
.B2(n_185),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_193),
.B1(n_188),
.B2(n_192),
.Y(n_196)
);

NAND3xp33_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_187),
.C(n_99),
.Y(n_197)
);


endmodule