module fake_aes_742_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_30;
wire n_16;
wire n_26;
wire n_25;
wire n_33;
wire n_13;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
BUFx6f_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_2), .Y(n_12) );
NOR2xp67_ASAP7_75t_L g13 ( .A(n_7), .B(n_1), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_5), .B(n_4), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_2), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
OR2x6_ASAP7_75t_L g20 ( .A(n_14), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_16), .B(n_3), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_11), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_12), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_16), .A2(n_3), .B1(n_5), .B2(n_6), .Y(n_24) );
AOI22xp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_11), .B1(n_17), .B2(n_15), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_20), .A2(n_11), .B1(n_18), .B2(n_15), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_19), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_26), .B(n_20), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND2xp5_ASAP7_75t_SL g31 ( .A(n_29), .B(n_27), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_20), .Y(n_32) );
INVx1_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
NAND2xp5_ASAP7_75t_L g34 ( .A(n_32), .B(n_25), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
OAI322xp33_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_24), .A3(n_18), .B1(n_22), .B2(n_13), .C1(n_25), .C2(n_8), .Y(n_36) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
OAI211xp5_ASAP7_75t_SL g38 ( .A1(n_36), .A2(n_24), .B(n_33), .C(n_22), .Y(n_38) );
INVx2_ASAP7_75t_L g39 ( .A(n_37), .Y(n_39) );
AOI22xp5_ASAP7_75t_SL g40 ( .A1(n_39), .A2(n_38), .B1(n_22), .B2(n_10), .Y(n_40) );
endmodule