module fake_jpeg_17144_n_385 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_385);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_385;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_43),
.Y(n_114)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_44),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_30),
.Y(n_52)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_33),
.A2(n_13),
.B1(n_1),
.B2(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_53),
.A2(n_37),
.B1(n_36),
.B2(n_19),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_23),
.Y(n_54)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_0),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_58),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_0),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_33),
.B1(n_20),
.B2(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_97),
.B1(n_42),
.B2(n_49),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_74),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_34),
.B(n_21),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_111),
.C(n_28),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_79),
.B(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_17),
.Y(n_80)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_14),
.Y(n_85)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_14),
.Y(n_87)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_28),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_90),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_98),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_95),
.B(n_96),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_45),
.B(n_21),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_33),
.B1(n_37),
.B2(n_22),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_17),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_99),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_32),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_18),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_109),
.A2(n_30),
.B(n_5),
.C(n_7),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_56),
.B(n_19),
.Y(n_111)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_83),
.B1(n_10),
.B2(n_11),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_97),
.B1(n_102),
.B2(n_75),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_122),
.A2(n_125),
.B1(n_140),
.B2(n_144),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_123),
.B(n_27),
.C(n_10),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_44),
.B1(n_64),
.B2(n_59),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_126),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_71),
.A2(n_36),
.B1(n_108),
.B2(n_31),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_127),
.A2(n_145),
.B1(n_167),
.B2(n_9),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_31),
.B1(n_36),
.B2(n_23),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_139),
.B1(n_168),
.B2(n_5),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_92),
.B1(n_100),
.B2(n_41),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_162),
.B1(n_105),
.B2(n_107),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_66),
.Y(n_130)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_24),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_135),
.B(n_138),
.C(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_27),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_143),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_24),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_75),
.A2(n_35),
.B1(n_25),
.B2(n_51),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_78),
.A2(n_65),
.B1(n_55),
.B2(n_40),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_29),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_102),
.A2(n_35),
.B1(n_25),
.B2(n_29),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_71),
.A2(n_13),
.B1(n_35),
.B2(n_25),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_29),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_157),
.Y(n_181)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_77),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_148),
.B(n_155),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_35),
.B1(n_29),
.B2(n_27),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_149),
.A2(n_150),
.B1(n_10),
.B2(n_11),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_84),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_30),
.B(n_29),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_66),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_156),
.Y(n_183)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_66),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_68),
.B(n_29),
.Y(n_157)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_160),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_68),
.Y(n_160)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_161),
.A2(n_164),
.B(n_120),
.C(n_155),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_30),
.B1(n_27),
.B2(n_7),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_98),
.A2(n_4),
.B(n_5),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_150),
.B(n_162),
.Y(n_198)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_108),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_100),
.A2(n_27),
.B1(n_7),
.B2(n_8),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_133),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_170),
.A2(n_176),
.B1(n_192),
.B2(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_138),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_194),
.C(n_130),
.Y(n_236)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_124),
.B(n_114),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_125),
.B(n_8),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_198),
.B(n_207),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_122),
.A2(n_106),
.B1(n_112),
.B2(n_101),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_114),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_105),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_142),
.B(n_91),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_118),
.B(n_91),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_131),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_121),
.B(n_82),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_134),
.B(n_9),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_204),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_121),
.B(n_132),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_148),
.Y(n_230)
);

O2A1O1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_161),
.A2(n_83),
.B(n_101),
.C(n_112),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_126),
.B1(n_130),
.B2(n_170),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_140),
.Y(n_232)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_141),
.B(n_9),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g225 ( 
.A(n_211),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_187),
.B1(n_196),
.B2(n_161),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_213),
.A2(n_154),
.B(n_120),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_157),
.B(n_11),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g241 ( 
.A(n_214),
.Y(n_241)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_228),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_224),
.A2(n_231),
.B1(n_244),
.B2(n_207),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_161),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_236),
.C(n_240),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_219),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_165),
.B1(n_144),
.B2(n_149),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_232),
.A2(n_235),
.B1(n_221),
.B2(n_255),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_234),
.A2(n_198),
.B(n_192),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_169),
.B(n_159),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_238),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_239),
.A2(n_232),
.B1(n_223),
.B2(n_233),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_181),
.C(n_194),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_250),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_187),
.A2(n_189),
.B1(n_182),
.B2(n_184),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_180),
.B(n_181),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_212),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_203),
.B(n_190),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_180),
.B(n_175),
.C(n_205),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_179),
.Y(n_274)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_178),
.Y(n_252)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_252),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_195),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_202),
.B(n_188),
.Y(n_256)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_213),
.B(n_216),
.C(n_236),
.D(n_240),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_257),
.A2(n_258),
.B(n_262),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_260),
.B(n_266),
.Y(n_309)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_268),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_184),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_263),
.A2(n_270),
.B1(n_248),
.B2(n_249),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_276),
.Y(n_299)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_207),
.B1(n_174),
.B2(n_185),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_242),
.A2(n_172),
.B1(n_210),
.B2(n_171),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_287),
.B1(n_288),
.B2(n_252),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_219),
.B(n_171),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_273),
.A2(n_277),
.B(n_282),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_281),
.C(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_172),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_185),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_280),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_231),
.A2(n_224),
.B1(n_227),
.B2(n_237),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_279),
.A2(n_283),
.B1(n_284),
.B2(n_270),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_233),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_216),
.A2(n_234),
.B(n_223),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_284),
.B(n_258),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_232),
.A2(n_222),
.B(n_220),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_246),
.Y(n_285)
);

OA22x2_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_267),
.B1(n_268),
.B2(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_286),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_221),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_247),
.Y(n_290)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_290),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_295),
.C(n_296),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_293),
.A2(n_286),
.B(n_289),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_241),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_218),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_248),
.C(n_249),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_298),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_225),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_269),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_308),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_302),
.B1(n_285),
.B2(n_269),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_247),
.B1(n_254),
.B2(n_288),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_303),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_305),
.B(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_260),
.C(n_280),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_307),
.B(n_315),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_290),
.Y(n_312)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_287),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_317),
.B(n_318),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_273),
.C(n_283),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_319),
.A2(n_323),
.B(n_324),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_320),
.A2(n_293),
.B1(n_302),
.B2(n_314),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_294),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_333),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_304),
.B(n_318),
.Y(n_324)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_313),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_334),
.B(n_337),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_292),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_335),
.B(n_308),
.Y(n_343)
);

XNOR2x1_ASAP7_75t_L g336 ( 
.A(n_311),
.B(n_275),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_336),
.B(n_315),
.Y(n_341)
);

INVxp33_ASAP7_75t_L g337 ( 
.A(n_306),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_334),
.B(n_278),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_340),
.B(n_346),
.Y(n_358)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_291),
.C(n_331),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_347),
.C(n_348),
.Y(n_359)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_311),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_296),
.C(n_297),
.Y(n_348)
);

OAI322xp33_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_309),
.A3(n_298),
.B1(n_310),
.B2(n_295),
.C1(n_307),
.C2(n_317),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_350),
.A2(n_355),
.B1(n_356),
.B2(n_345),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_326),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_353),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_309),
.C(n_264),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_325),
.A2(n_328),
.B1(n_320),
.B2(n_324),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_329),
.C(n_319),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_362),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_345),
.A2(n_325),
.B(n_337),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_361),
.A2(n_365),
.B(n_355),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_344),
.A2(n_327),
.B1(n_323),
.B2(n_339),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_344),
.A2(n_330),
.B1(n_338),
.B2(n_306),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_363),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_264),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_351),
.A2(n_329),
.B1(n_354),
.B2(n_349),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_367),
.B(n_353),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_342),
.C(n_348),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_372),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_371),
.A2(n_364),
.B(n_365),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_356),
.C(n_347),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_364),
.C(n_357),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_369),
.A2(n_358),
.B1(n_362),
.B2(n_366),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_376),
.C(n_377),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_376),
.B(n_369),
.C(n_370),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_379),
.B(n_374),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_380),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_381),
.A2(n_378),
.B(n_365),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_382),
.B(n_361),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_383),
.A2(n_363),
.B(n_341),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_384),
.B(n_346),
.Y(n_385)
);


endmodule