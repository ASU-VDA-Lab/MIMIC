module fake_jpeg_30519_n_318 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_318);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_4),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_46),
.B(n_50),
.Y(n_108)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_52),
.B(n_54),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_33),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_59),
.B(n_61),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_69),
.Y(n_86)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_70),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_30),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_30),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_28),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_65),
.B1(n_60),
.B2(n_56),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_35),
.B1(n_23),
.B2(n_42),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_23),
.B1(n_39),
.B2(n_40),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_35),
.B1(n_42),
.B2(n_24),
.Y(n_80)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_39),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_83),
.B(n_94),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_42),
.B1(n_24),
.B2(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_84),
.A2(n_88),
.B1(n_89),
.B2(n_101),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_40),
.B1(n_43),
.B2(n_41),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_43),
.B1(n_34),
.B2(n_28),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_34),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_15),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_24),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_45),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_22),
.B1(n_36),
.B2(n_2),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_111),
.Y(n_148)
);

CKINVDCx9p33_ASAP7_75t_R g105 ( 
.A(n_54),
.Y(n_105)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_51),
.A2(n_22),
.B1(n_1),
.B2(n_3),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_110),
.A2(n_113),
.B1(n_55),
.B2(n_64),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_24),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_117),
.B(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_98),
.B(n_13),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_127),
.Y(n_163)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_133),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_81),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_56),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_130),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_12),
.B(n_3),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_138),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_86),
.C(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_70),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_137),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_0),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_5),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_5),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_146),
.Y(n_183)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_75),
.B(n_53),
.C(n_49),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_6),
.Y(n_147)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_75),
.B(n_99),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_99),
.B(n_7),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_139),
.B1(n_117),
.B2(n_130),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_126),
.A2(n_51),
.B1(n_107),
.B2(n_114),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_128),
.A2(n_114),
.B1(n_107),
.B2(n_92),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_103),
.B(n_91),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_162),
.B(n_181),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_87),
.B(n_96),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_182),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_138),
.A2(n_87),
.B1(n_96),
.B2(n_10),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_175),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_9),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_133),
.B(n_153),
.Y(n_181)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_122),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_192),
.B(n_206),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_146),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_181),
.A2(n_131),
.B(n_133),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_203),
.B(n_154),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_143),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_157),
.B(n_116),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_143),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_204),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_133),
.B(n_119),
.Y(n_203)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_171),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_121),
.C(n_135),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_214),
.C(n_167),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_134),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_152),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_161),
.B(n_162),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_170),
.B(n_141),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_212),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_132),
.C(n_118),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_180),
.B(n_125),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_180),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_217),
.A2(n_231),
.B(n_234),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_222),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_206),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_SL g227 ( 
.A1(n_198),
.A2(n_175),
.B(n_155),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_227),
.A2(n_229),
.B(n_233),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_187),
.A2(n_210),
.B1(n_209),
.B2(n_213),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_168),
.Y(n_230)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_164),
.B(n_168),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_203),
.A2(n_188),
.B1(n_198),
.B2(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_207),
.B(n_195),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_172),
.B(n_185),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_196),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_214),
.C(n_205),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_246),
.C(n_251),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_199),
.C(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_258),
.B1(n_228),
.B2(n_216),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_191),
.C(n_215),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_189),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_224),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_189),
.C(n_211),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_218),
.C(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_216),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_172),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_223),
.Y(n_267)
);

NAND4xp25_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_223),
.C(n_169),
.D(n_124),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_257),
.A2(n_217),
.B(n_232),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_247),
.B(n_248),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_273),
.Y(n_278)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_272),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_231),
.C(n_222),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_251),
.C(n_256),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_204),
.B1(n_220),
.B2(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_236),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_246),
.B(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_252),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_268),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_276),
.B(n_281),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_265),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_247),
.C(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_260),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_286),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_248),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_280),
.B(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_266),
.C(n_272),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_271),
.C(n_262),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_263),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_295),
.C(n_275),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_265),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_296),
.A2(n_297),
.B(n_224),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_278),
.B(n_249),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_284),
.A3(n_276),
.B1(n_258),
.B2(n_245),
.C1(n_204),
.C2(n_243),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_300),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g300 ( 
.A(n_296),
.B(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_301),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_304),
.B(n_294),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_245),
.C(n_243),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_305),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_295),
.B1(n_190),
.B2(n_197),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_309),
.Y(n_313)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_200),
.B(n_202),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_310),
.B(n_188),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_312),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_308),
.A2(n_186),
.B1(n_178),
.B2(n_142),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_178),
.B(n_306),
.C(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_311),
.C(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_311),
.Y(n_318)
);


endmodule