module fake_netlist_5_2160_n_1833 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1833);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1833;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_43),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_127),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_1),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_46),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_141),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_14),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_28),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_21),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_19),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_158),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_28),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_87),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_93),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_60),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_33),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_77),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_121),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_139),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_35),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_59),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_4),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_34),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_53),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_21),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_34),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_110),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_114),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_123),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_69),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_116),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_32),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_8),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_17),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_74),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_29),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_18),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_108),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_166),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_3),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_4),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_68),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_62),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_79),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_40),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_86),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_3),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_48),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_151),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_63),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_26),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_99),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_133),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_19),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_142),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_78),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_113),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_103),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_85),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_132),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_171),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_5),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_102),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_64),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_1),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_44),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_163),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_161),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_37),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_100),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_29),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_26),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_91),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_73),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_160),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_80),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_43),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_106),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_27),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_57),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_152),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_136),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_96),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_67),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_41),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_47),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_55),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_2),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_140),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_76),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_18),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_14),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_130),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_170),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_65),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_56),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_24),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_167),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_173),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_137),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_9),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_0),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_70),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_95),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_145),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_107),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_31),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_38),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_72),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_83),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_88),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_11),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_155),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_46),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_92),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_101),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_176),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_148),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_90),
.B(n_172),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_94),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_7),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_61),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_104),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_52),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_22),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_144),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_89),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_7),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_33),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_49),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_52),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_154),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_0),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_115),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_51),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_71),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_17),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_42),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_111),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_31),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_20),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_36),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_6),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_45),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_81),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_128),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_134),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_165),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_39),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_55),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_150),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_212),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_219),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_193),
.B(n_2),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_227),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_232),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_214),
.B(n_6),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_245),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_214),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_214),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_246),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_354),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_200),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_274),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_247),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_242),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_214),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_263),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_214),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_261),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_204),
.B(n_8),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_241),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_214),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_274),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_290),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_214),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_267),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_316),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_214),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_193),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_197),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_279),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_222),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_281),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_197),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_185),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_250),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_250),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_274),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_329),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_329),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_282),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_351),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_275),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_338),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_210),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_254),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_211),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_213),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_338),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_287),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_317),
.B(n_9),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_254),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_297),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_301),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_195),
.B(n_10),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_254),
.Y(n_413)
);

INVx4_ASAP7_75t_R g414 ( 
.A(n_323),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_254),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_340),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_215),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_305),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_254),
.Y(n_419)
);

CKINVDCx16_ASAP7_75t_R g420 ( 
.A(n_340),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_306),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_201),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_256),
.B(n_323),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_203),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_218),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_216),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_192),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_308),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_221),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_228),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_194),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_238),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_328),
.B(n_10),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_185),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_239),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_319),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_188),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_243),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_194),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_206),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_203),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_188),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_270),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_189),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_272),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_223),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_427),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_427),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_403),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_378),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_365),
.B(n_328),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_190),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_381),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_384),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_419),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_431),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_376),
.B(n_203),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_362),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_431),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_187),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_R g472 ( 
.A(n_442),
.B(n_189),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_439),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_440),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_440),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_359),
.B(n_190),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_425),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_430),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_432),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_R g481 ( 
.A(n_442),
.B(n_191),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_359),
.B(n_230),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_443),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_445),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_385),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_412),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_367),
.A2(n_220),
.B1(n_229),
.B2(n_233),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_433),
.B(n_186),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g493 ( 
.A1(n_429),
.A2(n_273),
.B(n_206),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_390),
.B(n_230),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_392),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_393),
.B(n_264),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_424),
.B(n_231),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_444),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_377),
.B(n_196),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_395),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_401),
.B(n_264),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_406),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_391),
.B(n_283),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_283),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_369),
.B(n_296),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_444),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_357),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_296),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_357),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_402),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_358),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_358),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_379),
.B(n_324),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_360),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_360),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_361),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_361),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_363),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_363),
.B(n_179),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_366),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_366),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_234),
.B1(n_312),
.B2(n_273),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_487),
.B(n_180),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_457),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_468),
.B(n_370),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_487),
.B(n_370),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_487),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

AND3x2_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_355),
.C(n_509),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_450),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_457),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_452),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_467),
.B(n_388),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_452),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_487),
.B(n_181),
.Y(n_539)
);

BUFx6f_ASAP7_75t_SL g540 ( 
.A(n_508),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_493),
.B(n_182),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_487),
.B(n_183),
.Y(n_543)
);

BUFx4f_ASAP7_75t_L g544 ( 
.A(n_493),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_467),
.B(n_404),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_487),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_450),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_450),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_493),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_457),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_487),
.Y(n_552)
);

AO21x2_ASAP7_75t_L g553 ( 
.A1(n_468),
.A2(n_198),
.B(n_184),
.Y(n_553)
);

AOI21x1_ASAP7_75t_L g554 ( 
.A1(n_459),
.A2(n_453),
.B(n_468),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_451),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_451),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_508),
.B(n_441),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_492),
.B(n_405),
.Y(n_558)
);

BUFx10_ASAP7_75t_L g559 ( 
.A(n_499),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_499),
.B(n_420),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_487),
.A2(n_234),
.B1(n_312),
.B2(n_294),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_457),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_513),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_476),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_451),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_484),
.A2(n_476),
.B1(n_489),
.B2(n_493),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_513),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_455),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_455),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_498),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_515),
.B(n_373),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_515),
.B(n_288),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_455),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_472),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_373),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_484),
.A2(n_346),
.B1(n_291),
.B2(n_295),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_450),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_493),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_456),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_484),
.A2(n_313),
.B1(n_333),
.B2(n_300),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_461),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_456),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_463),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_510),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_451),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_463),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_484),
.A2(n_342),
.B1(n_343),
.B2(n_180),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_515),
.B(n_382),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_456),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_489),
.B(n_382),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_463),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_512),
.A2(n_446),
.B1(n_417),
.B2(n_426),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_515),
.B(n_387),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_484),
.B(n_387),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_451),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_509),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_493),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_517),
.B(n_389),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_463),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_451),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_464),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_464),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_490),
.B(n_368),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_451),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_471),
.B(n_389),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_464),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_471),
.B(n_398),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_398),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_464),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_451),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_476),
.B(n_407),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_493),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_517),
.B(n_407),
.Y(n_617)
);

INVxp33_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_476),
.A2(n_180),
.B1(n_253),
.B2(n_289),
.Y(n_619)
);

BUFx6f_ASAP7_75t_SL g620 ( 
.A(n_516),
.Y(n_620)
);

INVxp33_ASAP7_75t_SL g621 ( 
.A(n_490),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_451),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_458),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_447),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_522),
.B(n_410),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_472),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_522),
.B(n_410),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_458),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_458),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_460),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_512),
.B(n_411),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_517),
.B(n_411),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_514),
.B(n_418),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_517),
.B(n_180),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_522),
.B(n_418),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_523),
.B(n_421),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_447),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_523),
.B(n_421),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_460),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_489),
.A2(n_400),
.B1(n_428),
.B2(n_436),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_501),
.Y(n_641)
);

BUFx8_ASAP7_75t_SL g642 ( 
.A(n_510),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_509),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_488),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_501),
.Y(n_645)
);

NAND2xp33_ASAP7_75t_L g646 ( 
.A(n_489),
.B(n_180),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_447),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_488),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_501),
.Y(n_649)
);

INVxp33_ASAP7_75t_L g650 ( 
.A(n_490),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_506),
.B(n_428),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_501),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_516),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_506),
.B(n_436),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_501),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_506),
.B(n_224),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_514),
.A2(n_266),
.B1(n_396),
.B2(n_394),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_516),
.B(n_225),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_460),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_501),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_477),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_514),
.B(n_416),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_523),
.B(n_191),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_519),
.B(n_399),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_462),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_488),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_519),
.B(n_521),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_491),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_479),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_524),
.B(n_326),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_462),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_523),
.B(n_253),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_462),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_519),
.B(n_371),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_524),
.B(n_516),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_SL g676 ( 
.A1(n_453),
.A2(n_284),
.B(n_350),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_623),
.Y(n_677)
);

NOR2xp67_ASAP7_75t_L g678 ( 
.A(n_595),
.B(n_518),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_567),
.A2(n_524),
.B1(n_520),
.B2(n_521),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_662),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_600),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_623),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_548),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_520),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_545),
.B(n_518),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_609),
.B(n_524),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_564),
.B(n_520),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_526),
.B(n_520),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_611),
.B(n_520),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_L g690 ( 
.A(n_558),
.B(n_521),
.C(n_481),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_526),
.B(n_520),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_626),
.B(n_625),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_530),
.B(n_516),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_593),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_531),
.B(n_192),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_644),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_628),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_593),
.B(n_510),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_530),
.B(n_518),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_539),
.A2(n_516),
.B1(n_505),
.B2(n_511),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_544),
.B(n_518),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_531),
.B(n_192),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_547),
.B(n_518),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_544),
.B(n_518),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_628),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_644),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_547),
.B(n_504),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_539),
.A2(n_505),
.B1(n_504),
.B2(n_511),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_627),
.B(n_497),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_552),
.B(n_504),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_635),
.B(n_497),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_548),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_534),
.B(n_503),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_552),
.B(n_504),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_612),
.B(n_375),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_631),
.B(n_380),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_667),
.B(n_505),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_559),
.B(n_505),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_559),
.B(n_511),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_629),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_600),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_675),
.B(n_511),
.Y(n_722)
);

OAI22xp33_ASAP7_75t_L g723 ( 
.A1(n_528),
.A2(n_481),
.B1(n_383),
.B2(n_502),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_576),
.B(n_540),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_648),
.B(n_479),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_643),
.Y(n_726)
);

BUFx12f_ASAP7_75t_SL g727 ( 
.A(n_574),
.Y(n_727)
);

BUFx4f_ASAP7_75t_L g728 ( 
.A(n_653),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_648),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_633),
.B(n_507),
.C(n_495),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_666),
.B(n_479),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_578),
.A2(n_453),
.B1(n_495),
.B2(n_491),
.C(n_500),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_666),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_587),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_668),
.B(n_479),
.Y(n_735)
);

AND2x4_ASAP7_75t_SL g736 ( 
.A(n_546),
.B(n_231),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_668),
.B(n_479),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_549),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_559),
.B(n_507),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_544),
.B(n_253),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_643),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_539),
.B(n_486),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_629),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_L g744 ( 
.A(n_640),
.B(n_507),
.C(n_495),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_630),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_576),
.B(n_507),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_630),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_550),
.B(n_253),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_651),
.B(n_507),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_618),
.B(n_507),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_639),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_543),
.B(n_615),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_550),
.B(n_253),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_SL g754 ( 
.A1(n_621),
.A2(n_326),
.B1(n_330),
.B2(n_334),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_654),
.B(n_187),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_L g756 ( 
.A1(n_574),
.A2(n_577),
.B1(n_597),
.B2(n_663),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_560),
.B(n_199),
.Y(n_757)
);

NAND3xp33_ASAP7_75t_SL g758 ( 
.A(n_537),
.B(n_334),
.C(n_330),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_534),
.B(n_503),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_543),
.B(n_579),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_639),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_550),
.B(n_459),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_659),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_563),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_664),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_663),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_659),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_580),
.B(n_459),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_580),
.B(n_543),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_579),
.B(n_486),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_665),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_665),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_548),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_601),
.Y(n_774)
);

NAND3xp33_ASAP7_75t_L g775 ( 
.A(n_670),
.B(n_500),
.C(n_491),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_608),
.B(n_601),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_553),
.A2(n_486),
.B1(n_477),
.B2(n_255),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_580),
.B(n_477),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_SL g779 ( 
.A1(n_621),
.A2(n_345),
.B1(n_335),
.B2(n_336),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_674),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_670),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_671),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_671),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_616),
.B(n_477),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_616),
.B(n_486),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_574),
.B(n_486),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_653),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_673),
.Y(n_788)
);

INVxp33_ASAP7_75t_SL g789 ( 
.A(n_563),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_548),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_658),
.B(n_500),
.C(n_496),
.Y(n_791)
);

AND2x2_ASAP7_75t_SL g792 ( 
.A(n_525),
.B(n_646),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_673),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_548),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_568),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_574),
.B(n_486),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_527),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_653),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_542),
.B(n_192),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_527),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_669),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_653),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_554),
.B(n_477),
.Y(n_803)
);

CKINVDCx16_ASAP7_75t_R g804 ( 
.A(n_568),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_620),
.A2(n_260),
.B1(n_244),
.B2(n_240),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_620),
.A2(n_265),
.B1(n_235),
.B2(n_217),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_546),
.B(n_503),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_573),
.B(n_199),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_546),
.B(n_503),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_554),
.B(n_477),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_553),
.B(n_478),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_535),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_591),
.B(n_202),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_535),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_624),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_624),
.B(n_477),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_L g817 ( 
.A(n_542),
.B(n_192),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_641),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_604),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_641),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_596),
.B(n_494),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_551),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_542),
.B(n_624),
.Y(n_823)
);

INVx4_ASAP7_75t_L g824 ( 
.A(n_604),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_SL g825 ( 
.A(n_604),
.B(n_208),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_551),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_562),
.Y(n_827)
);

NAND3xp33_ASAP7_75t_L g828 ( 
.A(n_602),
.B(n_502),
.C(n_496),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_617),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_637),
.B(n_477),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_637),
.B(n_477),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_637),
.B(n_447),
.Y(n_832)
);

BUFx12f_ASAP7_75t_L g833 ( 
.A(n_634),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_634),
.B(n_192),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_SL g835 ( 
.A1(n_632),
.A2(n_335),
.B1(n_336),
.B2(n_345),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_647),
.B(n_447),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_647),
.B(n_447),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_636),
.B(n_202),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_553),
.A2(n_325),
.B1(n_322),
.B2(n_315),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_645),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_647),
.B(n_656),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_645),
.B(n_192),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_562),
.Y(n_843)
);

A2O1A1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_650),
.A2(n_502),
.B(n_496),
.C(n_494),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_565),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_649),
.B(n_652),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_765),
.B(n_557),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_762),
.A2(n_646),
.B(n_638),
.Y(n_848)
);

BUFx12f_ASAP7_75t_L g849 ( 
.A(n_795),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_709),
.A2(n_572),
.B1(n_620),
.B2(n_540),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_677),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_762),
.A2(n_614),
.B(n_604),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_686),
.B(n_619),
.Y(n_853)
);

AOI21xp33_ASAP7_75t_L g854 ( 
.A1(n_711),
.A2(n_757),
.B(n_716),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_768),
.A2(n_614),
.B(n_604),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_721),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_768),
.A2(n_614),
.B(n_556),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_801),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_789),
.B(n_764),
.Y(n_859)
);

INVx11_ASAP7_75t_L g860 ( 
.A(n_833),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_692),
.B(n_572),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_680),
.B(n_533),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_785),
.A2(n_652),
.B(n_649),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_760),
.A2(n_614),
.B(n_556),
.Y(n_864)
);

BUFx4f_ASAP7_75t_L g865 ( 
.A(n_746),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_689),
.A2(n_590),
.B1(n_561),
.B2(n_540),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_776),
.A2(n_614),
.B(n_556),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_717),
.B(n_583),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_679),
.A2(n_655),
.B1(n_660),
.B2(n_657),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_778),
.A2(n_566),
.B(n_555),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_778),
.A2(n_566),
.B(n_555),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_769),
.A2(n_752),
.B(n_823),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_769),
.A2(n_566),
.B(n_555),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_698),
.B(n_607),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_780),
.B(n_607),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_844),
.A2(n_676),
.B(n_494),
.C(n_603),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_844),
.A2(n_603),
.B(n_605),
.C(n_613),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_823),
.A2(n_598),
.B(n_588),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_688),
.A2(n_691),
.B1(n_693),
.B2(n_700),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_749),
.A2(n_655),
.B(n_660),
.C(n_310),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_688),
.A2(n_293),
.B1(n_299),
.B2(n_292),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_694),
.B(n_205),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_734),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_821),
.B(n_588),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_690),
.B(n_205),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_781),
.B(n_588),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_682),
.Y(n_887)
);

O2A1O1Ixp5_ASAP7_75t_L g888 ( 
.A1(n_691),
.A2(n_565),
.B(n_571),
.C(n_582),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_802),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_707),
.B(n_598),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_723),
.B(n_207),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_784),
.A2(n_622),
.B(n_598),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_784),
.A2(n_622),
.B(n_661),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_841),
.A2(n_622),
.B(n_661),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_740),
.A2(n_661),
.B(n_582),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_726),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_740),
.A2(n_661),
.B(n_584),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_808),
.A2(n_286),
.B(n_280),
.C(n_258),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_685),
.B(n_207),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_748),
.A2(n_661),
.B(n_584),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_710),
.B(n_605),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_748),
.A2(n_571),
.B(n_586),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_753),
.A2(n_586),
.B(n_589),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_813),
.A2(n_252),
.B(n_613),
.C(n_610),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_714),
.B(n_606),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_753),
.A2(n_589),
.B(n_594),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_766),
.B(n_606),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_SL g908 ( 
.A(n_789),
.B(n_642),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_722),
.B(n_610),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_838),
.A2(n_541),
.B(n_599),
.C(n_529),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_718),
.B(n_478),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_828),
.A2(n_541),
.B(n_599),
.C(n_529),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_684),
.B(n_594),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_687),
.B(n_532),
.Y(n_914)
);

OAI21xp33_ASAP7_75t_L g915 ( 
.A1(n_708),
.A2(n_719),
.B(n_715),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_755),
.B(n_532),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_741),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_739),
.B(n_209),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_678),
.B(n_209),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_774),
.A2(n_575),
.B(n_592),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_815),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_774),
.B(n_536),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_791),
.A2(n_569),
.B(n_592),
.C(n_585),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_774),
.A2(n_570),
.B(n_585),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_818),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_815),
.Y(n_926)
);

OR2x2_ASAP7_75t_L g927 ( 
.A(n_681),
.B(n_478),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_799),
.A2(n_581),
.B(n_575),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_802),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_829),
.B(n_268),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_799),
.A2(n_581),
.B(n_570),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_807),
.B(n_268),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_817),
.A2(n_569),
.B(n_538),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_809),
.B(n_536),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_699),
.A2(n_538),
.B1(n_332),
.B2(n_320),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_758),
.B(n_347),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_697),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_817),
.A2(n_448),
.B(n_449),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_SL g939 ( 
.A1(n_795),
.A2(n_347),
.B1(n_348),
.B2(n_349),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_802),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_792),
.A2(n_672),
.B1(n_634),
.B2(n_192),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_803),
.A2(n_449),
.B(n_454),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_742),
.A2(n_448),
.B(n_449),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_820),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_802),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_792),
.B(n_634),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_824),
.A2(n_448),
.B(n_454),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_756),
.A2(n_483),
.B(n_485),
.C(n_482),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_824),
.A2(n_448),
.B(n_454),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_824),
.A2(n_448),
.B(n_485),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_696),
.B(n_706),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_729),
.B(n_634),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_733),
.B(n_811),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_803),
.A2(n_810),
.B(n_811),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_811),
.B(n_634),
.Y(n_955)
);

CKINVDCx6p67_ASAP7_75t_R g956 ( 
.A(n_804),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_840),
.Y(n_957)
);

AO21x1_ASAP7_75t_L g958 ( 
.A1(n_699),
.A2(n_465),
.B(n_470),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_750),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_833),
.B(n_483),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_810),
.A2(n_465),
.B(n_474),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_701),
.A2(n_331),
.B1(n_320),
.B2(n_321),
.Y(n_962)
);

O2A1O1Ixp5_ASAP7_75t_L g963 ( 
.A1(n_842),
.A2(n_480),
.B(n_485),
.C(n_482),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_728),
.A2(n_448),
.B(n_485),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_815),
.B(n_321),
.Y(n_965)
);

O2A1O1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_732),
.A2(n_483),
.B(n_482),
.C(n_480),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_738),
.B(n_634),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_L g968 ( 
.A(n_744),
.B(n_672),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_713),
.B(n_672),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_728),
.A2(n_482),
.B(n_480),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_728),
.A2(n_480),
.B(n_465),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_697),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_705),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_736),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_701),
.A2(n_327),
.B1(n_331),
.B2(n_332),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_730),
.A2(n_672),
.B1(n_226),
.B2(n_304),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_835),
.B(n_348),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_724),
.B(n_736),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_764),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_775),
.B(n_327),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_713),
.A2(n_672),
.B1(n_311),
.B2(n_309),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_770),
.A2(n_466),
.B(n_475),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_786),
.A2(n_337),
.B(n_339),
.C(n_341),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_842),
.A2(n_475),
.B(n_474),
.C(n_473),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_846),
.A2(n_672),
.B(n_470),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_713),
.B(n_672),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_846),
.A2(n_470),
.B(n_475),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_705),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_703),
.A2(n_475),
.B(n_474),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_759),
.B(n_236),
.Y(n_990)
);

INVxp67_ASAP7_75t_SL g991 ( 
.A(n_819),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_839),
.A2(n_349),
.B(n_339),
.Y(n_992)
);

OAI321xp33_ASAP7_75t_L g993 ( 
.A1(n_754),
.A2(n_474),
.A3(n_473),
.B1(n_469),
.B2(n_466),
.C(n_307),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_787),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_683),
.A2(n_473),
.B(n_469),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_720),
.Y(n_996)
);

INVx11_ASAP7_75t_L g997 ( 
.A(n_727),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_683),
.A2(n_473),
.B(n_469),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_831),
.A2(n_469),
.B(n_466),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_727),
.B(n_337),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_720),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_759),
.Y(n_1002)
);

NOR2x2_ASAP7_75t_L g1003 ( 
.A(n_779),
.B(n_231),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_759),
.B(n_237),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_831),
.A2(n_466),
.B(n_356),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_743),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_683),
.A2(n_278),
.B(n_251),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_743),
.B(n_248),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_745),
.B(n_298),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_712),
.A2(n_285),
.B(n_259),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_773),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_704),
.B(n_353),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_796),
.Y(n_1013)
);

OAI21xp33_ASAP7_75t_L g1014 ( 
.A1(n_805),
.A2(n_777),
.B(n_806),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_745),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_751),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_725),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_751),
.B(n_763),
.Y(n_1018)
);

AO21x1_ASAP7_75t_L g1019 ( 
.A1(n_704),
.A2(n_249),
.B(n_307),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_712),
.A2(n_302),
.B(n_262),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_712),
.A2(n_303),
.B(n_269),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_763),
.B(n_314),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_L g1023 ( 
.A1(n_747),
.A2(n_761),
.B(n_767),
.C(n_772),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_771),
.B(n_318),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_771),
.B(n_277),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_787),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_731),
.B(n_352),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_782),
.B(n_257),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_798),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_782),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_735),
.A2(n_271),
.B(n_276),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_737),
.A2(n_819),
.B(n_832),
.Y(n_1032)
);

CKINVDCx16_ASAP7_75t_R g1033 ( 
.A(n_798),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_783),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_783),
.B(n_788),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_854),
.B(n_819),
.Y(n_1036)
);

AOI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_853),
.A2(n_793),
.B(n_702),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_R g1038 ( 
.A(n_1033),
.B(n_859),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_915),
.A2(n_837),
.B(n_836),
.C(n_695),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_959),
.B(n_794),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_994),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_865),
.B(n_819),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_994),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_874),
.B(n_249),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_851),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_861),
.B(n_794),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_959),
.B(n_797),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_883),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_875),
.A2(n_695),
.B1(n_702),
.B2(n_794),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_875),
.B(n_773),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_917),
.B(n_773),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_1014),
.A2(n_816),
.B(n_830),
.C(n_812),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_974),
.B(n_341),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_SL g1054 ( 
.A1(n_850),
.A2(n_344),
.B1(n_352),
.B2(n_353),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_872),
.A2(n_773),
.B(n_790),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_865),
.B(n_790),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_856),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_911),
.B(n_845),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1013),
.B(n_845),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_891),
.A2(n_936),
.B(n_885),
.C(n_898),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_858),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_954),
.A2(n_790),
.B(n_834),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1013),
.B(n_843),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_848),
.A2(n_843),
.B(n_797),
.C(n_827),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_922),
.A2(n_790),
.B(n_834),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_979),
.B(n_827),
.Y(n_1066)
);

OA21x2_ASAP7_75t_L g1067 ( 
.A1(n_863),
.A2(n_826),
.B(n_800),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_934),
.A2(n_826),
.B(n_822),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_856),
.B(n_822),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_868),
.A2(n_814),
.B1(n_812),
.B2(n_800),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_994),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_850),
.A2(n_879),
.B1(n_953),
.B2(n_941),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_896),
.B(n_814),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_936),
.A2(n_344),
.B(n_825),
.C(n_307),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_994),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_847),
.A2(n_249),
.B1(n_178),
.B2(n_168),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1017),
.B(n_11),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_896),
.B(n_12),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_862),
.B(n_978),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_909),
.A2(n_164),
.B(n_156),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_862),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_955),
.A2(n_143),
.B(n_138),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_SL g1083 ( 
.A1(n_946),
.A2(n_126),
.B(n_125),
.C(n_124),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_977),
.A2(n_13),
.B(n_15),
.C(n_16),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1017),
.B(n_13),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_849),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_914),
.A2(n_117),
.B(n_97),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_930),
.B(n_15),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_941),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_916),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_925),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_944),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_876),
.A2(n_23),
.B(n_25),
.C(n_27),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_957),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_973),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_1026),
.B(n_84),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_927),
.B(n_30),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_890),
.A2(n_82),
.B(n_75),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_968),
.A2(n_867),
.B(n_884),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_901),
.B(n_905),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_956),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_1000),
.B(n_30),
.Y(n_1102)
);

NAND2xp33_ASAP7_75t_SL g1103 ( 
.A(n_1026),
.B(n_1029),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_919),
.A2(n_66),
.B1(n_35),
.B2(n_36),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1000),
.B(n_32),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_977),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_1106)
);

INVx4_ASAP7_75t_L g1107 ( 
.A(n_1026),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_887),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_939),
.B(n_42),
.C(n_45),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_932),
.B(n_47),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_961),
.A2(n_48),
.B(n_49),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_882),
.B(n_50),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_993),
.B(n_50),
.C(n_51),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_960),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_907),
.B(n_53),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_SL g1116 ( 
.A(n_889),
.B(n_54),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_918),
.B(n_54),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_907),
.A2(n_56),
.B1(n_58),
.B2(n_1002),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_886),
.B(n_58),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_886),
.B(n_1027),
.Y(n_1120)
);

OA22x2_ASAP7_75t_L g1121 ( 
.A1(n_1003),
.A2(n_951),
.B1(n_992),
.B2(n_960),
.Y(n_1121)
);

AOI21x1_ASAP7_75t_SL g1122 ( 
.A1(n_967),
.A2(n_952),
.B(n_986),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_980),
.A2(n_983),
.B(n_965),
.C(n_869),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1027),
.B(n_1002),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_SL g1125 ( 
.A1(n_881),
.A2(n_966),
.B1(n_866),
.B2(n_877),
.C(n_948),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1026),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_965),
.B(n_921),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_913),
.A2(n_894),
.B(n_864),
.Y(n_1128)
);

NOR2x1_ASAP7_75t_L g1129 ( 
.A(n_889),
.B(n_929),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_921),
.B(n_926),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_926),
.B(n_991),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1012),
.A2(n_880),
.B(n_904),
.C(n_910),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1012),
.A2(n_975),
.B(n_962),
.C(n_935),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1006),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1019),
.A2(n_1004),
.B1(n_990),
.B2(n_1008),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_943),
.A2(n_1032),
.B(n_1023),
.C(n_963),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_937),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_908),
.B(n_1009),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1029),
.B(n_940),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1029),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_972),
.Y(n_1141)
);

INVx4_ASAP7_75t_L g1142 ( 
.A(n_1029),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_960),
.B(n_988),
.Y(n_1143)
);

AO32x2_ASAP7_75t_L g1144 ( 
.A1(n_929),
.A2(n_958),
.A3(n_888),
.B1(n_1023),
.B2(n_1005),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_940),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_996),
.B(n_1001),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_SL g1147 ( 
.A1(n_912),
.A2(n_923),
.B(n_969),
.C(n_899),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_991),
.A2(n_852),
.B(n_855),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1022),
.A2(n_1024),
.B1(n_1025),
.B2(n_1028),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_940),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1035),
.A2(n_1015),
.B(n_1034),
.C(n_963),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_928),
.A2(n_933),
.B(n_931),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1030),
.B(n_1018),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_940),
.Y(n_1155)
);

AND2x2_ASAP7_75t_SL g1156 ( 
.A(n_945),
.B(n_997),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_999),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_857),
.A2(n_893),
.B(n_873),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_860),
.B(n_1011),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_945),
.B(n_1031),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_945),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_945),
.B(n_987),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_870),
.A2(n_871),
.B(n_878),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_895),
.A2(n_897),
.B(n_900),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_976),
.B(n_1021),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_981),
.B(n_1020),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_SL g1167 ( 
.A(n_970),
.B(n_971),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_942),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_920),
.B(n_924),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_985),
.A2(n_984),
.B(n_888),
.C(n_1010),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1007),
.B(n_892),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_964),
.B(n_950),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_984),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_902),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_903),
.A2(n_906),
.B(n_938),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_989),
.A2(n_947),
.B(n_949),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_982),
.B(n_995),
.Y(n_1177)
);

AO21x1_ASAP7_75t_L g1178 ( 
.A1(n_998),
.A2(n_854),
.B(n_686),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_872),
.A2(n_774),
.B(n_550),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_854),
.B(n_865),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_856),
.Y(n_1181)
);

AO21x1_ASAP7_75t_L g1182 ( 
.A1(n_854),
.A2(n_686),
.B(n_689),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_883),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_858),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_854),
.A2(n_686),
.B(n_711),
.C(n_709),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_879),
.A2(n_888),
.B(n_946),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_854),
.B(n_765),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_854),
.B(n_686),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_883),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_959),
.B(n_694),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_872),
.A2(n_774),
.B(n_550),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_872),
.A2(n_774),
.B(n_550),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_915),
.B(n_686),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1182),
.A2(n_1136),
.A3(n_1178),
.B(n_1132),
.Y(n_1194)
);

AND2x4_ASAP7_75t_L g1195 ( 
.A(n_1190),
.B(n_1126),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1185),
.A2(n_1120),
.B(n_1188),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1187),
.B(n_1189),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1152),
.A2(n_1099),
.B(n_1100),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1100),
.A2(n_1128),
.B(n_1166),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1050),
.B(n_1190),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1193),
.B(n_1180),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1057),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1193),
.B(n_1058),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1069),
.B(n_1073),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1183),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1072),
.A2(n_1173),
.A3(n_1148),
.B(n_1158),
.Y(n_1206)
);

AOI221xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1105),
.A2(n_1054),
.B1(n_1084),
.B2(n_1118),
.C(n_1090),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1062),
.A2(n_1192),
.B(n_1124),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1186),
.A2(n_1125),
.B(n_1111),
.Y(n_1209)
);

NOR2xp67_ASAP7_75t_L g1210 ( 
.A(n_1048),
.B(n_1079),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1133),
.A2(n_1123),
.B(n_1049),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_1038),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1138),
.A2(n_1044),
.B1(n_1117),
.B2(n_1088),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1165),
.A2(n_1172),
.B(n_1055),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_1159),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1156),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1169),
.A2(n_1037),
.B(n_1163),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1181),
.B(n_1081),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1127),
.A2(n_1072),
.B(n_1060),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_1101),
.Y(n_1220)
);

AND2x6_ASAP7_75t_L g1221 ( 
.A(n_1150),
.B(n_1155),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1112),
.A2(n_1102),
.B1(n_1097),
.B2(n_1110),
.Y(n_1222)
);

OA21x2_ASAP7_75t_L g1223 ( 
.A1(n_1186),
.A2(n_1125),
.B(n_1135),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1093),
.A2(n_1090),
.B(n_1109),
.C(n_1118),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1091),
.A2(n_1184),
.B1(n_1094),
.B2(n_1092),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_SL g1226 ( 
.A1(n_1082),
.A2(n_1089),
.B(n_1098),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1043),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1169),
.A2(n_1037),
.B(n_1065),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1046),
.A2(n_1149),
.B(n_1115),
.C(n_1160),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1146),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1175),
.A2(n_1164),
.B(n_1176),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1078),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1095),
.Y(n_1233)
);

AND2x4_ASAP7_75t_L g1234 ( 
.A(n_1114),
.B(n_1143),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1121),
.A2(n_1089),
.B(n_1106),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1052),
.A2(n_1168),
.A3(n_1070),
.B(n_1064),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1147),
.A2(n_1039),
.B(n_1177),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1051),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_SL g1239 ( 
.A(n_1116),
.B(n_1107),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1063),
.B(n_1059),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1063),
.B(n_1085),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_1081),
.B(n_1121),
.Y(n_1242)
);

NOR2xp67_ASAP7_75t_L g1243 ( 
.A(n_1077),
.B(n_1107),
.Y(n_1243)
);

NAND2x1p5_ASAP7_75t_L g1244 ( 
.A(n_1041),
.B(n_1142),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1171),
.A2(n_1170),
.B(n_1036),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1068),
.A2(n_1157),
.B(n_1070),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1047),
.B(n_1040),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_1119),
.B(n_1047),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1040),
.B(n_1154),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1174),
.A2(n_1162),
.B(n_1151),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1066),
.B(n_1041),
.Y(n_1251)
);

AO22x2_ASAP7_75t_L g1252 ( 
.A1(n_1113),
.A2(n_1134),
.B1(n_1056),
.B2(n_1042),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1087),
.A2(n_1080),
.B(n_1131),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1174),
.A2(n_1103),
.B(n_1130),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1043),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1071),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1174),
.A2(n_1067),
.B(n_1139),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1067),
.A2(n_1153),
.B(n_1129),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1045),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1053),
.A2(n_1116),
.B1(n_1096),
.B2(n_1076),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1108),
.B(n_1141),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1137),
.A2(n_1142),
.B1(n_1104),
.B2(n_1075),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1174),
.A2(n_1083),
.B(n_1167),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1161),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1071),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1071),
.B(n_1075),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1075),
.Y(n_1267)
);

OAI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1074),
.A2(n_1145),
.B1(n_1140),
.B2(n_1150),
.C(n_1155),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1144),
.A2(n_1072),
.A3(n_1090),
.B1(n_1089),
.B2(n_1118),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1140),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1140),
.B(n_1155),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1150),
.Y(n_1272)
);

AOI221x1_ASAP7_75t_L g1273 ( 
.A1(n_1144),
.A2(n_854),
.B1(n_1185),
.B2(n_1093),
.C(n_1072),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1144),
.A2(n_728),
.B(n_1152),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1061),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1152),
.A2(n_728),
.B(n_1099),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1185),
.A2(n_854),
.B(n_711),
.C(n_709),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_L g1279 ( 
.A(n_1185),
.B(n_994),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1185),
.A2(n_686),
.B1(n_854),
.B2(n_1188),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1185),
.A2(n_854),
.B(n_711),
.C(n_709),
.Y(n_1281)
);

CKINVDCx11_ASAP7_75t_R g1282 ( 
.A(n_1086),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1122),
.A2(n_1191),
.B(n_1179),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_SL g1284 ( 
.A(n_1185),
.B(n_558),
.C(n_715),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1189),
.Y(n_1285)
);

AO22x2_ASAP7_75t_L g1286 ( 
.A1(n_1072),
.A2(n_1089),
.B1(n_1118),
.B2(n_1090),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1038),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1061),
.Y(n_1288)
);

BUFx5_ASAP7_75t_L g1289 ( 
.A(n_1168),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1290)
);

NOR4xp25_ASAP7_75t_L g1291 ( 
.A(n_1185),
.B(n_854),
.C(n_1084),
.D(n_1106),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1061),
.Y(n_1292)
);

AOI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1079),
.A2(n_716),
.B1(n_715),
.B2(n_875),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1156),
.Y(n_1294)
);

AO32x2_ASAP7_75t_L g1295 ( 
.A1(n_1072),
.A2(n_1090),
.A3(n_1089),
.B1(n_1118),
.B2(n_1070),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1185),
.A2(n_854),
.B(n_686),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1061),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1183),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1101),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1185),
.A2(n_686),
.B1(n_854),
.B2(n_1188),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1038),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1189),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1156),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1305)
);

NAND2x1p5_ASAP7_75t_L g1306 ( 
.A(n_1183),
.B(n_1189),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1187),
.B(n_854),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1185),
.A2(n_854),
.B(n_686),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1061),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1061),
.Y(n_1310)
);

AOI21x1_ASAP7_75t_SL g1311 ( 
.A1(n_1120),
.A2(n_1188),
.B(n_1119),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1182),
.A2(n_1136),
.A3(n_1178),
.B(n_1132),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1185),
.A2(n_854),
.B(n_686),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1185),
.A2(n_854),
.B(n_686),
.Y(n_1315)
);

NOR4xp25_ASAP7_75t_L g1316 ( 
.A(n_1185),
.B(n_854),
.C(n_1084),
.D(n_1106),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1182),
.A2(n_1136),
.A3(n_1178),
.B(n_1132),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1079),
.A2(n_716),
.B1(n_715),
.B2(n_875),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1079),
.A2(n_716),
.B1(n_715),
.B2(n_875),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1185),
.A2(n_686),
.B1(n_854),
.B2(n_1188),
.Y(n_1320)
);

AO31x2_ASAP7_75t_L g1321 ( 
.A1(n_1182),
.A2(n_1136),
.A3(n_1178),
.B(n_1132),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1322)
);

OR2x6_ASAP7_75t_L g1323 ( 
.A(n_1048),
.B(n_883),
.Y(n_1323)
);

A2O1A1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1185),
.A2(n_854),
.B(n_711),
.C(n_709),
.Y(n_1324)
);

AO32x2_ASAP7_75t_L g1325 ( 
.A1(n_1072),
.A2(n_1090),
.A3(n_1089),
.B1(n_1118),
.B2(n_1070),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1152),
.A2(n_728),
.B(n_1099),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1185),
.A2(n_854),
.B(n_686),
.Y(n_1327)
);

NAND2x1p5_ASAP7_75t_L g1328 ( 
.A(n_1183),
.B(n_1189),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1188),
.B(n_874),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1185),
.A2(n_854),
.B(n_711),
.C(n_709),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1188),
.B(n_874),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1185),
.B(n_854),
.C(n_558),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1182),
.A2(n_1136),
.A3(n_1178),
.B(n_1132),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1079),
.A2(n_716),
.B1(n_715),
.B2(n_875),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1188),
.B(n_1187),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1183),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1152),
.A2(n_728),
.B(n_1099),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1183),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1185),
.A2(n_854),
.B(n_711),
.C(n_709),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1185),
.A2(n_854),
.B(n_711),
.C(n_709),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1255),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1205),
.Y(n_1342)
);

BUFx12f_ASAP7_75t_L g1343 ( 
.A(n_1282),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1329),
.B(n_1331),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1307),
.A2(n_1284),
.B1(n_1286),
.B2(n_1332),
.Y(n_1345)
);

BUFx4f_ASAP7_75t_SL g1346 ( 
.A(n_1299),
.Y(n_1346)
);

INVx5_ASAP7_75t_L g1347 ( 
.A(n_1221),
.Y(n_1347)
);

INVx6_ASAP7_75t_L g1348 ( 
.A(n_1255),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_SL g1349 ( 
.A1(n_1286),
.A2(n_1239),
.B1(n_1219),
.B2(n_1290),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1220),
.Y(n_1350)
);

INVx8_ASAP7_75t_L g1351 ( 
.A(n_1221),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1293),
.A2(n_1334),
.B1(n_1318),
.B2(n_1319),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1280),
.A2(n_1320),
.B1(n_1301),
.B2(n_1308),
.Y(n_1353)
);

OAI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1213),
.A2(n_1222),
.B(n_1235),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1296),
.A2(n_1327),
.B1(n_1314),
.B2(n_1315),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1211),
.A2(n_1196),
.B1(n_1305),
.B2(n_1276),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1300),
.A2(n_1335),
.B1(n_1313),
.B2(n_1322),
.Y(n_1357)
);

CKINVDCx11_ASAP7_75t_R g1358 ( 
.A(n_1215),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1242),
.A2(n_1238),
.B1(n_1204),
.B2(n_1200),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1212),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1216),
.B(n_1294),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1201),
.A2(n_1223),
.B1(n_1241),
.B2(n_1252),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1223),
.A2(n_1252),
.B1(n_1248),
.B2(n_1197),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1215),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1260),
.A2(n_1226),
.B1(n_1203),
.B2(n_1237),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1230),
.A2(n_1240),
.B1(n_1279),
.B2(n_1232),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1210),
.A2(n_1330),
.B1(n_1324),
.B2(n_1281),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1287),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1302),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1224),
.A2(n_1278),
.B(n_1339),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1338),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1247),
.B(n_1340),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1275),
.A2(n_1310),
.B1(n_1309),
.B2(n_1292),
.Y(n_1373)
);

AOI22x1_ASAP7_75t_SL g1374 ( 
.A1(n_1264),
.A2(n_1233),
.B1(n_1297),
.B2(n_1288),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1216),
.A2(n_1294),
.B1(n_1304),
.B2(n_1249),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1229),
.A2(n_1218),
.B1(n_1303),
.B2(n_1243),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1225),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1234),
.B(n_1195),
.Y(n_1378)
);

CKINVDCx6p67_ASAP7_75t_R g1379 ( 
.A(n_1323),
.Y(n_1379)
);

INVx1_ASAP7_75t_SL g1380 ( 
.A(n_1202),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1195),
.B(n_1261),
.Y(n_1381)
);

INVx3_ASAP7_75t_SL g1382 ( 
.A(n_1323),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1259),
.A2(n_1207),
.B1(n_1209),
.B2(n_1291),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1306),
.A2(n_1328),
.B1(n_1268),
.B2(n_1262),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_1256),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_1298),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1316),
.B(n_1336),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1267),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1263),
.A2(n_1295),
.B1(n_1325),
.B2(n_1251),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1251),
.B(n_1265),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1270),
.B(n_1227),
.Y(n_1391)
);

BUFx12f_ASAP7_75t_L g1392 ( 
.A(n_1256),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1265),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1266),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1265),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1272),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1271),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1272),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1250),
.A2(n_1274),
.B1(n_1254),
.B2(n_1244),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1258),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1221),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1245),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1209),
.A2(n_1217),
.B1(n_1228),
.B2(n_1199),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1295),
.A2(n_1325),
.B1(n_1214),
.B2(n_1198),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1236),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1246),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1206),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1273),
.B(n_1194),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1194),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1311),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1206),
.Y(n_1411)
);

CKINVDCx14_ASAP7_75t_R g1412 ( 
.A(n_1269),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1253),
.A2(n_1269),
.B1(n_1208),
.B2(n_1257),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1194),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1206),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1312),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1277),
.A2(n_1337),
.B(n_1326),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1283),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1312),
.Y(n_1419)
);

BUFx4f_ASAP7_75t_SL g1420 ( 
.A(n_1333),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1333),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1333),
.Y(n_1422)
);

OAI21xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1231),
.A2(n_1269),
.B(n_1317),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1317),
.B(n_1321),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1317),
.A2(n_1321),
.B1(n_1307),
.B2(n_716),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1321),
.A2(n_1318),
.B1(n_1319),
.B2(n_1293),
.Y(n_1426)
);

INVx1_ASAP7_75t_SL g1427 ( 
.A(n_1285),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1282),
.Y(n_1428)
);

INVx6_ASAP7_75t_L g1429 ( 
.A(n_1255),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1255),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_SL g1431 ( 
.A(n_1205),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1293),
.A2(n_1318),
.B1(n_1319),
.B2(n_1334),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1205),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1281),
.A2(n_854),
.B(n_1185),
.Y(n_1434)
);

CKINVDCx11_ASAP7_75t_R g1435 ( 
.A(n_1282),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1285),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1255),
.Y(n_1437)
);

CKINVDCx6p67_ASAP7_75t_R g1438 ( 
.A(n_1282),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1307),
.A2(n_854),
.B1(n_1284),
.B2(n_1286),
.Y(n_1440)
);

BUFx5_ASAP7_75t_L g1441 ( 
.A(n_1221),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1255),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_SL g1443 ( 
.A1(n_1307),
.A2(n_716),
.B1(n_715),
.B2(n_545),
.Y(n_1443)
);

BUFx10_ASAP7_75t_L g1444 ( 
.A(n_1220),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1307),
.A2(n_854),
.B1(n_1284),
.B2(n_1286),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1282),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1307),
.A2(n_854),
.B1(n_1284),
.B2(n_1286),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1307),
.A2(n_854),
.B1(n_1284),
.B2(n_1286),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1307),
.A2(n_854),
.B1(n_1284),
.B2(n_1286),
.Y(n_1450)
);

BUFx4_ASAP7_75t_R g1451 ( 
.A(n_1215),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1293),
.A2(n_1318),
.B1(n_1319),
.B2(n_1334),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1276),
.B(n_1290),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1285),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1289),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1397),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1350),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1443),
.A2(n_1352),
.B1(n_1432),
.B2(n_1452),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1409),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1403),
.A2(n_1406),
.B(n_1399),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1380),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1416),
.Y(n_1464)
);

NAND2x1p5_ASAP7_75t_L g1465 ( 
.A(n_1402),
.B(n_1347),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_SL g1466 ( 
.A(n_1343),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1405),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1457),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1412),
.B(n_1345),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1419),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_L g1471 ( 
.A(n_1347),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1421),
.Y(n_1472)
);

NAND3xp33_ASAP7_75t_L g1473 ( 
.A(n_1352),
.B(n_1426),
.C(n_1440),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1394),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1422),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1403),
.A2(n_1417),
.B(n_1400),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1411),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1411),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1414),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1415),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1407),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1345),
.B(n_1389),
.Y(n_1482)
);

NAND2x1_ASAP7_75t_L g1483 ( 
.A(n_1365),
.B(n_1353),
.Y(n_1483)
);

INVxp67_ASAP7_75t_L g1484 ( 
.A(n_1436),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1408),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1413),
.A2(n_1434),
.B(n_1367),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1371),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1370),
.B(n_1404),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1387),
.A2(n_1377),
.B(n_1372),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1420),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1420),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1347),
.Y(n_1492)
);

BUFx6f_ASAP7_75t_L g1493 ( 
.A(n_1347),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1423),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1404),
.B(n_1363),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1359),
.A2(n_1374),
.B1(n_1384),
.B2(n_1376),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1439),
.B(n_1446),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1418),
.Y(n_1498)
);

OAI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1354),
.A2(n_1454),
.B1(n_1455),
.B2(n_1453),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1413),
.Y(n_1500)
);

AND2x2_ASAP7_75t_SL g1501 ( 
.A(n_1355),
.B(n_1353),
.Y(n_1501)
);

NAND4xp25_ASAP7_75t_SL g1502 ( 
.A(n_1440),
.B(n_1448),
.C(n_1450),
.D(n_1449),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1355),
.B(n_1425),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1427),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1410),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1383),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1365),
.A2(n_1383),
.B(n_1362),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1348),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1363),
.B(n_1362),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1357),
.A2(n_1448),
.B1(n_1450),
.B2(n_1449),
.Y(n_1510)
);

BUFx12f_ASAP7_75t_L g1511 ( 
.A(n_1435),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1373),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1373),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1356),
.B(n_1344),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1445),
.B(n_1356),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1445),
.B(n_1349),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1410),
.Y(n_1517)
);

INVxp33_ASAP7_75t_L g1518 ( 
.A(n_1378),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1388),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1366),
.B(n_1381),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1441),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1441),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1441),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1366),
.A2(n_1375),
.B(n_1391),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1348),
.Y(n_1525)
);

INVx5_ASAP7_75t_SL g1526 ( 
.A(n_1379),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1392),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1456),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1390),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1361),
.A2(n_1385),
.B(n_1398),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1341),
.B(n_1442),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1386),
.A2(n_1342),
.B(n_1433),
.Y(n_1532)
);

OA21x2_ASAP7_75t_L g1533 ( 
.A1(n_1401),
.A2(n_1451),
.B(n_1351),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1358),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1393),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1431),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1348),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1458),
.B(n_1382),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_1382),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1499),
.B(n_1398),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1460),
.A2(n_1431),
.B1(n_1442),
.B2(n_1341),
.C(n_1437),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1514),
.B(n_1438),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1476),
.A2(n_1396),
.B(n_1395),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1465),
.B(n_1343),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1473),
.B(n_1364),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1459),
.Y(n_1546)
);

A2O1A1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1483),
.A2(n_1430),
.B(n_1360),
.C(n_1368),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1518),
.B(n_1444),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1502),
.A2(n_1428),
.B1(n_1369),
.B2(n_1346),
.Y(n_1549)
);

INVxp33_ASAP7_75t_L g1550 ( 
.A(n_1463),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1483),
.A2(n_1429),
.B(n_1346),
.C(n_1444),
.Y(n_1551)
);

AOI221xp5_ASAP7_75t_L g1552 ( 
.A1(n_1503),
.A2(n_1510),
.B1(n_1482),
.B2(n_1516),
.C(n_1496),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1476),
.A2(n_1428),
.B(n_1447),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1554)
);

NAND2x1p5_ASAP7_75t_L g1555 ( 
.A(n_1533),
.B(n_1471),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_SL g1556 ( 
.A(n_1489),
.B(n_1471),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1501),
.A2(n_1465),
.B(n_1486),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1474),
.B(n_1520),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1516),
.A2(n_1501),
.B1(n_1515),
.B2(n_1488),
.Y(n_1560)
);

A2O1A1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1501),
.A2(n_1486),
.B(n_1503),
.C(n_1515),
.Y(n_1561)
);

OAI211xp5_ASAP7_75t_L g1562 ( 
.A1(n_1482),
.A2(n_1488),
.B(n_1509),
.C(n_1469),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1489),
.B(n_1484),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1481),
.Y(n_1564)
);

AO32x2_ASAP7_75t_L g1565 ( 
.A1(n_1494),
.A2(n_1489),
.A3(n_1508),
.B1(n_1525),
.B2(n_1537),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1481),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1461),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1507),
.A2(n_1532),
.B(n_1465),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1507),
.A2(n_1462),
.B(n_1517),
.Y(n_1569)
);

AO32x2_ASAP7_75t_L g1570 ( 
.A1(n_1494),
.A2(n_1508),
.A3(n_1537),
.B1(n_1525),
.B2(n_1467),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1517),
.B(n_1505),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1505),
.A2(n_1536),
.B1(n_1533),
.B2(n_1479),
.Y(n_1572)
);

OAI211xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1504),
.A2(n_1528),
.B(n_1512),
.C(n_1513),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1523),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1509),
.A2(n_1530),
.B(n_1512),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1485),
.B(n_1495),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1506),
.A2(n_1500),
.B(n_1493),
.C(n_1492),
.Y(n_1577)
);

OA21x2_ASAP7_75t_L g1578 ( 
.A1(n_1464),
.A2(n_1472),
.B(n_1475),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1578),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1563),
.B(n_1498),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1578),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1570),
.B(n_1475),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1570),
.B(n_1470),
.Y(n_1583)
);

AOI222xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1560),
.A2(n_1534),
.B1(n_1470),
.B2(n_1472),
.C1(n_1491),
.C2(n_1490),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1567),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1567),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_L g1587 ( 
.A(n_1552),
.B(n_1490),
.C(n_1491),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1570),
.B(n_1477),
.Y(n_1588)
);

OAI222xp33_ASAP7_75t_L g1589 ( 
.A1(n_1557),
.A2(n_1519),
.B1(n_1466),
.B2(n_1531),
.C1(n_1529),
.C2(n_1498),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1545),
.A2(n_1511),
.B1(n_1524),
.B2(n_1533),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1570),
.B(n_1477),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1564),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1573),
.B(n_1529),
.C(n_1519),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1538),
.Y(n_1594)
);

INVx5_ASAP7_75t_L g1595 ( 
.A(n_1574),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1565),
.B(n_1480),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1566),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1566),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1559),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1546),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1565),
.B(n_1480),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1546),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1576),
.B(n_1468),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1554),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1565),
.B(n_1478),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1575),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1579),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1595),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1593),
.A2(n_1561),
.B1(n_1562),
.B2(n_1590),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1587),
.A2(n_1545),
.B1(n_1541),
.B2(n_1561),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1599),
.B(n_1580),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1580),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1599),
.B(n_1597),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1596),
.B(n_1565),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1594),
.B(n_1550),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_R g1617 ( 
.A(n_1602),
.B(n_1511),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1569),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1601),
.B(n_1606),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1587),
.A2(n_1547),
.B1(n_1568),
.B2(n_1551),
.C(n_1549),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1585),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1585),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1604),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1606),
.B(n_1582),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1581),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1593),
.A2(n_1556),
.B(n_1577),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1586),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1583),
.B(n_1543),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1602),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1608),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1621),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1619),
.B(n_1607),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1618),
.B(n_1605),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1621),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1614),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1613),
.B(n_1607),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1613),
.B(n_1592),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1622),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1622),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1626),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1625),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1628),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1623),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1615),
.B(n_1591),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1612),
.B(n_1603),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1612),
.B(n_1592),
.Y(n_1651)
);

NAND2xp33_ASAP7_75t_SL g1652 ( 
.A(n_1617),
.B(n_1600),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1610),
.B(n_1572),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1604),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1626),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1598),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1633),
.B(n_1618),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1631),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1632),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1632),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1636),
.B(n_1653),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1635),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1635),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1637),
.B(n_1651),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1639),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1655),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1639),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1646),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1650),
.B(n_1616),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1650),
.B(n_1616),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1646),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1641),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1656),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1633),
.B(n_1618),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1656),
.Y(n_1678)
);

OAI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1644),
.A2(n_1611),
.B(n_1610),
.C(n_1627),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1641),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1624),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_SL g1682 ( 
.A(n_1654),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1642),
.B(n_1609),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1633),
.B(n_1629),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1654),
.B(n_1553),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1638),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1640),
.B(n_1629),
.Y(n_1688)
);

NAND2xp67_ASAP7_75t_L g1689 ( 
.A(n_1631),
.B(n_1548),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1638),
.B(n_1624),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1634),
.B(n_1594),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1654),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1643),
.B(n_1623),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_1611),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1654),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1645),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1642),
.B(n_1609),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1693),
.B(n_1642),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1679),
.A2(n_1620),
.B1(n_1663),
.B2(n_1584),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1693),
.B(n_1643),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1667),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1682),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1672),
.B(n_1673),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1666),
.B(n_1644),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1660),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1657),
.B(n_1643),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1683),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1671),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1661),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1666),
.B(n_1645),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1687),
.B(n_1647),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1657),
.B(n_1655),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1662),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1677),
.B(n_1655),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1662),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1676),
.B(n_1647),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1647),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1678),
.B(n_1648),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1674),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1692),
.B(n_1648),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1664),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1660),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1664),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1683),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1695),
.B(n_1648),
.Y(n_1726)
);

NOR2xp67_ASAP7_75t_L g1727 ( 
.A(n_1669),
.B(n_1627),
.Y(n_1727)
);

AND2x4_ASAP7_75t_SL g1728 ( 
.A(n_1683),
.B(n_1544),
.Y(n_1728)
);

NOR2x1_ASAP7_75t_SL g1729 ( 
.A(n_1694),
.B(n_1544),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1685),
.B(n_1649),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1691),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1649),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1669),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1720),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1699),
.A2(n_1620),
.B(n_1630),
.C(n_1547),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1699),
.B(n_1689),
.Y(n_1736)
);

NAND3xp33_ASAP7_75t_L g1737 ( 
.A(n_1701),
.B(n_1584),
.C(n_1665),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1705),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1702),
.A2(n_1590),
.B1(n_1630),
.B2(n_1685),
.Y(n_1739)
);

OAI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1702),
.A2(n_1659),
.B1(n_1690),
.B2(n_1681),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1725),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1709),
.B(n_1689),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1709),
.Y(n_1743)
);

NOR3xp33_ASAP7_75t_L g1744 ( 
.A(n_1703),
.B(n_1539),
.C(n_1542),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1703),
.B(n_1659),
.Y(n_1745)
);

INVxp67_ASAP7_75t_SL g1746 ( 
.A(n_1727),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_L g1747 ( 
.A(n_1701),
.B(n_1669),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1705),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1701),
.Y(n_1749)
);

NAND4xp25_ASAP7_75t_L g1750 ( 
.A(n_1727),
.B(n_1551),
.C(n_1571),
.D(n_1540),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1729),
.B(n_1684),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1731),
.B(n_1690),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1712),
.B(n_1684),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1704),
.A2(n_1617),
.B(n_1571),
.C(n_1589),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1728),
.A2(n_1685),
.B1(n_1553),
.B2(n_1544),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1704),
.B(n_1589),
.C(n_1459),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1729),
.A2(n_1600),
.B(n_1625),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1712),
.B(n_1681),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1721),
.B(n_1688),
.Y(n_1759)
);

O2A1O1Ixp33_ASAP7_75t_L g1760 ( 
.A1(n_1735),
.A2(n_1708),
.B(n_1725),
.C(n_1714),
.Y(n_1760)
);

INVxp67_ASAP7_75t_SL g1761 ( 
.A(n_1734),
.Y(n_1761)
);

INVxp67_ASAP7_75t_L g1762 ( 
.A(n_1749),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1743),
.B(n_1718),
.Y(n_1763)
);

AOI222xp33_ASAP7_75t_L g1764 ( 
.A1(n_1736),
.A2(n_1719),
.B1(n_1717),
.B2(n_1726),
.C1(n_1721),
.C2(n_1730),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1752),
.A2(n_1728),
.B(n_1708),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1754),
.A2(n_1728),
.B1(n_1717),
.B2(n_1719),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1757),
.A2(n_1708),
.B(n_1733),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1738),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1748),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1737),
.A2(n_1718),
.B1(n_1732),
.B2(n_1700),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1741),
.Y(n_1771)
);

OAI31xp33_ASAP7_75t_L g1772 ( 
.A1(n_1739),
.A2(n_1730),
.A3(n_1698),
.B(n_1726),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1740),
.B(n_1718),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1747),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1745),
.Y(n_1775)
);

AOI32xp33_ASAP7_75t_L g1776 ( 
.A1(n_1756),
.A2(n_1698),
.A3(n_1713),
.B1(n_1715),
.B2(n_1700),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1756),
.A2(n_1553),
.B1(n_1722),
.B2(n_1716),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1742),
.A2(n_1733),
.B(n_1714),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1751),
.Y(n_1779)
);

INVxp67_ASAP7_75t_L g1780 ( 
.A(n_1761),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1761),
.Y(n_1781)
);

NOR3x1_ASAP7_75t_L g1782 ( 
.A(n_1763),
.B(n_1773),
.C(n_1775),
.Y(n_1782)
);

AOI211x1_ASAP7_75t_L g1783 ( 
.A1(n_1765),
.A2(n_1758),
.B(n_1750),
.C(n_1753),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1762),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1762),
.Y(n_1785)
);

AND3x1_ASAP7_75t_L g1786 ( 
.A(n_1760),
.B(n_1755),
.C(n_1744),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1771),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1764),
.B(n_1744),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1759),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1768),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1770),
.B(n_1711),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1784),
.B(n_1785),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_L g1793 ( 
.A(n_1780),
.B(n_1772),
.C(n_1774),
.Y(n_1793)
);

AOI221xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1788),
.A2(n_1766),
.B1(n_1777),
.B2(n_1767),
.C(n_1778),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1781),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1787),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1791),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1790),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1789),
.B(n_1769),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1782),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1788),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1794),
.B(n_1786),
.C(n_1783),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1797),
.Y(n_1803)
);

O2A1O1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1800),
.A2(n_1801),
.B(n_1793),
.C(n_1799),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1800),
.A2(n_1799),
.B1(n_1792),
.B2(n_1795),
.C(n_1777),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1792),
.A2(n_1776),
.B1(n_1746),
.B2(n_1710),
.C(n_1724),
.Y(n_1806)
);

OA211x2_ASAP7_75t_L g1807 ( 
.A1(n_1805),
.A2(n_1746),
.B(n_1796),
.C(n_1798),
.Y(n_1807)
);

AOI211xp5_ASAP7_75t_L g1808 ( 
.A1(n_1802),
.A2(n_1710),
.B(n_1724),
.C(n_1716),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1803),
.A2(n_1698),
.B1(n_1722),
.B2(n_1715),
.Y(n_1809)
);

OAI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1804),
.A2(n_1711),
.B1(n_1715),
.B2(n_1713),
.Y(n_1810)
);

OAI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1806),
.A2(n_1723),
.B(n_1706),
.C(n_1527),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1803),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1812),
.Y(n_1813)
);

AO22x1_ASAP7_75t_L g1814 ( 
.A1(n_1810),
.A2(n_1713),
.B1(n_1683),
.B2(n_1697),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1809),
.B(n_1707),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1807),
.Y(n_1816)
);

NAND4xp75_ASAP7_75t_L g1817 ( 
.A(n_1811),
.B(n_1723),
.C(n_1706),
.D(n_1732),
.Y(n_1817)
);

OAI221xp5_ASAP7_75t_L g1818 ( 
.A1(n_1813),
.A2(n_1808),
.B1(n_1706),
.B2(n_1723),
.C(n_1669),
.Y(n_1818)
);

NOR4xp25_ASAP7_75t_L g1819 ( 
.A(n_1816),
.B(n_1686),
.C(n_1660),
.D(n_1696),
.Y(n_1819)
);

OAI31xp33_ASAP7_75t_L g1820 ( 
.A1(n_1815),
.A2(n_1686),
.A3(n_1697),
.B(n_1535),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1818),
.Y(n_1821)
);

NAND5xp2_ASAP7_75t_L g1822 ( 
.A(n_1821),
.B(n_1820),
.C(n_1817),
.D(n_1819),
.E(n_1814),
.Y(n_1822)
);

INVx4_ASAP7_75t_L g1823 ( 
.A(n_1822),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1822),
.Y(n_1824)
);

OA22x2_ASAP7_75t_L g1825 ( 
.A1(n_1823),
.A2(n_1686),
.B1(n_1697),
.B2(n_1665),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1824),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1826),
.A2(n_1686),
.B1(n_1675),
.B2(n_1696),
.C(n_1680),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1825),
.Y(n_1828)
);

AOI322xp5_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1732),
.A3(n_1707),
.B1(n_1697),
.B2(n_1668),
.C1(n_1680),
.C2(n_1675),
.Y(n_1829)
);

AO21x2_ASAP7_75t_L g1830 ( 
.A1(n_1829),
.A2(n_1827),
.B(n_1658),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1830),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_R g1832 ( 
.A1(n_1831),
.A2(n_1526),
.B1(n_1658),
.B2(n_1670),
.C(n_1668),
.Y(n_1832)
);

AOI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1832),
.A2(n_1535),
.B(n_1527),
.C(n_1487),
.Y(n_1833)
);


endmodule