module fake_jpeg_28170_n_237 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_237);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx2_ASAP7_75t_R g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_20),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_17),
.B1(n_18),
.B2(n_24),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_17),
.B1(n_24),
.B2(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_49),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_33),
.B1(n_32),
.B2(n_34),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_33),
.A2(n_24),
.B1(n_18),
.B2(n_22),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_27),
.B(n_25),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_20),
.B1(n_16),
.B2(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_48),
.A2(n_20),
.B1(n_16),
.B2(n_19),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_35),
.B1(n_34),
.B2(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_50),
.B(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_56),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_48),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx11_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_65),
.B1(n_27),
.B2(n_23),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_14),
.B1(n_19),
.B2(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_43),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_43),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_81),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_49),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_68),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_43),
.C(n_47),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_43),
.B1(n_35),
.B2(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_70),
.A2(n_43),
.B1(n_35),
.B2(n_39),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_71),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_31),
.C(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_98),
.B(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_104),
.B(n_92),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_87),
.B(n_74),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_108),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_52),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_112),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_36),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_28),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_114),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_14),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_59),
.B1(n_27),
.B2(n_23),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_118),
.A2(n_95),
.B1(n_23),
.B2(n_25),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_83),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_31),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_31),
.Y(n_145)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_123),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_80),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_124),
.B(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_135),
.B1(n_144),
.B2(n_114),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_13),
.B(n_15),
.C(n_97),
.D(n_77),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_SL g156 ( 
.A(n_131),
.B(n_133),
.C(n_140),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_26),
.B1(n_25),
.B2(n_97),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_111),
.A2(n_59),
.B1(n_97),
.B2(n_92),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_136),
.A2(n_61),
.B1(n_73),
.B2(n_2),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_15),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_86),
.B1(n_31),
.B2(n_15),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_138),
.A2(n_142),
.B1(n_110),
.B2(n_105),
.Y(n_159)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_117),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_13),
.B1(n_15),
.B2(n_10),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_148),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_99),
.A2(n_31),
.B1(n_62),
.B2(n_56),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_31),
.B1(n_11),
.B2(n_10),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_145),
.A2(n_123),
.B1(n_106),
.B2(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_133),
.A2(n_102),
.B(n_121),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_165),
.B(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_152),
.A2(n_166),
.B1(n_140),
.B2(n_128),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_163),
.Y(n_179)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_100),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_155),
.A2(n_132),
.B(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_157),
.B(n_158),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_127),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_138),
.B1(n_146),
.B2(n_61),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_101),
.Y(n_160)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_101),
.C(n_100),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_167),
.C(n_169),
.Y(n_184)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_147),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_120),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_136),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_109),
.B(n_115),
.Y(n_165)
);

OAI21x1_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_118),
.B(n_11),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_107),
.C(n_73),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_107),
.C(n_73),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_107),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_125),
.B1(n_147),
.B2(n_134),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_143),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_175),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_177),
.B(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_130),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_185),
.B(n_171),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_186),
.A2(n_154),
.B1(n_159),
.B2(n_164),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_190),
.A2(n_193),
.B1(n_178),
.B2(n_182),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_195),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_155),
.B1(n_150),
.B2(n_156),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_168),
.B(n_165),
.C(n_156),
.D(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_196),
.B(n_172),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_167),
.C(n_153),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_184),
.C(n_173),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_177),
.B(n_174),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_11),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_179),
.B1(n_185),
.B2(n_183),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_204),
.B1(n_200),
.B2(n_210),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_179),
.B1(n_181),
.B2(n_172),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_162),
.C(n_8),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_8),
.Y(n_219)
);

OA21x2_ASAP7_75t_SL g212 ( 
.A1(n_208),
.A2(n_195),
.B(n_191),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_217),
.B(n_207),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_202),
.B1(n_204),
.B2(n_201),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_209),
.A2(n_193),
.B(n_188),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_219),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_191),
.B(n_162),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_214),
.A2(n_206),
.B1(n_211),
.B2(n_205),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_224),
.C(n_225),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_206),
.B(n_1),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_223),
.B(n_215),
.C(n_216),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_228),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_217),
.B(n_1),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_0),
.B(n_2),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_230),
.A2(n_232),
.B1(n_4),
.B2(n_5),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_223),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_234),
.B(n_3),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_235),
.A2(n_4),
.B(n_5),
.Y(n_236)
);

XNOR2x2_ASAP7_75t_SL g237 ( 
.A(n_236),
.B(n_6),
.Y(n_237)
);


endmodule