module real_aes_6818_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_725;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g535 ( .A1(n_0), .A2(n_181), .B(n_536), .C(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_1), .B(n_486), .Y(n_540) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g193 ( .A(n_3), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_4), .B(n_153), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_5), .A2(n_459), .B(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_6), .A2(n_173), .B(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_7), .A2(n_35), .B1(n_147), .B2(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_8), .B(n_173), .Y(n_182) );
AND2x6_ASAP7_75t_L g165 ( .A(n_9), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_10), .A2(n_165), .B(n_464), .C(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_11), .B(n_36), .Y(n_126) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
INVx1_ASAP7_75t_L g186 ( .A(n_13), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_14), .B(n_151), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_15), .B(n_153), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_16), .B(n_139), .Y(n_257) );
AO32x2_ASAP7_75t_L g199 ( .A1(n_17), .A2(n_138), .A3(n_164), .B1(n_173), .B2(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_18), .B(n_147), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_19), .B(n_139), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_51), .B1(n_147), .B2(n_202), .Y(n_203) );
AOI22xp33_ASAP7_75t_SL g241 ( .A1(n_21), .A2(n_78), .B1(n_147), .B2(n_151), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_22), .B(n_147), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_23), .A2(n_164), .B(n_464), .C(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_24), .A2(n_56), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_24), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_25), .A2(n_164), .B(n_464), .C(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_26), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_27), .B(n_168), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_28), .A2(n_459), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_29), .B(n_168), .Y(n_216) );
INVx2_ASAP7_75t_L g149 ( .A(n_30), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_31), .A2(n_462), .B(n_472), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_32), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_33), .B(n_168), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_34), .B(n_223), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_36), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_37), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_38), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_39), .B(n_153), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_40), .B(n_459), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_41), .A2(n_101), .B1(n_114), .B2(n_757), .Y(n_100) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_42), .A2(n_462), .B(n_466), .C(n_472), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_43), .B(n_147), .Y(n_176) );
INVx1_ASAP7_75t_L g537 ( .A(n_44), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_45), .A2(n_89), .B1(n_202), .B2(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g467 ( .A(n_46), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_47), .B(n_147), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_48), .B(n_147), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_49), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_50), .B(n_159), .Y(n_180) );
AOI22xp33_ASAP7_75t_SL g255 ( .A1(n_52), .A2(n_57), .B1(n_147), .B2(n_151), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_53), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_54), .B(n_147), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_55), .B(n_147), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_56), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g447 ( .A1(n_56), .A2(n_130), .B1(n_131), .B2(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_58), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g166 ( .A(n_59), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_60), .B(n_459), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_61), .B(n_486), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_62), .A2(n_159), .B(n_189), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_63), .B(n_147), .Y(n_194) );
INVx1_ASAP7_75t_L g142 ( .A(n_64), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_66), .B(n_153), .Y(n_504) );
AO32x2_ASAP7_75t_L g237 ( .A1(n_67), .A2(n_164), .A3(n_173), .B1(n_238), .B2(n_242), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_68), .B(n_154), .Y(n_550) );
INVx1_ASAP7_75t_L g157 ( .A(n_69), .Y(n_157) );
INVx1_ASAP7_75t_L g211 ( .A(n_70), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_71), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_72), .B(n_469), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_73), .A2(n_464), .B(n_472), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_74), .B(n_151), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_75), .Y(n_481) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_77), .B(n_468), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g442 ( .A1(n_79), .A2(n_83), .B1(n_443), .B2(n_750), .C1(n_755), .C2(n_756), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_80), .B(n_202), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_81), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_82), .B(n_151), .Y(n_215) );
INVx1_ASAP7_75t_L g755 ( .A(n_83), .Y(n_755) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_85), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_86), .B(n_163), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_87), .B(n_151), .Y(n_177) );
INVx2_ASAP7_75t_L g110 ( .A(n_88), .Y(n_110) );
OR2x2_ASAP7_75t_L g123 ( .A(n_88), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g446 ( .A(n_88), .B(n_125), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_90), .A2(n_99), .B1(n_151), .B2(n_152), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_91), .B(n_459), .Y(n_500) );
INVx1_ASAP7_75t_L g503 ( .A(n_92), .Y(n_503) );
INVxp67_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_94), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_95), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g525 ( .A(n_96), .Y(n_525) );
INVx1_ASAP7_75t_L g546 ( .A(n_97), .Y(n_546) );
AND2x2_ASAP7_75t_L g474 ( .A(n_98), .B(n_168), .Y(n_474) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx3_ASAP7_75t_SL g759 ( .A(n_103), .Y(n_759) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .C(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g125 ( .A(n_109), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g451 ( .A(n_110), .B(n_125), .Y(n_451) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_110), .B(n_124), .Y(n_756) );
OA211x2_ASAP7_75t_L g114 ( .A1(n_111), .A2(n_115), .B(n_120), .C(n_439), .Y(n_114) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g441 ( .A(n_117), .Y(n_441) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_127), .B(n_435), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g438 ( .A(n_123), .Y(n_438) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_131), .Y(n_127) );
INVx1_ASAP7_75t_SL g448 ( .A(n_131), .Y(n_448) );
OR3x1_ASAP7_75t_L g131 ( .A(n_132), .B(n_363), .C(n_412), .Y(n_131) );
NAND5xp2_ASAP7_75t_L g132 ( .A(n_133), .B(n_278), .C(n_306), .D(n_336), .E(n_350), .Y(n_132) );
AOI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_196), .B1(n_228), .B2(n_233), .C(n_244), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_169), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_135), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g258 ( .A(n_136), .Y(n_258) );
AND2x2_ASAP7_75t_L g266 ( .A(n_136), .B(n_172), .Y(n_266) );
AND2x2_ASAP7_75t_L g289 ( .A(n_136), .B(n_171), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_136), .B(n_183), .Y(n_304) );
OR2x2_ASAP7_75t_L g313 ( .A(n_136), .B(n_251), .Y(n_313) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_136), .Y(n_316) );
AND2x2_ASAP7_75t_L g424 ( .A(n_136), .B(n_251), .Y(n_424) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_144), .B(n_167), .Y(n_136) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_137), .A2(n_184), .B(n_195), .Y(n_183) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_138), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_140), .B(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_156), .B(n_164), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_150), .B(n_153), .Y(n_145) );
INVx3_ASAP7_75t_L g210 ( .A(n_147), .Y(n_210) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_147), .Y(n_527) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
BUFx3_ASAP7_75t_L g240 ( .A(n_148), .Y(n_240) );
AND2x6_ASAP7_75t_L g464 ( .A(n_148), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g152 ( .A(n_149), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_149), .Y(n_160) );
INVx2_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_153), .A2(n_176), .B(n_177), .Y(n_175) );
INVx2_ASAP7_75t_L g181 ( .A(n_153), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_SL g209 ( .A1(n_153), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_153), .B(n_484), .Y(n_483) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_SL g238 ( .A1(n_154), .A2(n_163), .B1(n_239), .B2(n_241), .Y(n_238) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
INVx1_ASAP7_75t_L g223 ( .A(n_155), .Y(n_223) );
AND2x2_ASAP7_75t_L g460 ( .A(n_155), .B(n_160), .Y(n_460) );
INVx1_ASAP7_75t_L g465 ( .A(n_155), .Y(n_465) );
O2A1O1Ixp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_161), .C(n_162), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_158), .A2(n_181), .B(n_193), .C(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_158), .A2(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_162), .A2(n_225), .B(n_226), .Y(n_224) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_163), .A2(n_181), .B1(n_201), .B2(n_203), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_163), .A2(n_181), .B1(n_254), .B2(n_255), .Y(n_253) );
INVx4_ASAP7_75t_L g538 ( .A(n_163), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g277 ( .A(n_164), .B(n_252), .C(n_253), .Y(n_277) );
BUFx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_165), .A2(n_175), .B(n_178), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g184 ( .A1(n_165), .A2(n_185), .B(n_192), .Y(n_184) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_165), .A2(n_209), .B(n_213), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g218 ( .A1(n_165), .A2(n_219), .B(n_224), .Y(n_218) );
AND2x4_ASAP7_75t_L g459 ( .A(n_165), .B(n_460), .Y(n_459) );
INVx4_ASAP7_75t_SL g473 ( .A(n_165), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_165), .B(n_460), .Y(n_547) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_168), .A2(n_208), .B(n_216), .Y(n_207) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_168), .A2(n_218), .B(n_227), .Y(n_217) );
INVx2_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_168), .A2(n_458), .B(n_461), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_168), .A2(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g519 ( .A(n_168), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_169), .B(n_316), .Y(n_372) );
INVx2_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
OAI311xp33_ASAP7_75t_L g314 ( .A1(n_170), .A2(n_315), .A3(n_316), .B1(n_317), .C1(n_332), .Y(n_314) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_183), .Y(n_170) );
AND2x2_ASAP7_75t_L g275 ( .A(n_171), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g282 ( .A(n_171), .Y(n_282) );
AND2x2_ASAP7_75t_L g403 ( .A(n_171), .B(n_232), .Y(n_403) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_172), .B(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g259 ( .A(n_172), .B(n_183), .Y(n_259) );
AND2x2_ASAP7_75t_L g311 ( .A(n_172), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g325 ( .A(n_172), .B(n_258), .Y(n_325) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_182), .Y(n_172) );
INVx4_ASAP7_75t_L g252 ( .A(n_173), .Y(n_252) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_173), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_173), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B(n_181), .Y(n_178) );
INVx2_ASAP7_75t_L g232 ( .A(n_183), .Y(n_232) );
AND2x2_ASAP7_75t_L g274 ( .A(n_183), .B(n_258), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_188), .C(n_189), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_187), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_187), .A2(n_550), .B(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_189), .A2(n_525), .B(n_526), .C(n_527), .Y(n_524) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_190), .A2(n_214), .B(n_215), .Y(n_213) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g469 ( .A(n_191), .Y(n_469) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_204), .Y(n_196) );
OR2x2_ASAP7_75t_L g369 ( .A(n_197), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_197), .B(n_375), .Y(n_386) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_198), .B(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g243 ( .A(n_199), .Y(n_243) );
AND2x2_ASAP7_75t_L g310 ( .A(n_199), .B(n_237), .Y(n_310) );
AND2x2_ASAP7_75t_L g321 ( .A(n_199), .B(n_217), .Y(n_321) );
AND2x2_ASAP7_75t_L g330 ( .A(n_199), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_204), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_204), .B(n_271), .Y(n_315) );
INVx2_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g302 ( .A(n_205), .B(n_261), .Y(n_302) );
OR2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_217), .Y(n_205) );
INVx2_ASAP7_75t_L g235 ( .A(n_206), .Y(n_235) );
AND2x2_ASAP7_75t_L g329 ( .A(n_206), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
OR2x2_ASAP7_75t_L g346 ( .A(n_207), .B(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_207), .Y(n_409) );
AND2x2_ASAP7_75t_L g248 ( .A(n_217), .B(n_243), .Y(n_248) );
INVx1_ASAP7_75t_L g269 ( .A(n_217), .Y(n_269) );
AND2x2_ASAP7_75t_L g290 ( .A(n_217), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g331 ( .A(n_217), .Y(n_331) );
INVx1_ASAP7_75t_L g347 ( .A(n_217), .Y(n_347) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_217), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_230), .B(n_335), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_230), .A2(n_320), .B1(n_369), .B2(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OAI211xp5_ASAP7_75t_SL g412 ( .A1(n_231), .A2(n_413), .B(n_415), .C(n_433), .Y(n_412) );
INVx2_ASAP7_75t_L g265 ( .A(n_232), .Y(n_265) );
AND2x2_ASAP7_75t_L g323 ( .A(n_232), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g334 ( .A(n_232), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_233), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g307 ( .A(n_234), .B(n_271), .Y(n_307) );
BUFx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g339 ( .A(n_235), .B(n_330), .Y(n_339) );
AND2x2_ASAP7_75t_L g358 ( .A(n_235), .B(n_272), .Y(n_358) );
AND2x4_ASAP7_75t_L g294 ( .A(n_236), .B(n_268), .Y(n_294) );
AND2x2_ASAP7_75t_L g432 ( .A(n_236), .B(n_408), .Y(n_432) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_237), .Y(n_261) );
INVx1_ASAP7_75t_L g272 ( .A(n_237), .Y(n_272) );
INVx1_ASAP7_75t_L g371 ( .A(n_237), .Y(n_371) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_240), .Y(n_471) );
INVx2_ASAP7_75t_L g539 ( .A(n_240), .Y(n_539) );
INVx1_ASAP7_75t_L g516 ( .A(n_242), .Y(n_516) );
OR2x2_ASAP7_75t_L g262 ( .A(n_243), .B(n_247), .Y(n_262) );
AND2x2_ASAP7_75t_L g271 ( .A(n_243), .B(n_272), .Y(n_271) );
NOR2xp67_ASAP7_75t_L g291 ( .A(n_243), .B(n_292), .Y(n_291) );
OAI221xp5_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_249), .B1(n_260), .B2(n_263), .C(n_267), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_246), .A2(n_268), .B(n_270), .C(n_273), .Y(n_267) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g292 ( .A(n_247), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_247), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_247), .B(n_269), .Y(n_375) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_247), .Y(n_382) );
AND2x2_ASAP7_75t_L g300 ( .A(n_248), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g337 ( .A(n_248), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_259), .Y(n_249) );
INVx2_ASAP7_75t_L g328 ( .A(n_250), .Y(n_328) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_250), .A2(n_261), .B1(n_378), .B2(n_380), .C1(n_381), .C2(n_383), .Y(n_377) );
AND2x2_ASAP7_75t_L g434 ( .A(n_250), .B(n_403), .Y(n_434) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_258), .Y(n_250) );
INVx1_ASAP7_75t_L g324 ( .A(n_251), .Y(n_324) );
AO21x1_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B(n_256), .Y(n_251) );
INVx3_ASAP7_75t_L g486 ( .A(n_252), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_252), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_252), .A2(n_522), .B(n_529), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_252), .B(n_530), .Y(n_529) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_252), .A2(n_545), .B(n_552), .Y(n_544) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x4_ASAP7_75t_L g276 ( .A(n_257), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g362 ( .A(n_259), .B(n_296), .Y(n_362) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_260), .A2(n_374), .B(n_376), .Y(n_373) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_261), .B(n_268), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_261), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx3_ASAP7_75t_L g327 ( .A(n_265), .Y(n_327) );
OR2x2_ASAP7_75t_L g379 ( .A(n_265), .B(n_301), .Y(n_379) );
AND2x2_ASAP7_75t_L g295 ( .A(n_266), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g333 ( .A(n_266), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_266), .B(n_327), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_266), .B(n_323), .Y(n_349) );
AND2x2_ASAP7_75t_L g353 ( .A(n_266), .B(n_335), .Y(n_353) );
INVxp67_ASAP7_75t_L g285 ( .A(n_268), .Y(n_285) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_270), .A2(n_343), .B1(n_348), .B2(n_349), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_270), .B(n_375), .Y(n_405) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g391 ( .A(n_271), .B(n_382), .Y(n_391) );
AND2x2_ASAP7_75t_L g420 ( .A(n_271), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g425 ( .A(n_271), .B(n_375), .Y(n_425) );
INVx1_ASAP7_75t_L g338 ( .A(n_272), .Y(n_338) );
BUFx2_ASAP7_75t_L g344 ( .A(n_272), .Y(n_344) );
INVx1_ASAP7_75t_L g429 ( .A(n_273), .Y(n_429) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2x1p5_ASAP7_75t_L g280 ( .A(n_274), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g305 ( .A(n_275), .Y(n_305) );
NOR2x1_ASAP7_75t_L g281 ( .A(n_276), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g288 ( .A(n_276), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx3_ASAP7_75t_L g335 ( .A(n_276), .Y(n_335) );
OR2x2_ASAP7_75t_L g401 ( .A(n_276), .B(n_402), .Y(n_401) );
AOI211xp5_ASAP7_75t_L g278 ( .A1(n_279), .A2(n_283), .B(n_286), .C(n_298), .Y(n_278) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_279), .A2(n_416), .B1(n_423), .B2(n_425), .C(n_426), .Y(n_415) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_287), .B(n_293), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_289), .B(n_327), .Y(n_341) );
AND2x2_ASAP7_75t_L g383 ( .A(n_289), .B(n_323), .Y(n_383) );
INVx1_ASAP7_75t_SL g396 ( .A(n_290), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_290), .B(n_344), .Y(n_399) );
INVx1_ASAP7_75t_L g417 ( .A(n_291), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_295), .A2(n_385), .B1(n_387), .B2(n_391), .C(n_392), .Y(n_384) );
AND2x2_ASAP7_75t_L g411 ( .A(n_296), .B(n_403), .Y(n_411) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g395 ( .A(n_297), .Y(n_395) );
AOI21xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_302), .B(n_303), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g366 ( .A(n_301), .B(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g352 ( .A(n_302), .Y(n_352) );
INVx1_ASAP7_75t_L g380 ( .A(n_303), .Y(n_380) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_311), .C(n_314), .Y(n_306) );
OAI31xp33_ASAP7_75t_L g433 ( .A1(n_307), .A2(n_345), .A3(n_432), .B(n_434), .Y(n_433) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g407 ( .A(n_310), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g428 ( .A(n_310), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_312), .B(n_327), .Y(n_355) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g430 ( .A(n_313), .B(n_327), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_322), .B1(n_326), .B2(n_329), .Y(n_317) );
NAND2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_321), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g357 ( .A(n_321), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g360 ( .A(n_321), .B(n_344), .Y(n_360) );
AND2x2_ASAP7_75t_L g414 ( .A(n_321), .B(n_409), .Y(n_414) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx1_ASAP7_75t_L g389 ( .A(n_325), .Y(n_389) );
NOR2xp67_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
OAI32xp33_ASAP7_75t_L g392 ( .A1(n_327), .A2(n_361), .A3(n_393), .B1(n_395), .B2(n_396), .Y(n_392) );
INVx1_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_330), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g390 ( .A(n_334), .Y(n_390) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B(n_340), .C(n_342), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_338), .B(n_375), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_339), .A2(n_351), .B1(n_352), .B2(n_353), .C(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g351 ( .A(n_349), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_359), .B2(n_361), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND4xp25_ASAP7_75t_SL g416 ( .A(n_359), .B(n_417), .C(n_418), .D(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
NAND4xp25_ASAP7_75t_SL g363 ( .A(n_364), .B(n_377), .C(n_384), .D(n_397), .Y(n_363) );
O2A1O1Ixp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B(n_372), .C(n_373), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_SL g394 ( .A(n_370), .Y(n_394) );
INVx2_ASAP7_75t_L g418 ( .A(n_375), .Y(n_418) );
OR2x2_ASAP7_75t_L g427 ( .A(n_382), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_404), .Y(n_397) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g423 ( .A(n_403), .B(n_424), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_406), .B(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
CKINVDCx16_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_426) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND3xp33_ASAP7_75t_SL g439 ( .A(n_435), .B(n_440), .C(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_447), .B1(n_449), .B2(n_452), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g751 ( .A(n_445), .Y(n_751) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g752 ( .A(n_447), .Y(n_752) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g753 ( .A(n_450), .Y(n_753) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx4_ASAP7_75t_L g754 ( .A(n_452), .Y(n_754) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR5x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_623), .C(n_701), .D(n_725), .E(n_742), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_495), .B(n_541), .C(n_600), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_475), .Y(n_455) );
AND2x2_ASAP7_75t_L g554 ( .A(n_456), .B(n_477), .Y(n_554) );
INVx5_ASAP7_75t_SL g582 ( .A(n_456), .Y(n_582) );
AND2x2_ASAP7_75t_L g618 ( .A(n_456), .B(n_603), .Y(n_618) );
OR2x2_ASAP7_75t_L g657 ( .A(n_456), .B(n_476), .Y(n_657) );
OR2x2_ASAP7_75t_L g688 ( .A(n_456), .B(n_579), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_456), .B(n_592), .Y(n_724) );
AND2x2_ASAP7_75t_L g736 ( .A(n_456), .B(n_579), .Y(n_736) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_474), .Y(n_456) );
BUFx2_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_463), .A2(n_473), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_463), .A2(n_473), .B(n_534), .C(n_535), .Y(n_533) );
INVx5_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .C(n_471), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_468), .A2(n_471), .B(n_503), .C(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g735 ( .A(n_475), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g598 ( .A(n_476), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_477), .B(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_477), .Y(n_591) );
INVx3_ASAP7_75t_L g606 ( .A(n_477), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_477), .B(n_487), .Y(n_630) );
OR2x2_ASAP7_75t_L g639 ( .A(n_477), .B(n_582), .Y(n_639) );
AND2x2_ASAP7_75t_L g643 ( .A(n_477), .B(n_603), .Y(n_643) );
AND2x2_ASAP7_75t_L g649 ( .A(n_477), .B(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g686 ( .A(n_477), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_477), .B(n_544), .Y(n_700) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_486), .A2(n_532), .B(n_540), .Y(n_531) );
OR2x2_ASAP7_75t_L g592 ( .A(n_487), .B(n_544), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_487), .B(n_579), .Y(n_603) );
AND2x2_ASAP7_75t_L g615 ( .A(n_487), .B(n_606), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_487), .B(n_544), .Y(n_638) );
INVx1_ASAP7_75t_SL g650 ( .A(n_487), .Y(n_650) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g543 ( .A(n_488), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_488), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
AND2x2_ASAP7_75t_L g563 ( .A(n_497), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_497), .B(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g570 ( .A(n_497), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_497), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g595 ( .A(n_497), .B(n_586), .Y(n_595) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_497), .Y(n_614) );
AND2x2_ASAP7_75t_L g635 ( .A(n_497), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g645 ( .A(n_497), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g691 ( .A(n_497), .B(n_574), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_497), .B(n_597), .Y(n_718) );
INVx5_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g588 ( .A(n_498), .Y(n_588) );
AND2x2_ASAP7_75t_L g654 ( .A(n_498), .B(n_586), .Y(n_654) );
AND2x2_ASAP7_75t_L g738 ( .A(n_498), .B(n_606), .Y(n_738) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_507), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_507), .Y(n_727) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
AND2x2_ASAP7_75t_L g557 ( .A(n_508), .B(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g566 ( .A(n_508), .B(n_564), .Y(n_566) );
INVx5_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
AND2x2_ASAP7_75t_L g597 ( .A(n_508), .B(n_531), .Y(n_597) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_508), .Y(n_634) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_512), .B(n_516), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g675 ( .A(n_520), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_520), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g708 ( .A(n_520), .B(n_574), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_520), .A2(n_631), .B(n_738), .C(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
BUFx2_ASAP7_75t_L g558 ( .A(n_521), .Y(n_558) );
INVx2_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .Y(n_522) );
INVx2_ASAP7_75t_L g564 ( .A(n_531), .Y(n_564) );
AND2x2_ASAP7_75t_L g571 ( .A(n_531), .B(n_562), .Y(n_571) );
AND2x2_ASAP7_75t_L g662 ( .A(n_531), .B(n_574), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AOI211x1_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_555), .B(n_568), .C(n_593), .Y(n_541) );
INVx1_ASAP7_75t_L g659 ( .A(n_542), .Y(n_659) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_554), .Y(n_542) );
INVx5_ASAP7_75t_SL g579 ( .A(n_544), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_544), .B(n_649), .Y(n_648) );
AOI311xp33_ASAP7_75t_L g667 ( .A1(n_544), .A2(n_668), .A3(n_670), .B(n_671), .C(n_677), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_544), .A2(n_615), .B(n_703), .C(n_706), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
INVxp67_ASAP7_75t_L g622 ( .A(n_554), .Y(n_622) );
NAND4xp25_ASAP7_75t_SL g555 ( .A(n_556), .B(n_559), .C(n_565), .D(n_567), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_556), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g613 ( .A(n_557), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_560), .B(n_566), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_560), .B(n_573), .Y(n_693) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_561), .B(n_574), .Y(n_711) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
INVxp67_ASAP7_75t_L g621 ( .A(n_563), .Y(n_621) );
AND2x4_ASAP7_75t_L g573 ( .A(n_564), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g647 ( .A(n_564), .B(n_586), .Y(n_647) );
INVx1_ASAP7_75t_L g674 ( .A(n_564), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_564), .B(n_661), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_565), .B(n_635), .Y(n_655) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_566), .B(n_588), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_566), .B(n_635), .Y(n_734) );
INVx1_ASAP7_75t_L g745 ( .A(n_567), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B(n_575), .C(n_583), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_571), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g625 ( .A(n_571), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
AND2x2_ASAP7_75t_L g584 ( .A(n_573), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_573), .B(n_635), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_573), .B(n_654), .Y(n_678) );
OR2x2_ASAP7_75t_L g594 ( .A(n_574), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g626 ( .A(n_574), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_574), .B(n_586), .Y(n_641) );
AND2x2_ASAP7_75t_L g698 ( .A(n_574), .B(n_654), .Y(n_698) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_574), .Y(n_705) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_576), .A2(n_588), .B1(n_710), .B2(n_712), .C(n_715), .Y(n_709) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g599 ( .A(n_579), .B(n_582), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_579), .B(n_649), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_579), .B(n_606), .Y(n_714) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g699 ( .A(n_581), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g713 ( .A(n_581), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_582), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_582), .B(n_603), .Y(n_610) );
AND2x2_ASAP7_75t_L g680 ( .A(n_582), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_582), .B(n_629), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_582), .B(n_730), .Y(n_729) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_587), .B(n_589), .Y(n_583) );
INVx2_ASAP7_75t_L g616 ( .A(n_584), .Y(n_616) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g636 ( .A(n_586), .Y(n_636) );
OR2x2_ASAP7_75t_L g640 ( .A(n_588), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g743 ( .A(n_588), .B(n_711), .Y(n_743) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g747 ( .A(n_594), .Y(n_747) );
INVx2_ASAP7_75t_SL g661 ( .A(n_595), .Y(n_661) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_598), .A2(n_679), .B(n_743), .C(n_744), .Y(n_742) );
OAI322xp33_ASAP7_75t_SL g611 ( .A1(n_599), .A2(n_612), .A3(n_615), .B1(n_616), .B2(n_617), .C1(n_619), .C2(n_622), .Y(n_611) );
INVx2_ASAP7_75t_L g631 ( .A(n_599), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_607), .B1(n_608), .B2(n_610), .C(n_611), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp33_ASAP7_75t_SL g677 ( .A1(n_602), .A2(n_678), .B1(n_679), .B2(n_682), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_603), .B(n_606), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_603), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g676 ( .A(n_605), .B(n_638), .Y(n_676) );
INVx1_ASAP7_75t_L g666 ( .A(n_606), .Y(n_666) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_610), .A2(n_720), .B(n_722), .Y(n_719) );
AOI21xp33_ASAP7_75t_L g644 ( .A1(n_612), .A2(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp67_ASAP7_75t_SL g673 ( .A(n_614), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_614), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g730 ( .A(n_615), .Y(n_730) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_651), .C(n_667), .D(n_683), .Y(n_623) );
AOI211xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_632), .C(n_644), .Y(n_624) );
INVx1_ASAP7_75t_L g716 ( .A(n_625), .Y(n_716) );
AND2x2_ASAP7_75t_L g664 ( .A(n_626), .B(n_647), .Y(n_664) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_631), .B(n_666), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B1(n_640), .B2(n_642), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_634), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_635), .A2(n_674), .B(n_697), .C(n_699), .Y(n_696) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g681 ( .A(n_638), .Y(n_681) );
INVx1_ASAP7_75t_L g741 ( .A(n_639), .Y(n_741) );
NAND2xp33_ASAP7_75t_SL g731 ( .A(n_640), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g670 ( .A(n_649), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B(n_656), .C(n_658), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_663), .B2(n_665), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_661), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_666), .B(n_687), .Y(n_749) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_675), .B(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_689), .B1(n_692), .B2(n_694), .C(n_696), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_699), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g701 ( .A(n_702), .B(n_709), .C(n_719), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_728), .C(n_737), .Y(n_725) );
INVx1_ASAP7_75t_L g746 ( .A(n_726), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_733), .B2(n_735), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22x1_ASAP7_75t_SL g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_759), .Y(n_758) );
endmodule