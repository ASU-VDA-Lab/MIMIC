module fake_jpeg_14562_n_219 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_45),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_SL g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_0),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_3),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_19),
.B1(n_21),
.B2(n_24),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_19),
.B1(n_34),
.B2(n_32),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_41),
.B1(n_18),
.B2(n_32),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_35),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_22),
.B1(n_31),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_25),
.B1(n_22),
.B2(n_29),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_72),
.Y(n_120)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_37),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_86),
.B1(n_90),
.B2(n_93),
.Y(n_108)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_89),
.Y(n_112)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_71),
.B1(n_53),
.B2(n_54),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_46),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_42),
.B1(n_27),
.B2(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_44),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_94),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

OAI32xp33_ASAP7_75t_L g90 ( 
.A1(n_56),
.A2(n_27),
.A3(n_18),
.B1(n_44),
.B2(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_44),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_63),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_44),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_97),
.C(n_69),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_42),
.B1(n_18),
.B2(n_26),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_3),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_26),
.C(n_42),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_69),
.C(n_67),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_16),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_15),
.Y(n_105)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_61),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_109),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_70),
.B1(n_61),
.B2(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_121),
.B1(n_6),
.B2(n_7),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_105),
.B(n_117),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_113),
.B(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_15),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_77),
.B(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_118),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_54),
.B1(n_53),
.B2(n_63),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_81),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_14),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_87),
.B(n_5),
.Y(n_118)
);

OAI22x1_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_75),
.Y(n_128)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_89),
.Y(n_124)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_92),
.B(n_78),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_139),
.B(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_115),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_88),
.C(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_144),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_81),
.B1(n_85),
.B2(n_82),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_108),
.B1(n_119),
.B2(n_120),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_73),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_72),
.C(n_12),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_106),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_103),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_138),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_159),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_157),
.B(n_9),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_135),
.A2(n_104),
.B(n_100),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_118),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_158),
.B(n_10),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_127),
.Y(n_159)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_9),
.B(n_10),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_147),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_135),
.B1(n_133),
.B2(n_144),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_166),
.A2(n_178),
.B1(n_164),
.B2(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_134),
.C(n_125),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_189)
);

AND2x4_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_136),
.Y(n_170)
);

BUFx12f_ASAP7_75t_SL g190 ( 
.A(n_170),
.Y(n_190)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_142),
.A3(n_127),
.B1(n_126),
.B2(n_140),
.C1(n_133),
.C2(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_108),
.C(n_12),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_148),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_177),
.B(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_186),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_188),
.Y(n_194)
);

AOI31xp67_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_170),
.A3(n_178),
.B(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_145),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_190),
.A2(n_177),
.B(n_176),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_169),
.C(n_173),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_198),
.C(n_187),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_160),
.C(n_179),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_200),
.A2(n_204),
.B(n_196),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_180),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_201),
.A2(n_205),
.B(n_150),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_158),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g203 ( 
.A(n_193),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_206),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_185),
.B(n_176),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_155),
.B1(n_170),
.B2(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_210),
.Y(n_215)
);

AOI31xp67_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_191),
.A3(n_150),
.B(n_155),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_163),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_202),
.C(n_194),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_13),
.C(n_215),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_216),
.A2(n_212),
.B(n_13),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_217),
.Y(n_219)
);


endmodule