module real_aes_6413_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_453;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g263 ( .A(n_0), .Y(n_263) );
AOI21xp33_ASAP7_75t_L g205 ( .A1(n_1), .A2(n_206), .B(n_212), .Y(n_205) );
INVx1_ASAP7_75t_L g186 ( .A(n_2), .Y(n_186) );
AND2x6_ASAP7_75t_L g211 ( .A(n_2), .B(n_184), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_2), .B(n_516), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_3), .A2(n_166), .B1(n_172), .B2(n_173), .Y(n_165) );
INVx1_ASAP7_75t_L g172 ( .A(n_3), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_3), .A2(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g222 ( .A(n_4), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_5), .B(n_296), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_6), .Y(n_123) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_7), .A2(n_23), .B1(n_91), .B2(n_92), .Y(n_90) );
INVx1_ASAP7_75t_L g204 ( .A(n_8), .Y(n_204) );
INVx1_ASAP7_75t_L g310 ( .A(n_9), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_10), .B(n_251), .Y(n_325) );
AO22x2_ASAP7_75t_L g94 ( .A1(n_11), .A2(n_24), .B1(n_91), .B2(n_95), .Y(n_94) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_12), .B(n_206), .Y(n_275) );
AOI22xp5_ASAP7_75t_SL g511 ( .A1(n_12), .A2(n_80), .B1(n_81), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_12), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_13), .A2(n_167), .B1(n_168), .B2(n_169), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_13), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_14), .B(n_197), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g307 ( .A1(n_15), .A2(n_308), .B(n_309), .C(n_311), .Y(n_307) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_16), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_17), .B(n_220), .Y(n_265) );
XOR2xp5_ASAP7_75t_L g522 ( .A(n_18), .B(n_82), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g133 ( .A1(n_19), .A2(n_31), .B1(n_134), .B2(n_138), .Y(n_133) );
AOI22xp33_ASAP7_75t_SL g140 ( .A1(n_20), .A2(n_29), .B1(n_141), .B2(n_145), .Y(n_140) );
INVx1_ASAP7_75t_L g241 ( .A(n_21), .Y(n_241) );
INVx2_ASAP7_75t_L g209 ( .A(n_22), .Y(n_209) );
OAI221xp5_ASAP7_75t_L g177 ( .A1(n_24), .A2(n_40), .B1(n_50), .B2(n_178), .C(n_179), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_24), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_25), .A2(n_211), .B(n_215), .C(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g521 ( .A(n_25), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_26), .A2(n_33), .B1(n_107), .B2(n_113), .Y(n_106) );
INVx1_ASAP7_75t_L g239 ( .A(n_27), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_28), .B(n_220), .Y(n_324) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_30), .A2(n_35), .B1(n_170), .B2(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_30), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_32), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_34), .B(n_206), .Y(n_298) );
INVx1_ASAP7_75t_L g171 ( .A(n_35), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_36), .B(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_37), .A2(n_215), .B1(n_235), .B2(n_237), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_38), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_39), .Y(n_260) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_40), .A2(n_59), .B1(n_91), .B2(n_95), .Y(n_100) );
INVxp67_ASAP7_75t_L g181 ( .A(n_40), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_41), .A2(n_219), .B(n_221), .C(n_224), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_42), .Y(n_328) );
INVx1_ASAP7_75t_L g213 ( .A(n_43), .Y(n_213) );
INVx1_ASAP7_75t_L g184 ( .A(n_44), .Y(n_184) );
AOI22xp33_ASAP7_75t_SL g151 ( .A1(n_45), .A2(n_65), .B1(n_152), .B2(n_154), .Y(n_151) );
INVx1_ASAP7_75t_L g203 ( .A(n_46), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_47), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_48), .Y(n_101) );
AOI22xp33_ASAP7_75t_SL g157 ( .A1(n_49), .A2(n_52), .B1(n_158), .B2(n_162), .Y(n_157) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_50), .A2(n_66), .B1(n_91), .B2(n_92), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_51), .Y(n_85) );
A2O1A1Ixp33_ASAP7_75t_SL g250 ( .A1(n_53), .A2(n_224), .B(n_251), .C(n_252), .Y(n_250) );
INVxp67_ASAP7_75t_L g253 ( .A(n_54), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_55), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_56), .Y(n_126) );
INVx1_ASAP7_75t_L g321 ( .A(n_57), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_58), .A2(n_211), .B(n_215), .C(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_60), .B(n_264), .Y(n_278) );
INVx2_ASAP7_75t_L g201 ( .A(n_61), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_62), .A2(n_80), .B1(n_81), .B2(n_164), .Y(n_79) );
INVx1_ASAP7_75t_L g164 ( .A(n_62), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_63), .B(n_251), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_64), .A2(n_211), .B(n_215), .C(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_67), .B(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_68), .Y(n_268) );
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_69), .A2(n_211), .B(n_215), .C(n_293), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_70), .Y(n_300) );
INVx1_ASAP7_75t_L g249 ( .A(n_71), .Y(n_249) );
CKINVDCx16_ASAP7_75t_R g306 ( .A(n_72), .Y(n_306) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_73), .B(n_264), .Y(n_294) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
INVx1_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_75), .B(n_199), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_76), .A2(n_206), .B(n_248), .Y(n_247) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_174), .B1(n_187), .B2(n_506), .C(n_510), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_165), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
AND3x1_ASAP7_75t_L g82 ( .A(n_83), .B(n_132), .C(n_150), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_105), .C(n_122), .Y(n_83) );
OAI22xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_86), .B1(n_101), .B2(n_102), .Y(n_84) );
BUFx3_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_96), .Y(n_87) );
INVx2_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
OR2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
AND2x2_ASAP7_75t_L g104 ( .A(n_89), .B(n_94), .Y(n_104) );
AND2x2_ASAP7_75t_L g137 ( .A(n_89), .B(n_111), .Y(n_137) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g112 ( .A(n_90), .B(n_100), .Y(n_112) );
AND2x2_ASAP7_75t_L g119 ( .A(n_90), .B(n_94), .Y(n_119) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g95 ( .A(n_93), .Y(n_95) );
INVx2_ASAP7_75t_L g111 ( .A(n_94), .Y(n_111) );
INVx1_ASAP7_75t_L g148 ( .A(n_94), .Y(n_148) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
NAND2x1p5_ASAP7_75t_L g103 ( .A(n_97), .B(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g139 ( .A(n_97), .B(n_137), .Y(n_139) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_99), .Y(n_97) );
INVx1_ASAP7_75t_L g110 ( .A(n_98), .Y(n_110) );
INVx1_ASAP7_75t_L g121 ( .A(n_98), .Y(n_121) );
INVx1_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_98), .B(n_100), .Y(n_149) );
AND2x2_ASAP7_75t_L g120 ( .A(n_99), .B(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g144 ( .A(n_100), .B(n_131), .Y(n_144) );
BUFx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g143 ( .A(n_104), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g163 ( .A(n_104), .B(n_120), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_116), .Y(n_105) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
INVx1_ASAP7_75t_L g115 ( .A(n_110), .Y(n_115) );
INVx1_ASAP7_75t_L g125 ( .A(n_111), .Y(n_125) );
AND2x4_ASAP7_75t_L g114 ( .A(n_112), .B(n_115), .Y(n_114) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_112), .B(n_125), .Y(n_124) );
BUFx12f_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx1_ASAP7_75t_L g128 ( .A(n_119), .Y(n_128) );
AND2x2_ASAP7_75t_L g136 ( .A(n_120), .B(n_137), .Y(n_136) );
AND2x6_ASAP7_75t_L g160 ( .A(n_120), .B(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_126), .B2(n_127), .Y(n_122) );
OR2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_140), .Y(n_132) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g153 ( .A(n_137), .B(n_144), .Y(n_153) );
AND2x4_ASAP7_75t_L g155 ( .A(n_137), .B(n_156), .Y(n_155) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx8_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx6_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
OR2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_157), .Y(n_150) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx11_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_166), .Y(n_173) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_176), .Y(n_175) );
AND3x1_ASAP7_75t_SL g176 ( .A(n_177), .B(n_182), .C(n_185), .Y(n_176) );
INVxp67_ASAP7_75t_L g516 ( .A(n_177), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_182), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_182), .A2(n_215), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g526 ( .A(n_182), .Y(n_526) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_183), .B(n_186), .Y(n_520) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
OR2x2_ASAP7_75t_SL g525 ( .A(n_185), .B(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
HB1xp67_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND3x1_ASAP7_75t_L g191 ( .A(n_192), .B(n_428), .C(n_473), .Y(n_191) );
NOR4xp25_ASAP7_75t_L g192 ( .A(n_193), .B(n_351), .C(n_392), .D(n_409), .Y(n_192) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_255), .B(n_271), .C(n_313), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_229), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_195), .B(n_256), .Y(n_255) );
NOR4xp25_ASAP7_75t_L g375 ( .A(n_195), .B(n_369), .C(n_376), .D(n_382), .Y(n_375) );
AND2x2_ASAP7_75t_L g448 ( .A(n_195), .B(n_337), .Y(n_448) );
AND2x2_ASAP7_75t_L g467 ( .A(n_195), .B(n_413), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_195), .B(n_462), .Y(n_476) );
AND2x2_ASAP7_75t_L g489 ( .A(n_195), .B(n_270), .Y(n_489) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_SL g334 ( .A(n_196), .Y(n_334) );
AND2x2_ASAP7_75t_L g341 ( .A(n_196), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g391 ( .A(n_196), .B(n_230), .Y(n_391) );
AND2x2_ASAP7_75t_SL g402 ( .A(n_196), .B(n_337), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_196), .B(n_230), .Y(n_406) );
AND2x2_ASAP7_75t_L g415 ( .A(n_196), .B(n_340), .Y(n_415) );
BUFx2_ASAP7_75t_L g438 ( .A(n_196), .Y(n_438) );
AND2x2_ASAP7_75t_L g442 ( .A(n_196), .B(n_246), .Y(n_442) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_205), .B(n_227), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_198), .B(n_285), .Y(n_284) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_199), .A2(n_247), .B(n_254), .Y(n_246) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx1_ASAP7_75t_L g232 ( .A(n_200), .Y(n_232) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
AND2x2_ASAP7_75t_SL g228 ( .A(n_201), .B(n_202), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
BUFx2_ASAP7_75t_L g304 ( .A(n_206), .Y(n_304) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_211), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g243 ( .A(n_207), .B(n_211), .Y(n_243) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g216 ( .A(n_209), .Y(n_216) );
INVx1_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
INVx1_ASAP7_75t_L g217 ( .A(n_210), .Y(n_217) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_210), .Y(n_220) );
INVx3_ASAP7_75t_L g223 ( .A(n_210), .Y(n_223) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_210), .Y(n_238) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
INVx4_ASAP7_75t_SL g226 ( .A(n_211), .Y(n_226) );
BUFx3_ASAP7_75t_L g509 ( .A(n_211), .Y(n_509) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_218), .C(n_226), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_214), .A2(n_226), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_214), .A2(n_226), .B(n_306), .C(n_307), .Y(n_305) );
INVx5_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g508 ( .A(n_215), .B(n_509), .Y(n_508) );
AND2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_217), .Y(n_215) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_216), .Y(n_225) );
BUFx3_ASAP7_75t_L g282 ( .A(n_216), .Y(n_282) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx4_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_223), .B(n_253), .Y(n_252) );
INVx5_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_225), .Y(n_297) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_226), .A2(n_234), .B1(n_242), .B2(n_243), .Y(n_233) );
INVx1_ASAP7_75t_L g269 ( .A(n_228), .Y(n_269) );
INVx2_ASAP7_75t_L g290 ( .A(n_228), .Y(n_290) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_228), .A2(n_303), .B(n_312), .Y(n_302) );
OR2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_246), .Y(n_229) );
AND2x2_ASAP7_75t_L g270 ( .A(n_230), .B(n_246), .Y(n_270) );
BUFx2_ASAP7_75t_L g344 ( .A(n_230), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_230), .A2(n_377), .B1(n_379), .B2(n_380), .Y(n_376) );
OR2x2_ASAP7_75t_L g398 ( .A(n_230), .B(n_258), .Y(n_398) );
AND2x2_ASAP7_75t_L g462 ( .A(n_230), .B(n_340), .Y(n_462) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g330 ( .A(n_231), .B(n_258), .Y(n_330) );
AND2x2_ASAP7_75t_L g337 ( .A(n_231), .B(n_246), .Y(n_337) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_231), .Y(n_379) );
OR2x2_ASAP7_75t_L g414 ( .A(n_231), .B(n_257), .Y(n_414) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_244), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_232), .B(n_245), .Y(n_244) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_232), .A2(n_259), .B(n_267), .Y(n_258) );
INVx2_ASAP7_75t_L g283 ( .A(n_232), .Y(n_283) );
INVx2_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_SL g237 ( .A1(n_238), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_237) );
INVx2_ASAP7_75t_L g240 ( .A(n_238), .Y(n_240) );
INVx4_ASAP7_75t_L g308 ( .A(n_238), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_243), .A2(n_260), .B(n_261), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_243), .A2(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g333 ( .A(n_246), .Y(n_333) );
INVx3_ASAP7_75t_L g342 ( .A(n_246), .Y(n_342) );
BUFx2_ASAP7_75t_L g366 ( .A(n_246), .Y(n_366) );
AND2x2_ASAP7_75t_L g399 ( .A(n_246), .B(n_334), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_255), .A2(n_485), .B1(n_486), .B2(n_487), .Y(n_484) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_270), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_257), .B(n_342), .Y(n_346) );
INVx1_ASAP7_75t_L g374 ( .A(n_257), .Y(n_374) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g340 ( .A(n_258), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B(n_265), .C(n_266), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_269), .B(n_300), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_269), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g352 ( .A(n_270), .Y(n_352) );
NAND2x1_ASAP7_75t_SL g271 ( .A(n_272), .B(n_286), .Y(n_271) );
AND2x2_ASAP7_75t_L g350 ( .A(n_272), .B(n_301), .Y(n_350) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_272), .Y(n_424) );
AND2x2_ASAP7_75t_L g451 ( .A(n_272), .B(n_371), .Y(n_451) );
AND2x2_ASAP7_75t_L g459 ( .A(n_272), .B(n_421), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_272), .B(n_316), .Y(n_486) );
INVx3_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g335 ( .A(n_273), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g356 ( .A(n_273), .Y(n_356) );
INVx1_ASAP7_75t_L g362 ( .A(n_273), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_273), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g395 ( .A(n_273), .B(n_319), .Y(n_395) );
OR2x2_ASAP7_75t_L g433 ( .A(n_273), .B(n_388), .Y(n_433) );
AOI32xp33_ASAP7_75t_L g445 ( .A1(n_273), .A2(n_446), .A3(n_449), .B1(n_450), .B2(n_451), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_273), .B(n_421), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_273), .B(n_381), .Y(n_496) );
OR2x6_ASAP7_75t_L g273 ( .A(n_274), .B(n_284), .Y(n_273) );
AOI21xp5_ASAP7_75t_SL g274 ( .A1(n_275), .A2(n_276), .B(n_283), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_279), .B(n_280), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_280), .A2(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
INVx1_ASAP7_75t_L g326 ( .A(n_283), .Y(n_326) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g407 ( .A(n_287), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_301), .Y(n_287) );
INVx1_ASAP7_75t_L g369 ( .A(n_288), .Y(n_369) );
AND2x2_ASAP7_75t_L g371 ( .A(n_288), .B(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_288), .B(n_318), .Y(n_388) );
AND2x2_ASAP7_75t_L g421 ( .A(n_288), .B(n_397), .Y(n_421) );
AND2x2_ASAP7_75t_L g458 ( .A(n_288), .B(n_319), .Y(n_458) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g316 ( .A(n_289), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_289), .B(n_318), .Y(n_348) );
AND2x2_ASAP7_75t_L g355 ( .A(n_289), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g396 ( .A(n_289), .B(n_397), .Y(n_396) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_299), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_292), .B(n_298), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_295), .B(n_297), .Y(n_293) );
INVx2_ASAP7_75t_L g372 ( .A(n_301), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_301), .B(n_318), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_301), .B(n_363), .Y(n_444) );
INVx1_ASAP7_75t_L g466 ( .A(n_301), .Y(n_466) );
INVx1_ASAP7_75t_L g483 ( .A(n_301), .Y(n_483) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g336 ( .A(n_302), .B(n_318), .Y(n_336) );
AND2x2_ASAP7_75t_L g358 ( .A(n_302), .B(n_319), .Y(n_358) );
INVx1_ASAP7_75t_L g397 ( .A(n_302), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_308), .B(n_310), .Y(n_309) );
AOI221x1_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_329), .B1(n_335), .B2(n_337), .C(n_338), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_314), .A2(n_402), .B1(n_469), .B2(n_470), .Y(n_468) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
AND2x2_ASAP7_75t_L g360 ( .A(n_315), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g455 ( .A(n_315), .B(n_335), .Y(n_455) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g411 ( .A(n_316), .B(n_336), .Y(n_411) );
INVx1_ASAP7_75t_L g423 ( .A(n_317), .Y(n_423) );
AND2x2_ASAP7_75t_L g434 ( .A(n_317), .B(n_421), .Y(n_434) );
AND2x2_ASAP7_75t_L g501 ( .A(n_317), .B(n_396), .Y(n_501) );
INVx2_ASAP7_75t_L g363 ( .A(n_318), .Y(n_363) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_326), .B(n_327), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_330), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g453 ( .A(n_330), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_331), .B(n_414), .Y(n_417) );
INVx3_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_332), .A2(n_453), .B(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NOR2xp33_ASAP7_75t_SL g475 ( .A(n_335), .B(n_361), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_336), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g427 ( .A(n_336), .B(n_355), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_336), .B(n_362), .Y(n_504) );
AND2x2_ASAP7_75t_L g373 ( .A(n_337), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g440 ( .A(n_337), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_343), .B(n_347), .Y(n_338) );
NAND2x1_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_340), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g389 ( .A(n_340), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_SL g401 ( .A(n_340), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_340), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g425 ( .A(n_341), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_341), .B(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_341), .B(n_344), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AOI211xp5_ASAP7_75t_L g412 ( .A1(n_344), .A2(n_383), .B(n_413), .C(n_415), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_344), .A2(n_431), .B1(n_434), .B2(n_435), .C(n_439), .Y(n_430) );
AND2x2_ASAP7_75t_L g426 ( .A(n_345), .B(n_379), .Y(n_426) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g386 ( .A(n_350), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g457 ( .A(n_350), .B(n_458), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_359), .C(n_384), .Y(n_351) );
NAND3xp33_ASAP7_75t_SL g470 ( .A(n_352), .B(n_471), .C(n_472), .Y(n_470) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_357), .Y(n_353) );
OR2x2_ASAP7_75t_L g443 ( .A(n_354), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_364), .B1(n_367), .B2(n_373), .C(n_375), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_361), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_361), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g383 ( .A(n_366), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_366), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_422) );
OR2x2_ASAP7_75t_L g503 ( .A(n_366), .B(n_414), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVxp67_ASAP7_75t_L g477 ( .A(n_369), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_371), .B(n_492), .Y(n_491) );
INVxp67_ASAP7_75t_L g378 ( .A(n_372), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_374), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_374), .B(n_421), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_374), .B(n_441), .Y(n_480) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_378), .Y(n_404) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g494 ( .A(n_383), .B(n_414), .Y(n_494) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g472 ( .A(n_389), .Y(n_472) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI322xp33_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_403), .C1(n_405), .C2(n_407), .Y(n_392) );
OAI322xp33_ASAP7_75t_L g474 ( .A1(n_393), .A2(n_475), .A3(n_476), .B1(n_477), .B2(n_478), .C1(n_479), .C2(n_481), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx4_ASAP7_75t_L g408 ( .A(n_395), .Y(n_408) );
AND2x2_ASAP7_75t_L g469 ( .A(n_395), .B(n_421), .Y(n_469) );
AND2x2_ASAP7_75t_L g482 ( .A(n_395), .B(n_483), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_398), .Y(n_493) );
INVx1_ASAP7_75t_L g471 ( .A(n_399), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
OR2x2_ASAP7_75t_L g405 ( .A(n_401), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g488 ( .A(n_401), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_401), .B(n_442), .Y(n_499) );
OR2x2_ASAP7_75t_L g432 ( .A(n_404), .B(n_433), .Y(n_432) );
INVxp33_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
OAI221xp5_ASAP7_75t_SL g409 ( .A1(n_408), .A2(n_410), .B1(n_412), .B2(n_416), .C(n_418), .Y(n_409) );
NOR2xp67_ASAP7_75t_L g465 ( .A(n_408), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g492 ( .A(n_408), .Y(n_492) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx3_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
AOI322xp5_ASAP7_75t_L g456 ( .A1(n_415), .A2(n_440), .A3(n_457), .B1(n_459), .B2(n_460), .C1(n_463), .C2(n_467), .Y(n_456) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B1(n_426), .B2(n_427), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_452), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_430), .B(n_445), .Y(n_429) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_433), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
NAND2xp33_ASAP7_75t_SL g450 ( .A(n_436), .B(n_447), .Y(n_450) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
OAI322xp33_ASAP7_75t_L g490 ( .A1(n_438), .A2(n_491), .A3(n_493), .B1(n_494), .B2(n_495), .C1(n_497), .C2(n_500), .Y(n_490) );
AOI21xp33_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_441), .B(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_448), .B(n_496), .Y(n_505) );
OAI211xp5_ASAP7_75t_SL g452 ( .A1(n_453), .A2(n_454), .B(n_456), .C(n_468), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NOR4xp25_ASAP7_75t_L g473 ( .A(n_474), .B(n_484), .C(n_490), .D(n_502), .Y(n_473) );
INVxp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
CKINVDCx14_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
OAI21xp5_ASAP7_75t_SL g502 ( .A1(n_503), .A2(n_504), .B(n_505), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_508), .Y(n_507) );
OAI322xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_513), .A3(n_517), .B1(n_518), .B2(n_521), .C1(n_522), .C2(n_523), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
CKINVDCx16_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
endmodule