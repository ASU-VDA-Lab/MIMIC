module fake_jpeg_21255_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_4),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_49),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_46),
.A2(n_43),
.B1(n_38),
.B2(n_7),
.Y(n_60)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_36),
.B(n_1),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_51),
.Y(n_56)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_5),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_3),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_63),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_44),
.B1(n_40),
.B2(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_41),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_60),
.A2(n_38),
.B1(n_41),
.B2(n_35),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_65),
.A2(n_70),
.B1(n_73),
.B2(n_67),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_58),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_39),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_5),
.C(n_6),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_32),
.B1(n_15),
.B2(n_18),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_56),
.Y(n_76)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_81),
.C(n_7),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_65),
.A2(n_62),
.B1(n_55),
.B2(n_19),
.Y(n_80)
);

NOR2xp67_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_82),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_6),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_71),
.B(n_68),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_82),
.B(n_11),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_8),
.C(n_9),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_86),
.A2(n_68),
.B1(n_75),
.B2(n_8),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_91),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_90),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_85),
.Y(n_94)
);

AOI321xp33_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_92),
.A3(n_83),
.B1(n_14),
.B2(n_20),
.C(n_21),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_10),
.B(n_13),
.C(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_31),
.Y(n_98)
);


endmodule