module fake_jpeg_19052_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_1),
.B(n_11),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_70),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_60),
.Y(n_78)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_79),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_51),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_54),
.B(n_41),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_71),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_94),
.Y(n_109)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_75),
.A2(n_55),
.B1(n_42),
.B2(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_100),
.B1(n_43),
.B2(n_21),
.Y(n_104)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_0),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_2),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_57),
.B1(n_64),
.B2(n_63),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_50),
.B1(n_61),
.B2(n_59),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_103),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_49),
.B(n_41),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_102),
.A2(n_113),
.B(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_62),
.B1(n_48),
.B2(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_111),
.Y(n_124)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_0),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_1),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_25),
.B(n_4),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_115),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_113),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_108),
.C(n_114),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_2),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_120),
.B(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_127),
.B(n_125),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_129),
.B(n_121),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_124),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_123),
.C(n_109),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_119),
.B(n_122),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_36),
.B(n_16),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_10),
.C(n_18),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

BUFx24_ASAP7_75t_SL g139 ( 
.A(n_138),
.Y(n_139)
);

NAND2xp33_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_19),
.Y(n_140)
);


endmodule