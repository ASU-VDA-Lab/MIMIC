module fake_jpeg_28334_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_43),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_18),
.B(n_0),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_18),
.B1(n_25),
.B2(n_28),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_55),
.B1(n_64),
.B2(n_30),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_25),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_39),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_34),
.A2(n_23),
.B1(n_27),
.B2(n_16),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_59),
.Y(n_78)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_34),
.A2(n_31),
.B1(n_21),
.B2(n_29),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_24),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_30),
.Y(n_72)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_62),
.B1(n_38),
.B2(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_35),
.B1(n_53),
.B2(n_21),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_83),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_38),
.B1(n_40),
.B2(n_36),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_82),
.B1(n_88),
.B2(n_31),
.Y(n_111)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_86),
.B1(n_81),
.B2(n_76),
.Y(n_102)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_51),
.Y(n_101)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_40),
.B1(n_36),
.B2(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_47),
.B1(n_59),
.B2(n_40),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_90),
.A2(n_96),
.B1(n_104),
.B2(n_105),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_36),
.B1(n_47),
.B2(n_63),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_111),
.B1(n_68),
.B2(n_16),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_49),
.B1(n_51),
.B2(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_97),
.B(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_84),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_39),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_101),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_85),
.A2(n_53),
.B1(n_66),
.B2(n_50),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_72),
.A2(n_35),
.B1(n_50),
.B2(n_16),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_109),
.B1(n_68),
.B2(n_19),
.Y(n_129)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_87),
.B1(n_80),
.B2(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_16),
.B1(n_27),
.B2(n_29),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_118),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_75),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_122),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_46),
.C(n_70),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_119),
.C(n_126),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_106),
.C(n_101),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_46),
.C(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_129),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_24),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_71),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_128),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_46),
.C(n_87),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_71),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_22),
.B1(n_19),
.B2(n_26),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_22),
.B1(n_19),
.B2(n_26),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_116),
.A2(n_100),
.B(n_99),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_138),
.B(n_151),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_100),
.B(n_99),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_107),
.B1(n_104),
.B2(n_108),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_148),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_108),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_152),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_132),
.B1(n_121),
.B2(n_133),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_109),
.B1(n_103),
.B2(n_93),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_103),
.B1(n_71),
.B2(n_26),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_103),
.C(n_26),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_137),
.C(n_119),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_168),
.C(n_174),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_139),
.A2(n_118),
.B(n_116),
.Y(n_159)
);

NAND2xp67_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_161),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_130),
.B(n_129),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_141),
.A2(n_131),
.B(n_122),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_173),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_8),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_0),
.B(n_2),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_9),
.C(n_3),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_177),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_0),
.B(n_4),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_4),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_187),
.Y(n_209)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_188),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_152),
.B1(n_153),
.B2(n_146),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_195),
.B1(n_192),
.B2(n_165),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_137),
.C(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_176),
.C(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_149),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_163),
.B(n_181),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_136),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_166),
.A2(n_140),
.B1(n_144),
.B2(n_147),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_164),
.B1(n_172),
.B2(n_165),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_140),
.B1(n_143),
.B2(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_196),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_194),
.Y(n_197)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_197),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_182),
.B(n_186),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_185),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_205),
.C(n_210),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_201),
.A2(n_202),
.B1(n_184),
.B2(n_195),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_203),
.B(n_198),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_161),
.C(n_155),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_206),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_154),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_4),
.C(n_5),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_216),
.B1(n_204),
.B2(n_207),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_7),
.B(n_9),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_186),
.B1(n_182),
.B2(n_183),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_218),
.C(n_221),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_222),
.B(n_10),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_5),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_6),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_209),
.C(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_228),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_231),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_202),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_226),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_210),
.Y(n_227)
);

AOI31xp33_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_221),
.A3(n_11),
.B(n_12),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_6),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_199),
.C(n_9),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_15),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_10),
.B(n_11),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_219),
.B1(n_218),
.B2(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_234),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_13),
.B(n_14),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_12),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_223),
.C(n_228),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_240),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_236),
.B(n_232),
.C(n_15),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_241),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_248),
.B(n_244),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_14),
.Y(n_250)
);


endmodule