module fake_jpeg_10104_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_SL g7 ( 
.A(n_5),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_6),
.Y(n_11)
);

INVx3_ASAP7_75t_SL g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

OAI32xp33_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_8),
.B1(n_12),
.B2(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_11),
.B(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_4),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_7),
.B(n_12),
.C(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_27),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_9),
.B1(n_10),
.B2(n_8),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_13),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_13),
.C(n_15),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_27),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_29),
.C(n_33),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.C(n_34),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_21),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_41),
.Y(n_43)
);


endmodule