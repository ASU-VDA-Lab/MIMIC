module fake_jpeg_6205_n_75 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_75);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_75;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_74;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_35;
wire n_48;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_31),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_51),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_21),
.B1(n_1),
.B2(n_4),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_53),
.B1(n_42),
.B2(n_41),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_54),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_23),
.B1(n_10),
.B2(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_59),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_45),
.B(n_44),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_38),
.B(n_36),
.Y(n_62)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_0),
.B1(n_13),
.B2(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_64),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_63),
.A2(n_57),
.B1(n_56),
.B2(n_0),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_26),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_61),
.C(n_18),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_68),
.Y(n_69)
);

BUFx4f_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_15),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_27),
.B(n_28),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_32),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_33),
.Y(n_75)
);


endmodule