module fake_jpeg_16732_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_37),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_30),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_40),
.B1(n_20),
.B2(n_24),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_23),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_24),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_68),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_40),
.B1(n_37),
.B2(n_31),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_58),
.A2(n_41),
.B1(n_35),
.B2(n_34),
.Y(n_106)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_37),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_61),
.B(n_77),
.Y(n_99)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_81),
.B1(n_41),
.B2(n_51),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_66),
.A2(n_28),
.B1(n_50),
.B2(n_16),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_19),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_72),
.Y(n_97)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_32),
.CON(n_70),
.SN(n_70)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_16),
.B(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_79),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_29),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_36),
.B1(n_21),
.B2(n_29),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_78),
.B1(n_27),
.B2(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_26),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_38),
.B1(n_25),
.B2(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_22),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_82),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_25),
.B1(n_21),
.B2(n_18),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_16),
.Y(n_82)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_34),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_102),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_52),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_82),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_52),
.A3(n_38),
.B1(n_28),
.B2(n_34),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_66),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_106),
.B1(n_109),
.B2(n_3),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_100),
.Y(n_112)
);

OAI22x1_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_72),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_0),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_105),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_2),
.Y(n_105)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_34),
.B1(n_35),
.B2(n_5),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_61),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_118),
.B(n_90),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_SL g145 ( 
.A(n_113),
.B(n_128),
.C(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_119),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_129),
.C(n_103),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_83),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_92),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_89),
.B(n_76),
.Y(n_123)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_125),
.Y(n_140)
);

INVx13_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_65),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_133),
.Y(n_151)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_105),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_149),
.Y(n_156)
);

NOR3xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_97),
.C(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_142),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_106),
.B(n_95),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_154),
.B(n_155),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_116),
.C(n_132),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_112),
.A2(n_109),
.B1(n_90),
.B2(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_153),
.A2(n_130),
.B1(n_117),
.B2(n_119),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_113),
.A2(n_111),
.B(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_158),
.C(n_163),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_161),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_86),
.C(n_125),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_168),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_150),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_3),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_138),
.C(n_137),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_143),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_169),
.Y(n_195)
);

OA21x2_ASAP7_75t_SL g179 ( 
.A1(n_171),
.A2(n_146),
.B(n_145),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_173),
.B(n_156),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_163),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_162),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_182),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_135),
.C(n_153),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.C(n_166),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_145),
.C(n_148),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_165),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_189),
.C(n_193),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_190),
.A2(n_176),
.B(n_178),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_156),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_191),
.B(n_192),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_196),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_160),
.C(n_151),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_164),
.B(n_142),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_174),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_191),
.A2(n_183),
.B1(n_177),
.B2(n_175),
.Y(n_202)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_202),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_196),
.B(n_193),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_180),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_205),
.B(n_3),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_192),
.A2(n_147),
.B1(n_14),
.B2(n_12),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_187),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

OAI321xp33_ASAP7_75t_L g213 ( 
.A1(n_209),
.A2(n_201),
.A3(n_198),
.B1(n_199),
.B2(n_200),
.C(n_4),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_12),
.C(n_4),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_200),
.C(n_7),
.Y(n_214)
);

NOR3xp33_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_6),
.C(n_7),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_213),
.A2(n_215),
.B(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_219),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_212),
.C2(n_211),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_207),
.B(n_210),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_221),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_8),
.Y(n_223)
);


endmodule