module fake_jpeg_17206_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_62),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_42),
.C(n_53),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_77),
.B(n_81),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_51),
.B(n_50),
.C(n_40),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_79),
.B1(n_43),
.B2(n_1),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_48),
.B1(n_41),
.B2(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_84),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_0),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_41),
.B1(n_57),
.B2(n_44),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_92),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_90),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_66),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_79),
.B1(n_71),
.B2(n_58),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_93),
.A2(n_86),
.B1(n_85),
.B2(n_94),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_97),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_100),
.B(n_101),
.Y(n_114)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_108),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_4),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_111),
.A2(n_92),
.B(n_96),
.Y(n_120)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_103),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_120),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_111),
.B1(n_102),
.B2(n_99),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_87),
.B1(n_115),
.B2(n_99),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_126),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_23),
.C(n_33),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_124),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_122),
.B(n_22),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_21),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_131),
.A2(n_24),
.B1(n_32),
.B2(n_8),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_19),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_25),
.B(n_31),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_17),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_15),
.C(n_29),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_13),
.Y(n_137)
);


endmodule