module fake_jpeg_19173_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_36),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_36),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_54),
.B1(n_33),
.B2(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_53),
.B1(n_36),
.B2(n_33),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_24),
.B1(n_32),
.B2(n_19),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_23),
.B1(n_19),
.B2(n_27),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_R g59 ( 
.A(n_39),
.B(n_20),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_55),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_73),
.B(n_74),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_48),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_18),
.Y(n_105)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_34),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_44),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_89),
.B1(n_46),
.B2(n_57),
.Y(n_109)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_88),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_42),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_99),
.B1(n_100),
.B2(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_80),
.C(n_82),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_21),
.C(n_28),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_71),
.B1(n_77),
.B2(n_62),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_72),
.A2(n_34),
.B1(n_57),
.B2(n_46),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_57),
.B1(n_46),
.B2(n_49),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_21),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_63),
.B(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_105),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_57),
.B1(n_51),
.B2(n_47),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_46),
.B1(n_81),
.B2(n_68),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_28),
.B(n_21),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_87),
.B(n_2),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_121),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_67),
.B1(n_65),
.B2(n_70),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_47),
.B1(n_101),
.B2(n_66),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_64),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_46),
.B1(n_69),
.B2(n_93),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_28),
.B(n_21),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_126),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_92),
.B(n_14),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_135),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_132),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_133),
.C(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_86),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_131),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_105),
.C(n_96),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_90),
.B(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_91),
.B(n_79),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_141),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_113),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_97),
.B(n_2),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_85),
.Y(n_142)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_99),
.B1(n_94),
.B2(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_158),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_169),
.C(n_131),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_134),
.A2(n_107),
.B1(n_94),
.B2(n_116),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_112),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_154),
.A2(n_167),
.B(n_168),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_155),
.A2(n_128),
.B1(n_127),
.B2(n_135),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_101),
.B1(n_66),
.B2(n_85),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_101),
.B1(n_66),
.B2(n_114),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_97),
.B1(n_31),
.B2(n_16),
.Y(n_163)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_170),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_138),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_124),
.A2(n_21),
.B(n_97),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_140),
.A2(n_17),
.B(n_2),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_31),
.C(n_16),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_140),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_16),
.B1(n_17),
.B2(n_9),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_122),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_178),
.B(n_186),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_130),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_181),
.C(n_197),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_121),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_158),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_184),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_173),
.B1(n_163),
.B2(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_118),
.C(n_119),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_195),
.Y(n_217)
);

BUFx6f_ASAP7_75t_SL g184 ( 
.A(n_157),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_120),
.Y(n_186)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_149),
.A2(n_172),
.B1(n_152),
.B2(n_168),
.C(n_170),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_191),
.B(n_160),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_167),
.A2(n_132),
.B1(n_136),
.B2(n_123),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_136),
.B1(n_123),
.B2(n_139),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g195 ( 
.A1(n_146),
.A2(n_118),
.B(n_137),
.C(n_17),
.D(n_9),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_7),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_169),
.C(n_153),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_207),
.C(n_212),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_148),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_148),
.C(n_154),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_159),
.B1(n_164),
.B2(n_145),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_210),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_174),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_154),
.C(n_145),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_215),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_161),
.C(n_166),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_194),
.C(n_193),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_150),
.B1(n_3),
.B2(n_4),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_190),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_182),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_226),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_216),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_197),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_227),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_196),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_186),
.C(n_150),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_214),
.C(n_207),
.Y(n_235)
);

OA21x2_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_195),
.B(n_179),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_200),
.B(n_198),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_205),
.B(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_238),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_224),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_237),
.Y(n_255)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_198),
.B(n_200),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_240),
.A2(n_244),
.B(n_228),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_243),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_217),
.B(n_184),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_229),
.B1(n_189),
.B2(n_233),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_8),
.B1(n_13),
.B2(n_4),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_226),
.B1(n_230),
.B2(n_225),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_1),
.B(n_3),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_254),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_219),
.B(n_3),
.C(n_4),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_245),
.B(n_236),
.Y(n_257)
);

AOI21x1_ASAP7_75t_SL g268 ( 
.A1(n_257),
.A2(n_258),
.B(n_261),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_250),
.A2(n_245),
.B(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_255),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_267),
.A3(n_268),
.B1(n_5),
.B2(n_6),
.C1(n_220),
.C2(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_255),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_251),
.B1(n_253),
.B2(n_6),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_269),
.A2(n_251),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

AOI321xp33_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_256),
.A3(n_251),
.B1(n_6),
.B2(n_5),
.C(n_3),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_273),
.Y(n_275)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_271),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_269),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_274),
.Y(n_278)
);


endmodule