module fake_jpeg_21693_n_102 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_19),
.B(n_22),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_4),
.B1(n_6),
.B2(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_23),
.B1(n_18),
.B2(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_21),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_26),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_50),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_28),
.B1(n_24),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_57),
.B1(n_29),
.B2(n_22),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_27),
.B(n_15),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_56),
.B(n_26),
.Y(n_62)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_23),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_58),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_15),
.B(n_26),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_13),
.B1(n_29),
.B2(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_8),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_9),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_71),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_10),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_70),
.A2(n_48),
.B1(n_45),
.B2(n_64),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_49),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_55),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_80),
.B(n_73),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_43),
.CI(n_53),
.CON(n_75),
.SN(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_77),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_43),
.C(n_61),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_87),
.B(n_71),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_90),
.B(n_91),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_62),
.B(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_84),
.A2(n_77),
.B1(n_76),
.B2(n_75),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_85),
.C(n_84),
.Y(n_93)
);

OAI21x1_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_67),
.B(n_63),
.Y(n_98)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_75),
.C(n_69),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_95),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_66),
.C(n_68),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_46),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_99),
.B(n_46),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_100),
.A2(n_60),
.B1(n_97),
.B2(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_46),
.Y(n_102)
);


endmodule