module fake_jpeg_29095_n_132 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_26),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_32),
.Y(n_41)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_13),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_47),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_29),
.A2(n_25),
.B1(n_15),
.B2(n_12),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_46),
.B1(n_31),
.B2(n_17),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_12),
.B2(n_17),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_20),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_28),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_50),
.A2(n_25),
.B1(n_36),
.B2(n_15),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_25),
.B1(n_36),
.B2(n_30),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_55),
.B(n_28),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_36),
.B1(n_14),
.B2(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_60),
.Y(n_74)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_48),
.A2(n_47),
.B1(n_45),
.B2(n_27),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_67),
.Y(n_85)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_13),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_69),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_65),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_68),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_19),
.C(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_20),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g82 ( 
.A(n_71),
.B(n_73),
.C(n_10),
.Y(n_82)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_24),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_83),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_82),
.B(n_71),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_62),
.A2(n_23),
.B1(n_18),
.B2(n_16),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_61),
.C(n_67),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_63),
.B1(n_65),
.B2(n_64),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_93),
.A2(n_95),
.B(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_59),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_100),
.B(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_57),
.B1(n_56),
.B2(n_72),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_75),
.B(n_83),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_85),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_103),
.C(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_85),
.C(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_108),
.Y(n_115)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_111),
.C(n_114),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_92),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_101),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_103),
.A2(n_92),
.B(n_76),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_113),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_86),
.B(n_92),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

NAND4xp25_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_82),
.C(n_60),
.D(n_95),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_77),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_113),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_124),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_117),
.A2(n_110),
.B1(n_111),
.B2(n_3),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_37),
.B(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_120),
.B(n_124),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_128),
.C(n_18),
.Y(n_130)
);

OAI21x1_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_1),
.B(n_2),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_3),
.Y(n_132)
);


endmodule