module fake_ariane_2404_n_2048 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2048);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2048;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_1733;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx2_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_43),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_15),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_152),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_135),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_24),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_70),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_38),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_11),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_103),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_48),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_89),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_180),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_80),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_120),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_64),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_161),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_17),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_47),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_84),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_71),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_149),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_142),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_143),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_133),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_96),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_65),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_95),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_51),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_24),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_148),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_186),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_106),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_150),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_76),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_30),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_145),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_90),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_126),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_44),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_102),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_118),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_127),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_114),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_119),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_98),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_68),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_64),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_54),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_69),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_188),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_74),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_108),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_47),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_112),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_81),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_159),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_113),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_179),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_59),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_30),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_11),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_171),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_92),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_42),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_21),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_172),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_184),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_175),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_181),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_151),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_8),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_4),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_176),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_167),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_79),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_155),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_28),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_195),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_63),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_153),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_109),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_59),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_65),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_191),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_132),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_33),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_67),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_54),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_44),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_36),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_18),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_48),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_10),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_57),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_125),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_78),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_185),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_26),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_29),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_190),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_15),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_168),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_117),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_182),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_165),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_82),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_55),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_1),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_60),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_3),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_53),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_158),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_28),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_157),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_55),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_60),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_136),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_38),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_189),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_37),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_29),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_19),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_23),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_73),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_110),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_162),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_43),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_56),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_53),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_122),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_41),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_7),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_19),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_14),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_51),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_105),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_68),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_52),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_5),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_7),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_72),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_32),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_17),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_35),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_66),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_13),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_1),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_45),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_61),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_104),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_91),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_36),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_115),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_130),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_173),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_8),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_101),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_99),
.Y(n_374)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_178),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_9),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_88),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_124),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_58),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_94),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_86),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_10),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_87),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_177),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_58),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_39),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_0),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_198),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_174),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_57),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_42),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_49),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_201),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_31),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_156),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_197),
.Y(n_396)
);

BUFx8_ASAP7_75t_SL g397 ( 
.A(n_25),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_129),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_0),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_9),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_93),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_147),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_121),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_141),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_397),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_281),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_335),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_388),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_294),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_273),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_249),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_213),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_333),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_213),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_384),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_277),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_277),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_277),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_377),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_377),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_377),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_216),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_R g428 ( 
.A(n_251),
.B(n_202),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_325),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_206),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_274),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_256),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_204),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_205),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_274),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_262),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_211),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_329),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_329),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_206),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_360),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_207),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_263),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_208),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_381),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_223),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_238),
.B(n_2),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_395),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_240),
.B(n_2),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_258),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_269),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_299),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_304),
.B(n_5),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_207),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_302),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_317),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_344),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_309),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_360),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_353),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_214),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_323),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_331),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_336),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_337),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_347),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_350),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_351),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_209),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_362),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_214),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_236),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_209),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_236),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_212),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_212),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_318),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_215),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_296),
.B(n_6),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_221),
.B(n_6),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_215),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_363),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_304),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_304),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_218),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_365),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_218),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_318),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_375),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_219),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_375),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_208),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_315),
.B(n_12),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_219),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_360),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_372),
.B(n_12),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_404),
.B(n_13),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_210),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_368),
.Y(n_501)
);

INVxp33_ASAP7_75t_SL g502 ( 
.A(n_210),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_376),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_224),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_217),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_360),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_391),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_426),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_461),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_429),
.B(n_412),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_443),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_494),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_458),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_497),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_497),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_R g518 ( 
.A(n_422),
.B(n_432),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_482),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_435),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_507),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_414),
.B(n_392),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_455),
.B(n_360),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_439),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_448),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_417),
.B(n_217),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_411),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_455),
.B(n_260),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_434),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_229),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_438),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_454),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_457),
.Y(n_536)
);

HB1xp67_ASAP7_75t_L g537 ( 
.A(n_425),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_460),
.Y(n_538)
);

NOR2xp67_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_285),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_445),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_464),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_465),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_505),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_467),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_468),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_447),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_431),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_472),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_484),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_488),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_424),
.B(n_233),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_503),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_427),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_430),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_449),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_459),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_499),
.B(n_235),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_451),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_406),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_433),
.B(n_220),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_495),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_432),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_450),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_437),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_440),
.B(n_220),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_406),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_462),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_442),
.B(n_261),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_463),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_416),
.B(n_224),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_405),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_481),
.Y(n_578)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_473),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_441),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_416),
.B(n_244),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_419),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_485),
.B(n_285),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_442),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_444),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_444),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_419),
.B(n_247),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_486),
.B(n_203),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_R g589 ( 
.A(n_456),
.B(n_268),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_537),
.B(n_407),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_582),
.B(n_566),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_520),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_203),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_530),
.A2(n_413),
.B1(n_415),
.B2(n_409),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_582),
.B(n_566),
.Y(n_595)
);

INVx4_ASAP7_75t_SL g596 ( 
.A(n_523),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_523),
.B(n_226),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_519),
.B(n_420),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_582),
.B(n_456),
.Y(n_599)
);

OR2x6_ASAP7_75t_L g600 ( 
.A(n_523),
.B(n_226),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_530),
.B(n_548),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_582),
.B(n_471),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_537),
.B(n_407),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_585),
.Y(n_604)
);

AND3x2_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_312),
.C(n_246),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_584),
.B(n_408),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_569),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_519),
.B(n_420),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_582),
.B(n_471),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_512),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_566),
.B(n_475),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_421),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_566),
.B(n_475),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_557),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_557),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_561),
.A2(n_413),
.B1(n_415),
.B2(n_409),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_561),
.A2(n_502),
.B1(n_500),
.B2(n_428),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_558),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_512),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_581),
.B(n_477),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_558),
.Y(n_622)
);

AND3x4_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_408),
.C(n_231),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_509),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_583),
.A2(n_504),
.B1(n_496),
.B2(n_477),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_523),
.B(n_583),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_520),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_520),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_514),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_584),
.B(n_311),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_578),
.B(n_421),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_581),
.B(n_478),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_559),
.B(n_246),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_587),
.B(n_478),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_524),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_578),
.B(n_423),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_587),
.B(n_480),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_520),
.Y(n_639)
);

NAND3xp33_ASAP7_75t_L g640 ( 
.A(n_586),
.B(n_483),
.C(n_480),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_588),
.B(n_474),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_543),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_520),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_524),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_532),
.B(n_423),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_533),
.Y(n_646)
);

AND2x6_ASAP7_75t_L g647 ( 
.A(n_583),
.B(n_312),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g648 ( 
.A(n_518),
.B(n_483),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_532),
.B(n_576),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_510),
.B(n_487),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_589),
.B(n_573),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_559),
.B(n_487),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_543),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_510),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_527),
.B(n_319),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_516),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_527),
.A2(n_504),
.B1(n_496),
.B2(n_489),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_559),
.B(n_489),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_559),
.B(n_492),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_533),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_588),
.A2(n_559),
.B1(n_492),
.B2(n_562),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_559),
.B(n_476),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_524),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_588),
.B(n_479),
.Y(n_665)
);

AND3x2_ASAP7_75t_L g666 ( 
.A(n_563),
.B(n_328),
.C(n_319),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_533),
.B(n_311),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_588),
.B(n_250),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_533),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_533),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_538),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_516),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_526),
.Y(n_673)
);

INVx4_ASAP7_75t_SL g674 ( 
.A(n_538),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_538),
.Y(n_675)
);

INVx6_ASAP7_75t_L g676 ( 
.A(n_538),
.Y(n_676)
);

BUFx8_ASAP7_75t_SL g677 ( 
.A(n_577),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_517),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_538),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_562),
.A2(n_493),
.B1(n_491),
.B2(n_490),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_538),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_562),
.A2(n_345),
.B1(n_307),
.B2(n_382),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_222),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_569),
.B(n_222),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_526),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_517),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_541),
.Y(n_687)
);

AO22x2_ASAP7_75t_L g688 ( 
.A1(n_565),
.A2(n_567),
.B1(n_570),
.B2(n_564),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_575),
.Y(n_689)
);

BUFx4f_ASAP7_75t_L g690 ( 
.A(n_541),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_541),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_526),
.A2(n_354),
.B1(n_386),
.B2(n_390),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_579),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_580),
.B(n_231),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_541),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_511),
.B(n_253),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_541),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_541),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_528),
.B(n_234),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_546),
.A2(n_352),
.B1(n_357),
.B2(n_239),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_546),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_543),
.B(n_225),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_564),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_552),
.B(n_254),
.Y(n_704)
);

AND2x2_ASAP7_75t_SL g705 ( 
.A(n_571),
.B(n_328),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_515),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_552),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_543),
.B(n_553),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_548),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_546),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_521),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_553),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_521),
.Y(n_715)
);

INVx1_ASAP7_75t_SL g716 ( 
.A(n_560),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_552),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_511),
.B(n_255),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_553),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_525),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_525),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_529),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_529),
.Y(n_724)
);

BUFx6f_ASAP7_75t_SL g725 ( 
.A(n_565),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_553),
.B(n_225),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_574),
.A2(n_361),
.B1(n_324),
.B2(n_400),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_572),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_567),
.B(n_227),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_535),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_535),
.B(n_227),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_536),
.B(n_228),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_536),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_580),
.B(n_542),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_542),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_545),
.B(n_228),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_545),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_549),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_549),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_550),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_508),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_550),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_645),
.B(n_574),
.Y(n_743)
);

NOR2x1p5_ASAP7_75t_L g744 ( 
.A(n_640),
.B(n_531),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_610),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_607),
.B(n_570),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_619),
.Y(n_747)
);

AND2x2_ASAP7_75t_SL g748 ( 
.A(n_705),
.B(n_266),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_705),
.B(n_580),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_634),
.Y(n_750)
);

BUFx8_ASAP7_75t_L g751 ( 
.A(n_604),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_649),
.B(n_528),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_607),
.B(n_552),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_683),
.B(n_522),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_626),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_655),
.A2(n_556),
.B1(n_554),
.B2(n_551),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_652),
.B(n_230),
.Y(n_757)
);

NOR2xp67_ASAP7_75t_L g758 ( 
.A(n_718),
.B(n_551),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_634),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_659),
.B(n_598),
.Y(n_760)
);

NAND2xp33_ASAP7_75t_L g761 ( 
.A(n_593),
.B(n_311),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_634),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_630),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_632),
.A2(n_338),
.B1(n_334),
.B2(n_327),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_656),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_684),
.B(n_522),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_627),
.B(n_554),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_634),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_653),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_627),
.B(n_556),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_621),
.B(n_513),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_641),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_627),
.B(n_555),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_694),
.B(n_596),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_656),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_630),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_636),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_637),
.A2(n_349),
.B1(n_234),
.B2(n_245),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_592),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_627),
.B(n_734),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_655),
.A2(n_555),
.B1(n_539),
.B2(n_338),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_655),
.A2(n_539),
.B1(n_245),
.B2(n_324),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_621),
.B(n_534),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_672),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_627),
.B(n_230),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_627),
.B(n_232),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_672),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_678),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_678),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_686),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_686),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_596),
.B(n_544),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_624),
.B(n_232),
.Y(n_793)
);

NOR2x1_ASAP7_75t_L g794 ( 
.A(n_651),
.B(n_267),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_596),
.B(n_544),
.Y(n_795)
);

BUFx8_ASAP7_75t_L g796 ( 
.A(n_725),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_633),
.B(n_568),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_624),
.B(n_237),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_601),
.B(n_540),
.Y(n_799)
);

INVxp67_ASAP7_75t_SL g800 ( 
.A(n_662),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_644),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_655),
.A2(n_326),
.B1(n_349),
.B2(n_356),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_696),
.B(n_237),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_650),
.B(n_719),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_642),
.B(n_241),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_608),
.B(n_241),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_614),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_664),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_615),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_633),
.B(n_635),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_591),
.B(n_242),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_591),
.B(n_595),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_661),
.B(n_242),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_647),
.B(n_243),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_618),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_592),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_647),
.B(n_243),
.Y(n_817)
);

INVxp33_ASAP7_75t_L g818 ( 
.A(n_590),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_653),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_617),
.A2(n_327),
.B1(n_334),
.B2(n_326),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_673),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_647),
.B(n_252),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_647),
.B(n_252),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_685),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_R g825 ( 
.A(n_603),
.B(n_547),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_635),
.B(n_314),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_622),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_647),
.B(n_278),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_701),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_677),
.Y(n_830)
);

NAND2xp33_ASAP7_75t_L g831 ( 
.A(n_593),
.B(n_311),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_647),
.B(n_278),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_714),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_595),
.B(n_320),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_712),
.B(n_320),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_658),
.A2(n_276),
.B(n_398),
.C(n_389),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_706),
.B(n_314),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_599),
.B(n_321),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_638),
.B(n_348),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_715),
.B(n_321),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_721),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_710),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_722),
.B(n_340),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_641),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_641),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_723),
.B(n_340),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_724),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_730),
.B(n_341),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_697),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_733),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_638),
.B(n_348),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_735),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_655),
.A2(n_403),
.B1(n_401),
.B2(n_396),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_697),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_717),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_737),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_738),
.B(n_341),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_286),
.B(n_290),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_739),
.B(n_346),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_714),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_740),
.B(n_346),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_742),
.B(n_366),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_599),
.B(n_366),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_720),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_655),
.B(n_370),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_612),
.B(n_370),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_606),
.B(n_371),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_597),
.B(n_301),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_720),
.Y(n_869)
);

NAND2xp33_ASAP7_75t_L g870 ( 
.A(n_593),
.B(n_602),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_703),
.B(n_371),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_709),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_629),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_654),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_717),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_629),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_629),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_709),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_688),
.B(n_356),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_611),
.B(n_359),
.Y(n_880)
);

NOR2xp67_ASAP7_75t_L g881 ( 
.A(n_657),
.B(n_403),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_611),
.B(n_613),
.Y(n_882)
);

O2A1O1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_658),
.A2(n_316),
.B(n_369),
.C(n_373),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_716),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_676),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_602),
.B(n_393),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_688),
.B(n_393),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_688),
.B(n_396),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_613),
.B(n_401),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_592),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_639),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_597),
.B(n_322),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_625),
.B(n_359),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_639),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_597),
.B(n_361),
.Y(n_895)
);

BUFx12f_ASAP7_75t_SL g896 ( 
.A(n_597),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_600),
.B(n_364),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_665),
.B(n_364),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_639),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_609),
.B(n_257),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_609),
.B(n_259),
.Y(n_901)
);

NAND2x1p5_ASAP7_75t_L g902 ( 
.A(n_620),
.B(n_330),
.Y(n_902)
);

NOR3xp33_ASAP7_75t_L g903 ( 
.A(n_648),
.B(n_400),
.C(n_399),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_731),
.B(n_264),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_646),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_732),
.B(n_265),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_736),
.B(n_275),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_646),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_690),
.B(n_592),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_702),
.B(n_279),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_690),
.B(n_660),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_804),
.B(n_651),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_760),
.A2(n_631),
.B(n_690),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_810),
.A2(n_631),
.B(n_616),
.C(n_648),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_884),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_752),
.A2(n_727),
.B(n_726),
.C(n_729),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_779),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_748),
.B(n_623),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_804),
.B(n_600),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_760),
.A2(n_663),
.B(n_646),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_896),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_882),
.A2(n_594),
.B(n_663),
.C(n_713),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_812),
.A2(n_669),
.B(n_663),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_812),
.A2(n_670),
.B(n_669),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_800),
.B(n_600),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_780),
.A2(n_670),
.B(n_669),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_769),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_749),
.B(n_600),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_748),
.B(n_709),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_876),
.A2(n_671),
.B(n_670),
.Y(n_930)
);

O2A1O1Ixp33_ASAP7_75t_L g931 ( 
.A1(n_893),
.A2(n_699),
.B(n_668),
.C(n_713),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_749),
.B(n_668),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_743),
.A2(n_623),
.B1(n_741),
.B2(n_725),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_803),
.A2(n_679),
.B(n_713),
.C(n_707),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_745),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_807),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_876),
.A2(n_671),
.B(n_679),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_877),
.A2(n_671),
.B(n_679),
.Y(n_938)
);

BUFx12f_ASAP7_75t_L g939 ( 
.A(n_830),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_826),
.B(n_680),
.C(n_682),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_839),
.A2(n_707),
.B(n_695),
.C(n_681),
.Y(n_941)
);

OAI21x1_ASAP7_75t_L g942 ( 
.A1(n_902),
.A2(n_681),
.B(n_695),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_877),
.A2(n_695),
.B(n_681),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_769),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_891),
.A2(n_707),
.B(n_711),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_792),
.Y(n_946)
);

AOI21x1_ASAP7_75t_L g947 ( 
.A1(n_909),
.A2(n_704),
.B(n_378),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_880),
.A2(n_725),
.B1(n_593),
.B2(n_676),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_767),
.A2(n_770),
.B(n_773),
.Y(n_949)
);

BUFx12f_ASAP7_75t_L g950 ( 
.A(n_830),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_818),
.B(n_689),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_867),
.A2(n_628),
.B1(n_711),
.B2(n_675),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_779),
.B(n_816),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_818),
.B(n_693),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_851),
.A2(n_898),
.B(n_797),
.C(n_783),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_885),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_754),
.B(n_700),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_754),
.B(n_692),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_809),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_766),
.B(n_593),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_891),
.A2(n_620),
.B(n_711),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_766),
.B(n_728),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_792),
.B(n_605),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_795),
.B(n_666),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_771),
.A2(n_704),
.B(n_667),
.C(n_342),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_772),
.B(n_620),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_779),
.B(n_660),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_772),
.B(n_628),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_819),
.A2(n_698),
.B(n_691),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_820),
.A2(n_667),
.B(n_399),
.C(n_394),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_879),
.A2(n_593),
.B1(n_691),
.B2(n_687),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_746),
.B(n_628),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_779),
.B(n_816),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_844),
.B(n_643),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_779),
.B(n_660),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_774),
.B(n_643),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_816),
.B(n_660),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_815),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_833),
.A2(n_698),
.B(n_691),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_844),
.B(n_674),
.Y(n_980)
);

AO22x1_ASAP7_75t_L g981 ( 
.A1(n_751),
.A2(n_677),
.B1(n_394),
.B2(n_310),
.Y(n_981)
);

NAND2xp33_ASAP7_75t_L g982 ( 
.A(n_816),
.B(n_280),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_845),
.B(n_674),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_757),
.A2(n_282),
.B(n_287),
.C(n_288),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_795),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_811),
.A2(n_698),
.B(n_687),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_750),
.B(n_643),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_774),
.A2(n_676),
.B1(n_675),
.B2(n_687),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_827),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_811),
.A2(n_675),
.B(n_270),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_747),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_834),
.A2(n_374),
.B(n_297),
.Y(n_992)
);

INVx11_ASAP7_75t_L g993 ( 
.A(n_751),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_816),
.B(n_674),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_866),
.A2(n_303),
.B1(n_387),
.B2(n_385),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_879),
.A2(n_293),
.B1(n_295),
.B2(n_298),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_834),
.A2(n_271),
.B(n_383),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_751),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_905),
.A2(n_272),
.B(n_380),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_905),
.A2(n_283),
.B(n_284),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_902),
.A2(n_367),
.B(n_311),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_909),
.A2(n_911),
.B(n_757),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_911),
.A2(n_289),
.B(n_291),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_841),
.B(n_305),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_847),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_873),
.A2(n_292),
.B(n_300),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_765),
.A2(n_379),
.B(n_355),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_894),
.A2(n_313),
.B(n_402),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_845),
.B(n_306),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_850),
.B(n_308),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_799),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_764),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_860),
.A2(n_402),
.B1(n_248),
.B2(n_21),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_872),
.B(n_16),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_778),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_899),
.A2(n_402),
.B(n_248),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_896),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_852),
.B(n_20),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_874),
.B(n_22),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_860),
.A2(n_856),
.B1(n_756),
.B2(n_805),
.Y(n_1020)
);

OAI22x1_ASAP7_75t_L g1021 ( 
.A1(n_895),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_1021)
);

O2A1O1Ixp5_ASAP7_75t_L g1022 ( 
.A1(n_838),
.A2(n_311),
.B(n_367),
.C(n_33),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_908),
.A2(n_753),
.B(n_910),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_883),
.A2(n_402),
.B(n_248),
.C(n_34),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_802),
.B(n_402),
.C(n_248),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_775),
.A2(n_311),
.B(n_367),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_784),
.A2(n_311),
.B(n_367),
.Y(n_1027)
);

OAI21xp33_ASAP7_75t_L g1028 ( 
.A1(n_871),
.A2(n_248),
.B(n_32),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_806),
.A2(n_27),
.B(n_34),
.C(n_35),
.Y(n_1029)
);

INVxp67_ASAP7_75t_SL g1030 ( 
.A(n_750),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_758),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_885),
.Y(n_1032)
);

NOR3xp33_ASAP7_75t_L g1033 ( 
.A(n_806),
.B(n_41),
.C(n_45),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_904),
.B(n_46),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_838),
.A2(n_367),
.B(n_128),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_759),
.B(n_762),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_863),
.A2(n_367),
.B(n_123),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_890),
.B(n_367),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_906),
.B(n_46),
.Y(n_1039)
);

INVx1_ASAP7_75t_SL g1040 ( 
.A(n_837),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_863),
.A2(n_886),
.B(n_849),
.Y(n_1041)
);

BUFx12f_ASAP7_75t_L g1042 ( 
.A(n_796),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_787),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_1043)
);

AOI22x1_ASAP7_75t_L g1044 ( 
.A1(n_864),
.A2(n_367),
.B1(n_61),
.B2(n_62),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_788),
.A2(n_134),
.B(n_199),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_759),
.B(n_131),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_789),
.A2(n_137),
.B(n_196),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_892),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_890),
.B(n_50),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_790),
.A2(n_116),
.B(n_193),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_907),
.B(n_62),
.Y(n_1051)
);

BUFx4f_ASAP7_75t_L g1052 ( 
.A(n_872),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_890),
.B(n_63),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_SL g1054 ( 
.A(n_796),
.B(n_66),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_892),
.A2(n_67),
.B1(n_69),
.B2(n_75),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_892),
.A2(n_77),
.B1(n_85),
.B2(n_97),
.Y(n_1056)
);

OAI321xp33_ASAP7_75t_L g1057 ( 
.A1(n_781),
.A2(n_100),
.A3(n_107),
.B1(n_138),
.B2(n_139),
.C(n_140),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_791),
.A2(n_146),
.B(n_154),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_794),
.A2(n_163),
.B(n_166),
.C(n_169),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_886),
.A2(n_192),
.B(n_200),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_762),
.B(n_768),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_849),
.A2(n_875),
.B(n_855),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_854),
.A2(n_875),
.B(n_855),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_793),
.B(n_798),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_SL g1065 ( 
.A1(n_889),
.A2(n_869),
.B(n_900),
.C(n_901),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_768),
.B(n_890),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_881),
.A2(n_858),
.B(n_853),
.C(n_870),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_878),
.B(n_895),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_744),
.B(n_892),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_868),
.B(n_878),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_785),
.A2(n_786),
.B1(n_840),
.B2(n_859),
.Y(n_1071)
);

INVx2_ASAP7_75t_SL g1072 ( 
.A(n_837),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_796),
.Y(n_1073)
);

HB1xp67_ASAP7_75t_L g1074 ( 
.A(n_825),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_755),
.Y(n_1075)
);

O2A1O1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_835),
.A2(n_846),
.B(n_843),
.C(n_848),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_890),
.B(n_902),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_777),
.A2(n_824),
.B(n_821),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_763),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_868),
.B(n_862),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_857),
.A2(n_861),
.B1(n_813),
.B2(n_782),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_868),
.B(n_776),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_854),
.A2(n_870),
.B(n_776),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_777),
.A2(n_829),
.B(n_801),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_801),
.B(n_829),
.Y(n_1085)
);

AOI21x1_ASAP7_75t_L g1086 ( 
.A1(n_808),
.A2(n_824),
.B(n_842),
.Y(n_1086)
);

BUFx4f_ASAP7_75t_L g1087 ( 
.A(n_897),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_808),
.B(n_842),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_821),
.A2(n_865),
.B1(n_814),
.B2(n_817),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_897),
.B(n_888),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_887),
.B(n_822),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_823),
.B(n_828),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_L g1093 ( 
.A(n_832),
.B(n_903),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_761),
.A2(n_831),
.B(n_836),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_761),
.B(n_752),
.C(n_893),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1001),
.A2(n_831),
.B(n_1083),
.Y(n_1096)
);

AO31x2_ASAP7_75t_L g1097 ( 
.A1(n_941),
.A2(n_1089),
.A3(n_1091),
.B(n_1092),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_922),
.A2(n_1076),
.B(n_913),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_936),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_941),
.A2(n_1091),
.A3(n_1092),
.B(n_1071),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1064),
.A2(n_1081),
.B(n_924),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1095),
.B(n_955),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1041),
.A2(n_926),
.B(n_1002),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1020),
.A2(n_972),
.B(n_923),
.Y(n_1104)
);

AO21x1_ASAP7_75t_L g1105 ( 
.A1(n_1045),
.A2(n_1050),
.B(n_1047),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_918),
.A2(n_1068),
.B1(n_933),
.B2(n_962),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1086),
.A2(n_942),
.B(n_1062),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1063),
.A2(n_1084),
.B(n_1078),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_914),
.A2(n_916),
.B(n_918),
.C(n_912),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_920),
.A2(n_947),
.B(n_1023),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1011),
.B(n_958),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1011),
.B(n_932),
.Y(n_1112)
);

AOI21xp33_ASAP7_75t_L g1113 ( 
.A1(n_940),
.A2(n_1040),
.B(n_984),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1065),
.A2(n_934),
.B(n_945),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1065),
.A2(n_1039),
.B(n_1034),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_959),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_SL g1117 ( 
.A1(n_949),
.A2(n_1037),
.B(n_1035),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_993),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1051),
.A2(n_1094),
.B(n_937),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_931),
.A2(n_1067),
.B(n_1080),
.C(n_1028),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1012),
.A2(n_1015),
.B(n_1033),
.C(n_1029),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_917),
.B(n_1068),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1038),
.A2(n_1077),
.B(n_1027),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_SL g1124 ( 
.A1(n_1058),
.A2(n_925),
.B(n_1026),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_980),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_SL g1126 ( 
.A1(n_1060),
.A2(n_1018),
.B(n_960),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_953),
.A2(n_973),
.B(n_938),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_930),
.A2(n_943),
.B(n_961),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_1085),
.A2(n_1088),
.B(n_975),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1033),
.B(n_1031),
.C(n_1055),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_957),
.B(n_919),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_952),
.A2(n_977),
.B(n_967),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_967),
.A2(n_975),
.B(n_977),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_986),
.A2(n_969),
.B(n_979),
.Y(n_1134)
);

AO21x1_ASAP7_75t_L g1135 ( 
.A1(n_1049),
.A2(n_1053),
.B(n_1046),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1072),
.B(n_978),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_917),
.B(n_976),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_989),
.B(n_1005),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_SL g1139 ( 
.A1(n_1044),
.A2(n_1070),
.B(n_1056),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1074),
.B(n_929),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_1066),
.A2(n_994),
.B(n_1046),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_SL g1142 ( 
.A1(n_1090),
.A2(n_1007),
.B(n_948),
.Y(n_1142)
);

OR2x6_ASAP7_75t_L g1143 ( 
.A(n_998),
.B(n_1042),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1066),
.A2(n_994),
.B(n_1008),
.Y(n_1144)
);

NOR2x1_ASAP7_75t_SL g1145 ( 
.A(n_917),
.B(n_1082),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1074),
.B(n_929),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1075),
.A2(n_1079),
.B(n_1016),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_L g1148 ( 
.A1(n_1022),
.A2(n_1049),
.B(n_1053),
.C(n_1024),
.Y(n_1148)
);

INVx4_ASAP7_75t_L g1149 ( 
.A(n_939),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_985),
.B(n_928),
.Y(n_1150)
);

CKINVDCx20_ASAP7_75t_R g1151 ( 
.A(n_950),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_917),
.A2(n_990),
.B(n_974),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_946),
.B(n_1009),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1009),
.B(n_1030),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_983),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1087),
.B(n_954),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1024),
.A2(n_965),
.A3(n_1013),
.B(n_991),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_966),
.A2(n_974),
.B(n_968),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1087),
.B(n_951),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1030),
.B(n_915),
.Y(n_1160)
);

AOI21xp33_ASAP7_75t_L g1161 ( 
.A1(n_995),
.A2(n_970),
.B(n_996),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_966),
.A2(n_968),
.B(n_1057),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_996),
.A2(n_1010),
.B(n_1004),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1043),
.A2(n_1022),
.B(n_982),
.C(n_1014),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1036),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1093),
.A2(n_1000),
.B(n_999),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1006),
.A2(n_1052),
.B(n_971),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1014),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_987),
.A2(n_971),
.B(n_1061),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1048),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_1036),
.A2(n_1061),
.B(n_988),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1019),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1052),
.A2(n_927),
.B(n_944),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_927),
.A2(n_944),
.B(n_956),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_1073),
.Y(n_1175)
);

NAND2xp33_ASAP7_75t_SL g1176 ( 
.A(n_956),
.B(n_1032),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1032),
.A2(n_1069),
.B(n_1003),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_921),
.B(n_1017),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_921),
.Y(n_1179)
);

OAI21xp33_ASAP7_75t_L g1180 ( 
.A1(n_1054),
.A2(n_997),
.B(n_992),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1017),
.B(n_963),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1059),
.A2(n_1025),
.B(n_1021),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_964),
.A2(n_780),
.B(n_922),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_981),
.A2(n_955),
.B1(n_1095),
.B2(n_748),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1185)
);

OR2x6_ASAP7_75t_L g1186 ( 
.A(n_998),
.B(n_1042),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1095),
.B(n_955),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_980),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_962),
.B(n_752),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_935),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_955),
.B(n_804),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_918),
.A2(n_752),
.B1(n_748),
.B2(n_825),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_918),
.A2(n_893),
.B(n_530),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_962),
.B(n_752),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_L g1198 ( 
.A(n_1011),
.B(n_884),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_955),
.A2(n_882),
.B(n_810),
.C(n_1095),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_936),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_1011),
.B(n_985),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_955),
.B(n_804),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1011),
.B(n_985),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_922),
.A2(n_780),
.B(n_760),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_955),
.A2(n_1095),
.B1(n_748),
.B2(n_912),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1210)
);

AO221x2_ASAP7_75t_L g1211 ( 
.A1(n_1021),
.A2(n_1043),
.B1(n_1095),
.B2(n_940),
.C(n_820),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_962),
.B(n_752),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1040),
.B(n_706),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_993),
.Y(n_1217)
);

NOR2x1_ASAP7_75t_L g1218 ( 
.A(n_998),
.B(n_912),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_918),
.A2(n_893),
.B(n_530),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_922),
.A2(n_780),
.B(n_760),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_912),
.B(n_748),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_936),
.Y(n_1222)
);

AO21x2_ASAP7_75t_L g1223 ( 
.A1(n_1026),
.A2(n_1027),
.B(n_941),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_922),
.A2(n_780),
.B(n_760),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_915),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_955),
.B(n_804),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_955),
.B(n_804),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_955),
.B(n_804),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_955),
.A2(n_1095),
.B1(n_748),
.B2(n_912),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_962),
.B(n_752),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_962),
.B(n_752),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1011),
.B(n_985),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_SL g1241 ( 
.A1(n_1002),
.A2(n_1041),
.B(n_924),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_922),
.A2(n_780),
.B(n_760),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_955),
.A2(n_1095),
.B1(n_748),
.B2(n_912),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1001),
.A2(n_1083),
.B(n_1086),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_962),
.B(n_752),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1076),
.A2(n_760),
.B(n_1064),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_955),
.A2(n_1095),
.B(n_914),
.C(n_810),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1011),
.B(n_985),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_918),
.A2(n_752),
.B1(n_748),
.B2(n_825),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1099),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1227),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1181),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1214),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1143),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1194),
.A2(n_1249),
.B(n_1195),
.C(n_1219),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1105),
.A2(n_1189),
.B(n_1102),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_L g1258 ( 
.A(n_1200),
.B(n_1247),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1193),
.A2(n_1230),
.B1(n_1206),
.B2(n_1234),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1103),
.A2(n_1119),
.B(n_1098),
.Y(n_1261)
);

OR2x6_ASAP7_75t_SL g1262 ( 
.A(n_1184),
.B(n_1153),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1125),
.B(n_1155),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1116),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1151),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1203),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1156),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1221),
.B(n_1231),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1212),
.B(n_1236),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_L g1270 ( 
.A(n_1247),
.B(n_1121),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1109),
.B(n_1112),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1125),
.B(n_1155),
.Y(n_1272)
);

AND2x6_ASAP7_75t_SL g1273 ( 
.A(n_1143),
.B(n_1186),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1163),
.A2(n_1161),
.B(n_1130),
.C(n_1164),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1102),
.A2(n_1189),
.B(n_1158),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1121),
.A2(n_1243),
.B(n_1235),
.C(n_1209),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1118),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1190),
.B(n_1159),
.Y(n_1278)
);

CKINVDCx20_ASAP7_75t_R g1279 ( 
.A(n_1217),
.Y(n_1279)
);

OR2x4_ASAP7_75t_L g1280 ( 
.A(n_1178),
.B(n_1172),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1187),
.B(n_1188),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1160),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1158),
.A2(n_1124),
.B(n_1104),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1162),
.A2(n_1134),
.B(n_1101),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_1138),
.B1(n_1245),
.B2(n_1238),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1143),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1205),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1186),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1222),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1115),
.A2(n_1117),
.B(n_1119),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_SL g1291 ( 
.A(n_1149),
.B(n_1186),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_1190),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1211),
.A2(n_1154),
.B1(n_1111),
.B2(n_1113),
.Y(n_1293)
);

A2O1A1Ixp33_ASAP7_75t_SL g1294 ( 
.A1(n_1115),
.A2(n_1166),
.B(n_1237),
.C(n_1229),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1205),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1187),
.B(n_1188),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1140),
.B(n_1146),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1218),
.B(n_1169),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_SL g1299 ( 
.A(n_1173),
.B(n_1183),
.Y(n_1299)
);

OA22x2_ASAP7_75t_L g1300 ( 
.A1(n_1168),
.A2(n_1170),
.B1(n_1248),
.B2(n_1207),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1199),
.B(n_1202),
.Y(n_1301)
);

HB1xp67_ASAP7_75t_L g1302 ( 
.A(n_1136),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1134),
.A2(n_1162),
.B(n_1128),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1211),
.A2(n_1248),
.B1(n_1239),
.B2(n_1207),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1128),
.A2(n_1246),
.B(n_1199),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1175),
.A2(n_1149),
.B1(n_1178),
.B2(n_1179),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1239),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1202),
.A2(n_1246),
.B(n_1213),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1175),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1210),
.B(n_1213),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1198),
.B(n_1150),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1210),
.A2(n_1226),
.B(n_1216),
.Y(n_1312)
);

OR2x2_ASAP7_75t_SL g1313 ( 
.A(n_1165),
.B(n_1182),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1122),
.B(n_1216),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1122),
.B(n_1225),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1142),
.A2(n_1180),
.B1(n_1135),
.B2(n_1139),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1225),
.B(n_1240),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1226),
.B(n_1240),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1177),
.Y(n_1319)
);

INVx4_ASAP7_75t_SL g1320 ( 
.A(n_1157),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1229),
.B(n_1237),
.Y(n_1321)
);

OR2x6_ASAP7_75t_L g1322 ( 
.A(n_1173),
.B(n_1167),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1145),
.B(n_1100),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1100),
.B(n_1208),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_L g1325 ( 
.A(n_1166),
.B(n_1167),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1120),
.B(n_1220),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1224),
.B(n_1242),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1164),
.B(n_1126),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1137),
.Y(n_1329)
);

BUFx3_ASAP7_75t_L g1330 ( 
.A(n_1174),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1141),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1114),
.A2(n_1132),
.A3(n_1171),
.B(n_1152),
.Y(n_1332)
);

CKINVDCx8_ASAP7_75t_R g1333 ( 
.A(n_1176),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1132),
.A2(n_1137),
.B1(n_1114),
.B2(n_1152),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1129),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1100),
.B(n_1097),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1133),
.B(n_1144),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1223),
.A2(n_1241),
.B(n_1096),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1223),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1157),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1148),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1127),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1157),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1157),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1147),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1097),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1148),
.A2(n_1097),
.B1(n_1123),
.B2(n_1110),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1108),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1107),
.B(n_1185),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1197),
.A2(n_1244),
.B(n_1204),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1201),
.B(n_1215),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1233),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1228),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1232),
.A2(n_1105),
.B(n_1102),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1099),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1099),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1214),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1099),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1143),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1195),
.A2(n_748),
.B1(n_940),
.B2(n_705),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1192),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1105),
.A2(n_1158),
.B(n_1102),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1195),
.A2(n_748),
.B1(n_940),
.B2(n_705),
.Y(n_1365)
);

INVx5_ASAP7_75t_L g1366 ( 
.A(n_1125),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1193),
.A2(n_1039),
.B(n_1034),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1227),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1105),
.A2(n_1189),
.B(n_1102),
.Y(n_1371)
);

INVx3_ASAP7_75t_SL g1372 ( 
.A(n_1143),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1194),
.A2(n_955),
.B(n_1095),
.C(n_1249),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1105),
.A2(n_1189),
.B(n_1102),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1143),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1099),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1194),
.A2(n_1249),
.B1(n_955),
.B2(n_1095),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1200),
.A2(n_955),
.B(n_1247),
.C(n_1219),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1194),
.A2(n_1249),
.B1(n_918),
.B2(n_748),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_1160),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1125),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_SL g1389 ( 
.A1(n_1098),
.A2(n_606),
.B(n_659),
.C(n_652),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1194),
.B(n_1249),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1393)
);

AO32x1_ASAP7_75t_L g1394 ( 
.A1(n_1184),
.A2(n_1209),
.A3(n_1243),
.B1(n_1235),
.B2(n_1043),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1105),
.A2(n_1189),
.B(n_1102),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1143),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1227),
.Y(n_1397)
);

OAI221xp5_ASAP7_75t_L g1398 ( 
.A1(n_1194),
.A2(n_955),
.B1(n_1249),
.B2(n_752),
.C(n_1219),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1194),
.A2(n_955),
.B(n_1095),
.C(n_1249),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1105),
.A2(n_1189),
.B(n_1102),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1191),
.B(n_1196),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1105),
.A2(n_1189),
.B(n_1102),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1221),
.B(n_1131),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1099),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1398),
.A2(n_1382),
.B1(n_1285),
.B2(n_1341),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1336),
.B(n_1324),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1265),
.Y(n_1409)
);

NAND2x1p5_ASAP7_75t_L g1410 ( 
.A(n_1299),
.B(n_1292),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1250),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1279),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1264),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1350),
.A2(n_1303),
.B(n_1338),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1266),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1303),
.A2(n_1305),
.B(n_1283),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1289),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1251),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1350),
.A2(n_1305),
.B(n_1308),
.Y(n_1419)
);

BUFx2_ASAP7_75t_R g1420 ( 
.A(n_1372),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1355),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1282),
.Y(n_1422)
);

AOI21xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1306),
.A2(n_1276),
.B(n_1285),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1392),
.A2(n_1361),
.B1(n_1365),
.B2(n_1384),
.Y(n_1424)
);

AO21x1_ASAP7_75t_L g1425 ( 
.A1(n_1382),
.A2(n_1270),
.B(n_1383),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1356),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1358),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1322),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1346),
.B(n_1268),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1360),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1398),
.A2(n_1293),
.B1(n_1300),
.B2(n_1362),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1381),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1277),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1300),
.A2(n_1362),
.B1(n_1370),
.B2(n_1373),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1375),
.A2(n_1399),
.B1(n_1280),
.B2(n_1333),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1343),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1268),
.B(n_1314),
.Y(n_1437)
);

INVxp33_ASAP7_75t_L g1438 ( 
.A(n_1368),
.Y(n_1438)
);

BUFx2_ASAP7_75t_SL g1439 ( 
.A(n_1360),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1309),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1335),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1277),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1344),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1315),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1280),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1406),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1259),
.B(n_1370),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1281),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1253),
.B(n_1269),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1281),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1296),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1259),
.A2(n_1405),
.B1(n_1373),
.B2(n_1374),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1369),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1322),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1258),
.A2(n_1405),
.B1(n_1402),
.B2(n_1393),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1330),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1322),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1374),
.A2(n_1385),
.B1(n_1402),
.B2(n_1393),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1380),
.B(n_1385),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1380),
.B(n_1297),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1312),
.A2(n_1284),
.B(n_1354),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1292),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1274),
.A2(n_1256),
.B1(n_1262),
.B2(n_1271),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1376),
.A2(n_1388),
.B1(n_1378),
.B2(n_1401),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1325),
.A2(n_1354),
.B(n_1364),
.Y(n_1465)
);

INVx1_ASAP7_75t_SL g1466 ( 
.A(n_1254),
.Y(n_1466)
);

BUFx8_ASAP7_75t_SL g1467 ( 
.A(n_1397),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1317),
.B(n_1390),
.Y(n_1468)
);

AOI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1312),
.A2(n_1404),
.B(n_1400),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1260),
.A2(n_1326),
.B1(n_1271),
.B2(n_1311),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1391),
.A2(n_1403),
.B1(n_1359),
.B2(n_1363),
.Y(n_1471)
);

OAI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1304),
.A2(n_1291),
.B1(n_1252),
.B2(n_1328),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1337),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1302),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1275),
.A2(n_1257),
.B1(n_1371),
.B2(n_1395),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1273),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1257),
.A2(n_1371),
.B(n_1377),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1334),
.A2(n_1347),
.B(n_1275),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1386),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1347),
.A2(n_1395),
.B(n_1377),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1323),
.B(n_1320),
.Y(n_1481)
);

INVxp67_ASAP7_75t_L g1482 ( 
.A(n_1295),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_SL g1483 ( 
.A(n_1286),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1260),
.A2(n_1287),
.B1(n_1267),
.B2(n_1307),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1296),
.A2(n_1321),
.B(n_1310),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1329),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1301),
.A2(n_1321),
.B(n_1318),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1313),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1320),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1255),
.A2(n_1396),
.B1(n_1379),
.B2(n_1288),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1327),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1327),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1357),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_1278),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1394),
.A2(n_1278),
.B1(n_1292),
.B2(n_1366),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1301),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1310),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1318),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1263),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1272),
.Y(n_1500)
);

INVx3_ASAP7_75t_L g1501 ( 
.A(n_1342),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1320),
.B(n_1261),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1298),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1345),
.A2(n_1294),
.B(n_1352),
.Y(n_1504)
);

INVx6_ASAP7_75t_L g1505 ( 
.A(n_1292),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1339),
.A2(n_1387),
.B1(n_1366),
.B2(n_1316),
.Y(n_1506)
);

CKINVDCx11_ASAP7_75t_R g1507 ( 
.A(n_1331),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1366),
.B(n_1387),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1366),
.B(n_1387),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1334),
.A2(n_1319),
.B(n_1367),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1394),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1331),
.A2(n_1389),
.B1(n_1290),
.B2(n_1319),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1332),
.B(n_1290),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1351),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1348),
.Y(n_1515)
);

INVx6_ASAP7_75t_L g1516 ( 
.A(n_1349),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1353),
.A2(n_748),
.B1(n_1211),
.B2(n_601),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1274),
.A2(n_955),
.B(n_1095),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1350),
.A2(n_1303),
.B(n_1338),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1322),
.Y(n_1520)
);

AO21x1_ASAP7_75t_SL g1521 ( 
.A1(n_1316),
.A2(n_1296),
.B(n_1281),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1259),
.B(n_1191),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1340),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1251),
.Y(n_1524)
);

INVxp33_ASAP7_75t_L g1525 ( 
.A(n_1368),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1384),
.A2(n_1249),
.B1(n_1194),
.B2(n_601),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1350),
.A2(n_1303),
.B(n_1338),
.Y(n_1527)
);

AO21x1_ASAP7_75t_L g1528 ( 
.A1(n_1382),
.A2(n_1392),
.B(n_1276),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1336),
.B(n_1324),
.Y(n_1529)
);

BUFx8_ASAP7_75t_SL g1530 ( 
.A(n_1265),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1336),
.B(n_1324),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1250),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1259),
.B(n_1191),
.Y(n_1533)
);

NOR2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1360),
.B(n_998),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1250),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1250),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_SL g1537 ( 
.A1(n_1276),
.A2(n_1383),
.B(n_1283),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1335),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1335),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1265),
.Y(n_1540)
);

NAND2x1p5_ASAP7_75t_L g1541 ( 
.A(n_1299),
.B(n_1169),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1392),
.A2(n_748),
.B1(n_1219),
.B2(n_1195),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1449),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1523),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1468),
.B(n_1437),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1419),
.A2(n_1519),
.B(n_1414),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1496),
.B(n_1497),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_L g1549 ( 
.A(n_1428),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1468),
.B(n_1437),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1420),
.B(n_1409),
.Y(n_1551)
);

CKINVDCx14_ASAP7_75t_R g1552 ( 
.A(n_1409),
.Y(n_1552)
);

INVx4_ASAP7_75t_L g1553 ( 
.A(n_1507),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1408),
.B(n_1529),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1422),
.Y(n_1555)
);

AOI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1469),
.A2(n_1475),
.B(n_1487),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1429),
.B(n_1408),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1507),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1460),
.B(n_1447),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1530),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1486),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1531),
.B(n_1444),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1527),
.A2(n_1469),
.B(n_1510),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1460),
.B(n_1459),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1458),
.B(n_1452),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1514),
.Y(n_1567)
);

INVxp67_ASAP7_75t_SL g1568 ( 
.A(n_1479),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1444),
.B(n_1454),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1429),
.B(n_1448),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1418),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1463),
.A2(n_1435),
.B1(n_1537),
.B2(n_1518),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1454),
.B(n_1520),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1498),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1540),
.B(n_1530),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1448),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1450),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1485),
.Y(n_1578)
);

AO21x2_ASAP7_75t_L g1579 ( 
.A1(n_1537),
.A2(n_1511),
.B(n_1526),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1520),
.B(n_1521),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1524),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1450),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1467),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1540),
.B(n_1412),
.Y(n_1584)
);

OR2x6_ASAP7_75t_L g1585 ( 
.A(n_1489),
.B(n_1481),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1478),
.A2(n_1487),
.B(n_1541),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1445),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1451),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1451),
.B(n_1485),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1485),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1436),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1436),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1516),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1412),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1474),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1521),
.B(n_1473),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1514),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1443),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1443),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1477),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1514),
.B(n_1457),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1477),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1455),
.B(n_1522),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1493),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1513),
.B(n_1457),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1457),
.B(n_1516),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1411),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1413),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1415),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1516),
.B(n_1480),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_1442),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1417),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1533),
.B(n_1434),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1421),
.Y(n_1614)
);

CKINVDCx20_ASAP7_75t_R g1615 ( 
.A(n_1467),
.Y(n_1615)
);

BUFx3_ASAP7_75t_L g1616 ( 
.A(n_1488),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1426),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1427),
.B(n_1432),
.Y(n_1618)
);

OA21x2_ASAP7_75t_L g1619 ( 
.A1(n_1515),
.A2(n_1425),
.B(n_1528),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1446),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1532),
.B(n_1535),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1441),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1536),
.Y(n_1623)
);

OA21x2_ASAP7_75t_L g1624 ( 
.A1(n_1515),
.A2(n_1425),
.B(n_1528),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1491),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_R g1626 ( 
.A(n_1442),
.B(n_1433),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1492),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1517),
.A2(n_1407),
.B1(n_1424),
.B2(n_1542),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1482),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1502),
.B(n_1416),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1441),
.B(n_1539),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1416),
.A2(n_1461),
.B(n_1410),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1441),
.B(n_1539),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1493),
.Y(n_1635)
);

AO21x1_ASAP7_75t_SL g1636 ( 
.A1(n_1506),
.A2(n_1431),
.B(n_1503),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1504),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1504),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1499),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1544),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1578),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1548),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1548),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1545),
.B(n_1416),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1545),
.B(n_1461),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1544),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1552),
.B(n_1453),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1546),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1550),
.B(n_1461),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1546),
.Y(n_1652)
);

BUFx2_ASAP7_75t_SL g1653 ( 
.A(n_1559),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1556),
.A2(n_1564),
.B(n_1547),
.Y(n_1654)
);

INVx1_ASAP7_75t_SL g1655 ( 
.A(n_1631),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1610),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1550),
.B(n_1465),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1590),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1554),
.B(n_1558),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1632),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1634),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1554),
.B(n_1465),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1568),
.B(n_1470),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1557),
.B(n_1538),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_SL g1665 ( 
.A1(n_1566),
.A2(n_1476),
.B1(n_1423),
.B2(n_1494),
.Y(n_1665)
);

OR2x6_ASAP7_75t_L g1666 ( 
.A(n_1585),
.B(n_1538),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_L g1667 ( 
.A(n_1553),
.B(n_1456),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1632),
.A2(n_1484),
.B(n_1508),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1586),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1628),
.A2(n_1476),
.B1(n_1471),
.B2(n_1472),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1572),
.A2(n_1525),
.B1(n_1438),
.B2(n_1464),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1603),
.A2(n_1494),
.B1(n_1505),
.B2(n_1495),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1619),
.A2(n_1410),
.B(n_1512),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1557),
.B(n_1589),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1558),
.B(n_1501),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1559),
.Y(n_1676)
);

INVx2_ASAP7_75t_SL g1677 ( 
.A(n_1634),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1630),
.B(n_1410),
.Y(n_1678)
);

NAND3xp33_ASAP7_75t_L g1679 ( 
.A(n_1619),
.B(n_1500),
.C(n_1453),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1589),
.B(n_1440),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1586),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1634),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1590),
.Y(n_1683)
);

BUFx3_ASAP7_75t_L g1684 ( 
.A(n_1559),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1630),
.B(n_1462),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1570),
.B(n_1466),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1549),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1570),
.B(n_1439),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1574),
.B(n_1439),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1563),
.B(n_1462),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1613),
.A2(n_1534),
.B1(n_1483),
.B2(n_1490),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1692)
);

NAND3xp33_ASAP7_75t_L g1693 ( 
.A(n_1642),
.B(n_1587),
.C(n_1562),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1667),
.B(n_1580),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1654),
.A2(n_1602),
.B(n_1600),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_L g1696 ( 
.A(n_1642),
.B(n_1592),
.C(n_1591),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1647),
.B(n_1575),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1659),
.B(n_1555),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.B(n_1596),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1659),
.B(n_1581),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1659),
.B(n_1680),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1641),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1680),
.B(n_1560),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1662),
.B(n_1580),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1674),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1657),
.B(n_1573),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1643),
.B(n_1598),
.C(n_1599),
.Y(n_1707)
);

NAND3xp33_ASAP7_75t_L g1708 ( 
.A(n_1643),
.B(n_1598),
.C(n_1599),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1680),
.B(n_1565),
.Y(n_1709)
);

OAI211xp5_ASAP7_75t_L g1710 ( 
.A1(n_1665),
.A2(n_1571),
.B(n_1553),
.C(n_1629),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1657),
.B(n_1595),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_SL g1712 ( 
.A(n_1663),
.B(n_1561),
.C(n_1611),
.Y(n_1712)
);

OAI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1665),
.A2(n_1616),
.B1(n_1551),
.B2(n_1612),
.C(n_1608),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1672),
.A2(n_1553),
.B1(n_1604),
.B2(n_1635),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1667),
.B(n_1593),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1672),
.A2(n_1553),
.B1(n_1543),
.B2(n_1594),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1663),
.B(n_1619),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1689),
.A2(n_1607),
.B(n_1639),
.C(n_1625),
.Y(n_1718)
);

NAND4xp25_ASAP7_75t_L g1719 ( 
.A(n_1689),
.B(n_1671),
.C(n_1651),
.D(n_1650),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_SL g1720 ( 
.A1(n_1679),
.A2(n_1624),
.B1(n_1619),
.B2(n_1673),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1657),
.B(n_1618),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1644),
.B(n_1645),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1653),
.B(n_1626),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1644),
.B(n_1618),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1691),
.A2(n_1583),
.B(n_1584),
.Y(n_1725)
);

NAND3xp33_ASAP7_75t_L g1726 ( 
.A(n_1679),
.B(n_1592),
.C(n_1591),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1644),
.B(n_1621),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_L g1728 ( 
.A(n_1658),
.B(n_1625),
.C(n_1627),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1687),
.B(n_1593),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1645),
.B(n_1621),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1645),
.B(n_1563),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1670),
.A2(n_1601),
.B1(n_1624),
.B2(n_1627),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1676),
.B(n_1626),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1649),
.B(n_1573),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1649),
.B(n_1605),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1686),
.A2(n_1614),
.B1(n_1617),
.B2(n_1608),
.C(n_1620),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1691),
.A2(n_1606),
.B(n_1633),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1658),
.B(n_1624),
.C(n_1574),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1649),
.B(n_1576),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1675),
.B(n_1605),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1671),
.A2(n_1579),
.B1(n_1616),
.B2(n_1624),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1675),
.B(n_1606),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1686),
.B(n_1576),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1673),
.A2(n_1633),
.B(n_1631),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1653),
.A2(n_1601),
.B1(n_1567),
.B2(n_1597),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1683),
.B(n_1638),
.C(n_1637),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1674),
.B(n_1577),
.Y(n_1747)
);

OAI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1668),
.A2(n_1616),
.B1(n_1609),
.B2(n_1620),
.C(n_1623),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1676),
.B(n_1433),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1675),
.B(n_1569),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1685),
.B(n_1682),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1674),
.B(n_1577),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1688),
.B(n_1582),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_SL g1754 ( 
.A(n_1661),
.B(n_1615),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1685),
.B(n_1569),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1688),
.B(n_1582),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1655),
.B(n_1588),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1717),
.B(n_1683),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1705),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1735),
.B(n_1692),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1695),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1717),
.A2(n_1636),
.B1(n_1579),
.B2(n_1668),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1728),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1739),
.B(n_1640),
.Y(n_1764)
);

INVx3_ASAP7_75t_L g1765 ( 
.A(n_1695),
.Y(n_1765)
);

AND2x4_ASAP7_75t_SL g1766 ( 
.A(n_1740),
.B(n_1666),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1692),
.B(n_1682),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1695),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1711),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1736),
.B(n_1640),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1722),
.B(n_1724),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1699),
.B(n_1685),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1747),
.B(n_1646),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1699),
.B(n_1678),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1752),
.B(n_1646),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1757),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1723),
.B(n_1666),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1753),
.B(n_1648),
.Y(n_1778)
);

AND2x2_ASAP7_75t_SL g1779 ( 
.A(n_1741),
.B(n_1650),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1756),
.B(n_1648),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1702),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1696),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1704),
.B(n_1678),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1727),
.B(n_1730),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1732),
.A2(n_1636),
.B1(n_1579),
.B2(n_1668),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1738),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1707),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1704),
.B(n_1678),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1706),
.B(n_1690),
.Y(n_1789)
);

NAND3xp33_ASAP7_75t_L g1790 ( 
.A(n_1720),
.B(n_1612),
.C(n_1609),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1708),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1706),
.B(n_1690),
.Y(n_1792)
);

AND2x4_ASAP7_75t_L g1793 ( 
.A(n_1740),
.B(n_1666),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1721),
.B(n_1652),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1743),
.B(n_1652),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1701),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1734),
.B(n_1690),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1734),
.B(n_1661),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1726),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1731),
.B(n_1651),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1746),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1698),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1751),
.B(n_1661),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1751),
.B(n_1666),
.Y(n_1804)
);

INVxp67_ASAP7_75t_SL g1805 ( 
.A(n_1748),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1750),
.B(n_1677),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1694),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1755),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1719),
.B(n_1703),
.Y(n_1809)
);

OR2x6_ASAP7_75t_L g1810 ( 
.A(n_1790),
.B(n_1737),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1795),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1782),
.B(n_1787),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1771),
.B(n_1700),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1779),
.A2(n_1716),
.B1(n_1714),
.B2(n_1713),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1771),
.B(n_1709),
.Y(n_1815)
);

BUFx2_ASAP7_75t_L g1816 ( 
.A(n_1782),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1787),
.B(n_1718),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1771),
.B(n_1664),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1795),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1765),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1778),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1778),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1780),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1793),
.B(n_1676),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1784),
.B(n_1664),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1760),
.B(n_1755),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1780),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1766),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1765),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1793),
.B(n_1684),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1799),
.A2(n_1710),
.B(n_1725),
.C(n_1744),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1770),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1760),
.B(n_1793),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1793),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1760),
.B(n_1742),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1763),
.B(n_1693),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1765),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1799),
.A2(n_1754),
.B(n_1694),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1763),
.B(n_1750),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1784),
.B(n_1664),
.Y(n_1840)
);

NOR2x1p5_ASAP7_75t_SL g1841 ( 
.A(n_1761),
.B(n_1600),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1770),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1784),
.B(n_1742),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1793),
.B(n_1684),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1759),
.B(n_1677),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1786),
.B(n_1801),
.C(n_1805),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1773),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1765),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1791),
.B(n_1614),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1791),
.B(n_1697),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1802),
.B(n_1677),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1802),
.B(n_1656),
.Y(n_1852)
);

OAI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1790),
.A2(n_1712),
.B(n_1754),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1849),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1833),
.B(n_1807),
.Y(n_1855)
);

OAI21xp33_ASAP7_75t_SL g1856 ( 
.A1(n_1810),
.A2(n_1779),
.B(n_1807),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1811),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1812),
.B(n_1810),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1819),
.Y(n_1859)
);

NOR2x1_ASAP7_75t_L g1860 ( 
.A(n_1846),
.B(n_1801),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1833),
.B(n_1805),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1821),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1816),
.B(n_1786),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1835),
.B(n_1826),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1832),
.B(n_1809),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1822),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1828),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1835),
.B(n_1807),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1823),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1826),
.B(n_1789),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1827),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1810),
.A2(n_1779),
.B1(n_1785),
.B2(n_1762),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1842),
.B(n_1809),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1820),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1850),
.B(n_1809),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1843),
.B(n_1815),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1850),
.B(n_1836),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1817),
.B(n_1769),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1847),
.B(n_1769),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1824),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1839),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1825),
.Y(n_1882)
);

NOR2x1_ASAP7_75t_R g1883 ( 
.A(n_1824),
.B(n_1684),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1813),
.B(n_1758),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1828),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1844),
.B(n_1789),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1831),
.B(n_1758),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1845),
.Y(n_1888)
);

NOR2x1p5_ASAP7_75t_L g1889 ( 
.A(n_1834),
.B(n_1759),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1844),
.B(n_1789),
.Y(n_1890)
);

INVx3_ASAP7_75t_L g1891 ( 
.A(n_1824),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1838),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1830),
.B(n_1853),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1840),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1831),
.B(n_1776),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1834),
.B(n_1830),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1818),
.B(n_1776),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1820),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1829),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1864),
.B(n_1830),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1857),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1872),
.A2(n_1785),
.B1(n_1762),
.B2(n_1814),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1860),
.B(n_1837),
.C(n_1829),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1860),
.A2(n_1768),
.B1(n_1761),
.B2(n_1765),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1877),
.B(n_1852),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1875),
.B(n_1796),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1868),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1895),
.B(n_1796),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1892),
.Y(n_1909)
);

NOR2x1_ASAP7_75t_L g1910 ( 
.A(n_1858),
.B(n_1837),
.Y(n_1910)
);

BUFx3_ASAP7_75t_L g1911 ( 
.A(n_1867),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1857),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1864),
.B(n_1792),
.Y(n_1913)
);

INVx1_ASAP7_75t_SL g1914 ( 
.A(n_1858),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1889),
.B(n_1834),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1859),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1870),
.B(n_1792),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1859),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1856),
.A2(n_1777),
.B1(n_1848),
.B2(n_1761),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1868),
.Y(n_1920)
);

CKINVDCx16_ASAP7_75t_R g1921 ( 
.A(n_1893),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1893),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1876),
.B(n_1773),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1863),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1870),
.B(n_1792),
.Y(n_1925)
);

INVxp67_ASAP7_75t_SL g1926 ( 
.A(n_1878),
.Y(n_1926)
);

INVx1_ASAP7_75t_SL g1927 ( 
.A(n_1867),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1855),
.B(n_1797),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1876),
.B(n_1775),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1889),
.B(n_1848),
.Y(n_1930)
);

AOI222xp33_ASAP7_75t_L g1931 ( 
.A1(n_1887),
.A2(n_1841),
.B1(n_1768),
.B2(n_1656),
.C1(n_1781),
.C2(n_1777),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1862),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1862),
.Y(n_1933)
);

INVxp67_ASAP7_75t_L g1934 ( 
.A(n_1885),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1866),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1898),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1855),
.B(n_1797),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1921),
.B(n_1861),
.Y(n_1938)
);

OAI222xp33_ASAP7_75t_L g1939 ( 
.A1(n_1902),
.A2(n_1873),
.B1(n_1865),
.B2(n_1861),
.C1(n_1856),
.C2(n_1885),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1914),
.B(n_1881),
.Y(n_1940)
);

AOI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1909),
.A2(n_1861),
.B1(n_1854),
.B2(n_1866),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1901),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1921),
.B(n_1861),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1909),
.A2(n_1931),
.B1(n_1919),
.B2(n_1903),
.Y(n_1944)
);

O2A1O1Ixp33_ASAP7_75t_L g1945 ( 
.A1(n_1903),
.A2(n_1888),
.B(n_1869),
.C(n_1871),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1926),
.B(n_1854),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1900),
.B(n_1880),
.Y(n_1947)
);

NOR3xp33_ASAP7_75t_L g1948 ( 
.A(n_1924),
.B(n_1891),
.C(n_1880),
.Y(n_1948)
);

OAI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1919),
.A2(n_1891),
.B1(n_1880),
.B2(n_1884),
.Y(n_1949)
);

OAI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1904),
.A2(n_1891),
.B1(n_1880),
.B2(n_1896),
.Y(n_1950)
);

NOR3xp33_ASAP7_75t_L g1951 ( 
.A(n_1922),
.B(n_1891),
.C(n_1871),
.Y(n_1951)
);

OAI221xp5_ASAP7_75t_L g1952 ( 
.A1(n_1908),
.A2(n_1869),
.B1(n_1768),
.B2(n_1879),
.C(n_1894),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1927),
.B(n_1882),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1905),
.B(n_1882),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1907),
.A2(n_1896),
.B1(n_1894),
.B2(n_1890),
.Y(n_1955)
);

OAI33xp33_ASAP7_75t_L g1956 ( 
.A1(n_1934),
.A2(n_1901),
.A3(n_1912),
.B1(n_1935),
.B2(n_1933),
.B3(n_1932),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1907),
.A2(n_1896),
.B1(n_1890),
.B2(n_1886),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1900),
.B(n_1886),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1920),
.B(n_1928),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1920),
.B(n_1896),
.Y(n_1960)
);

AOI21xp33_ASAP7_75t_L g1961 ( 
.A1(n_1910),
.A2(n_1874),
.B(n_1898),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1911),
.B(n_1884),
.Y(n_1962)
);

OAI22xp33_ASAP7_75t_SL g1963 ( 
.A1(n_1910),
.A2(n_1899),
.B1(n_1898),
.B2(n_1874),
.Y(n_1963)
);

AOI311xp33_ASAP7_75t_L g1964 ( 
.A1(n_1912),
.A2(n_1800),
.A3(n_1733),
.B(n_1897),
.C(n_1749),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1911),
.B(n_1883),
.Y(n_1965)
);

INVx1_ASAP7_75t_SL g1966 ( 
.A(n_1938),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1963),
.B(n_1915),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1944),
.A2(n_1937),
.B1(n_1928),
.B2(n_1923),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1956),
.A2(n_1936),
.B1(n_1918),
.B2(n_1935),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1942),
.Y(n_1970)
);

NOR2xp33_ASAP7_75t_L g1971 ( 
.A(n_1943),
.B(n_1916),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1940),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1938),
.B(n_1937),
.Y(n_1973)
);

NAND2x1p5_ASAP7_75t_L g1974 ( 
.A(n_1943),
.B(n_1915),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1953),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1959),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1946),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1958),
.B(n_1913),
.Y(n_1978)
);

NAND3xp33_ASAP7_75t_L g1979 ( 
.A(n_1948),
.B(n_1918),
.C(n_1916),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1951),
.B(n_1913),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1954),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1947),
.B(n_1960),
.Y(n_1982)
);

OR2x2_ASAP7_75t_L g1983 ( 
.A(n_1962),
.B(n_1923),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1949),
.B(n_1915),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1941),
.B(n_1917),
.Y(n_1985)
);

INVxp67_ASAP7_75t_L g1986 ( 
.A(n_1965),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1966),
.B(n_1965),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1968),
.A2(n_1939),
.B1(n_1949),
.B2(n_1952),
.C(n_1945),
.Y(n_1988)
);

OAI211xp5_ASAP7_75t_L g1989 ( 
.A1(n_1984),
.A2(n_1964),
.B(n_1941),
.C(n_1961),
.Y(n_1989)
);

AOI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1967),
.A2(n_1936),
.B1(n_1930),
.B2(n_1950),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1982),
.B(n_1983),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1967),
.A2(n_1930),
.B1(n_1915),
.B2(n_1933),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_SL g1993 ( 
.A(n_1986),
.B(n_1883),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1984),
.A2(n_1955),
.B1(n_1957),
.B2(n_1906),
.Y(n_1994)
);

AOI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1969),
.A2(n_1932),
.B1(n_1930),
.B2(n_1899),
.C(n_1929),
.Y(n_1995)
);

AOI211xp5_ASAP7_75t_SL g1996 ( 
.A1(n_1972),
.A2(n_1930),
.B(n_1929),
.C(n_1925),
.Y(n_1996)
);

OAI211xp5_ASAP7_75t_L g1997 ( 
.A1(n_1969),
.A2(n_1899),
.B(n_1925),
.C(n_1917),
.Y(n_1997)
);

NOR2xp67_ASAP7_75t_L g1998 ( 
.A(n_1976),
.B(n_1845),
.Y(n_1998)
);

AOI221xp5_ASAP7_75t_L g1999 ( 
.A1(n_1971),
.A2(n_1623),
.B1(n_1617),
.B2(n_1775),
.C(n_1660),
.Y(n_1999)
);

NOR2x1_ASAP7_75t_L g2000 ( 
.A(n_1989),
.B(n_1979),
.Y(n_2000)
);

OA22x2_ASAP7_75t_L g2001 ( 
.A1(n_1994),
.A2(n_1985),
.B1(n_1975),
.B2(n_1973),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1991),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1996),
.B(n_1973),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1997),
.B(n_1980),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1987),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1995),
.Y(n_2006)
);

AOI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1988),
.A2(n_1971),
.B1(n_1977),
.B2(n_1981),
.C(n_1970),
.Y(n_2007)
);

AND5x1_ASAP7_75t_L g2008 ( 
.A(n_1993),
.B(n_1999),
.C(n_1990),
.D(n_1992),
.E(n_1974),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1998),
.B(n_1978),
.Y(n_2009)
);

NOR3x1_ASAP7_75t_L g2010 ( 
.A(n_1989),
.B(n_1974),
.C(n_1851),
.Y(n_2010)
);

NOR3xp33_ASAP7_75t_L g2011 ( 
.A(n_1989),
.B(n_1794),
.C(n_1764),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1993),
.B(n_1764),
.Y(n_2012)
);

NOR3xp33_ASAP7_75t_L g2013 ( 
.A(n_2000),
.B(n_1794),
.C(n_1509),
.Y(n_2013)
);

OAI221xp5_ASAP7_75t_L g2014 ( 
.A1(n_2008),
.A2(n_1715),
.B1(n_1808),
.B2(n_1745),
.C(n_1638),
.Y(n_2014)
);

NOR3x1_ASAP7_75t_L g2015 ( 
.A(n_2004),
.B(n_1715),
.C(n_1800),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_2009),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2003),
.B(n_1808),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_2001),
.A2(n_1729),
.B(n_1772),
.Y(n_2018)
);

AOI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_2006),
.A2(n_1637),
.B1(n_1660),
.B2(n_1681),
.C(n_1669),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2016),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2017),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2015),
.Y(n_2022)
);

NAND3xp33_ASAP7_75t_SL g2023 ( 
.A(n_2013),
.B(n_2007),
.C(n_2006),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2018),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_2019),
.B(n_2002),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_2014),
.B(n_2005),
.Y(n_2026)
);

AOI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_2023),
.A2(n_2011),
.B1(n_2012),
.B2(n_2010),
.C(n_1660),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_2020),
.Y(n_2028)
);

NOR2x1p5_ASAP7_75t_L g2029 ( 
.A(n_2022),
.B(n_1808),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_2021),
.B(n_1797),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2024),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_2026),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2030),
.B(n_2025),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_2028),
.B(n_1772),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2030),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2032),
.B(n_1798),
.Y(n_2036)
);

XNOR2x1_ASAP7_75t_L g2037 ( 
.A(n_2033),
.B(n_2029),
.Y(n_2037)
);

XNOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2035),
.B(n_2031),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2038),
.Y(n_2039)
);

AOI21xp33_ASAP7_75t_SL g2040 ( 
.A1(n_2039),
.A2(n_2037),
.B(n_2036),
.Y(n_2040)
);

OAI22x1_ASAP7_75t_L g2041 ( 
.A1(n_2039),
.A2(n_2034),
.B1(n_2027),
.B2(n_1804),
.Y(n_2041)
);

NAND3xp33_ASAP7_75t_SL g2042 ( 
.A(n_2040),
.B(n_2034),
.C(n_1483),
.Y(n_2042)
);

OR2x6_ASAP7_75t_L g2043 ( 
.A(n_2041),
.B(n_1430),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_2043),
.B(n_1772),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2044),
.Y(n_2045)
);

AOI322xp5_ASAP7_75t_L g2046 ( 
.A1(n_2045),
.A2(n_2042),
.A3(n_1774),
.B1(n_1783),
.B2(n_1788),
.C1(n_1804),
.C2(n_1767),
.Y(n_2046)
);

OAI221xp5_ASAP7_75t_R g2047 ( 
.A1(n_2046),
.A2(n_1767),
.B1(n_1798),
.B2(n_1803),
.C(n_1806),
.Y(n_2047)
);

AOI211xp5_ASAP7_75t_L g2048 ( 
.A1(n_2047),
.A2(n_1483),
.B(n_1729),
.C(n_1462),
.Y(n_2048)
);


endmodule