module fake_jpeg_31813_n_382 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_8),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_52),
.Y(n_86)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_41),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_13),
.Y(n_52)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_12),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_60),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_36),
.B(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_17),
.Y(n_118)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_34),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_15),
.B1(n_26),
.B2(n_37),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_70),
.A2(n_85),
.B1(n_88),
.B2(n_91),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_23),
.B1(n_31),
.B2(n_22),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_72),
.A2(n_87),
.B1(n_110),
.B2(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_20),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_73),
.B(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_28),
.B1(n_29),
.B2(n_20),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_75),
.A2(n_90),
.B1(n_96),
.B2(n_100),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_44),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_82),
.B(n_94),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_23),
.B1(n_30),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_15),
.B1(n_31),
.B2(n_21),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_14),
.B1(n_30),
.B2(n_32),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_64),
.A2(n_34),
.B1(n_21),
.B2(n_29),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_20),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_16),
.B1(n_21),
.B2(n_34),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_39),
.B(n_30),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_98),
.B(n_5),
.C(n_7),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_51),
.A2(n_33),
.B1(n_32),
.B2(n_16),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_39),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_102),
.B(n_117),
.Y(n_148)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_59),
.A2(n_32),
.B1(n_33),
.B2(n_3),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_9),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_45),
.A2(n_33),
.B1(n_17),
.B2(n_3),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_41),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_110)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_53),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_113),
.B(n_78),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_49),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_49),
.B(n_2),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_17),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_121),
.B(n_131),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_122),
.B(n_155),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_61),
.B1(n_60),
.B2(n_67),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_140),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_69),
.A2(n_57),
.B1(n_103),
.B2(n_85),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

NOR4xp25_ASAP7_75t_SL g129 ( 
.A(n_116),
.B(n_86),
.C(n_91),
.D(n_87),
.Y(n_129)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_129),
.A2(n_138),
.B(n_94),
.Y(n_213)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_130),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_57),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_135),
.B(n_142),
.Y(n_210)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_83),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_145),
.B1(n_151),
.B2(n_154),
.Y(n_181)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_7),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g211 ( 
.A(n_143),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_72),
.A2(n_9),
.B1(n_88),
.B2(n_70),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_149),
.B(n_161),
.Y(n_172)
);

CKINVDCx12_ASAP7_75t_R g150 ( 
.A(n_112),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_150),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_9),
.B1(n_109),
.B2(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_81),
.A2(n_114),
.B1(n_71),
.B2(n_89),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_156),
.Y(n_185)
);

INVx6_ASAP7_75t_SL g157 ( 
.A(n_74),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_141),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_81),
.A2(n_114),
.B1(n_89),
.B2(n_97),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_125),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_84),
.A2(n_97),
.B1(n_105),
.B2(n_101),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_105),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_165),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_101),
.A2(n_104),
.B1(n_120),
.B2(n_99),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_132),
.B1(n_151),
.B2(n_157),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_56),
.B1(n_45),
.B2(n_44),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_82),
.B(n_75),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_166),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_83),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_82),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_169),
.B(n_170),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_82),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_145),
.B(n_131),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_194),
.B(n_209),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_179),
.B(n_196),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_170),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_180),
.B(n_187),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_186),
.A2(n_198),
.B1(n_185),
.B2(n_174),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_134),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_188),
.A2(n_208),
.B1(n_185),
.B2(n_195),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_121),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_201),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_132),
.A2(n_136),
.B(n_135),
.Y(n_194)
);

OA22x2_ASAP7_75t_SL g195 ( 
.A1(n_136),
.A2(n_168),
.B1(n_124),
.B2(n_161),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_147),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_147),
.A2(n_144),
.B1(n_166),
.B2(n_153),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_162),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_215),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_160),
.A2(n_123),
.B(n_171),
.C(n_144),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_203),
.B(n_214),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g208 ( 
.A1(n_146),
.A2(n_152),
.B1(n_143),
.B2(n_137),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_130),
.A2(n_126),
.B(n_145),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_213),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_133),
.B(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_170),
.B(n_169),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_233),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_188),
.B1(n_177),
.B2(n_202),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_219),
.A2(n_248),
.B1(n_189),
.B2(n_205),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_196),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_227),
.C(n_218),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_223),
.B(n_231),
.Y(n_275)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_176),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_202),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_178),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_228),
.B(n_234),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_207),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_172),
.B(n_199),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_197),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_238),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_179),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_181),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_237),
.B(n_241),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_212),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_240),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_191),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_191),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_242),
.A2(n_253),
.B1(n_252),
.B2(n_239),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_173),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_245),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_184),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_208),
.Y(n_249)
);

NAND2x1_ASAP7_75t_SL g270 ( 
.A(n_249),
.B(n_211),
.Y(n_270)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_216),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_174),
.A2(n_184),
.B1(n_182),
.B2(n_203),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_189),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_176),
.B(n_183),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_254),
.Y(n_269)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_175),
.B(n_201),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_257),
.A2(n_259),
.B(n_283),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_260),
.A2(n_261),
.B1(n_284),
.B2(n_236),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_219),
.A2(n_205),
.B1(n_175),
.B2(n_211),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_229),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_230),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_270),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_274),
.B(n_278),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_220),
.A2(n_211),
.B(n_241),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_276),
.A2(n_255),
.B(n_250),
.Y(n_300)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XNOR2x1_ASAP7_75t_L g278 ( 
.A(n_227),
.B(n_211),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_258),
.B1(n_259),
.B2(n_256),
.Y(n_287)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_244),
.B(n_242),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_232),
.A2(n_237),
.B1(n_226),
.B2(n_249),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_256),
.C(n_224),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_225),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_287),
.A2(n_298),
.B1(n_308),
.B2(n_261),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_217),
.C(n_230),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_290),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_289),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_294),
.B(n_301),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_233),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_296),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_256),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_297),
.A2(n_283),
.B1(n_282),
.B2(n_257),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_259),
.A2(n_247),
.B1(n_231),
.B2(n_223),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_277),
.Y(n_299)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_299),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_302),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_272),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_284),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_278),
.C(n_286),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_304),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_276),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_306),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_262),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_243),
.Y(n_307)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_262),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_281),
.Y(n_309)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_274),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_311),
.B(n_320),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_318),
.B1(n_298),
.B2(n_300),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_313),
.B(n_317),
.C(n_324),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_282),
.C(n_260),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_302),
.A2(n_270),
.B1(n_264),
.B2(n_285),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_264),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_287),
.B(n_295),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_269),
.C(n_267),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_326),
.A2(n_309),
.B(n_292),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_271),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_290),
.B(n_301),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_329),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_323),
.Y(n_335)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

A2O1A1O1Ixp25_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_299),
.B(n_291),
.C(n_307),
.D(n_304),
.Y(n_337)
);

NOR2x1_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_318),
.Y(n_356)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_338),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_325),
.A2(n_294),
.B(n_310),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_339),
.B(n_343),
.Y(n_350)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_322),
.A2(n_291),
.B(n_297),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_341),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_321),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_344),
.Y(n_354)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_347),
.B(n_348),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

AOI21x1_ASAP7_75t_SL g352 ( 
.A1(n_341),
.A2(n_328),
.B(n_330),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_359),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_356),
.A2(n_349),
.B1(n_352),
.B2(n_355),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_342),
.B(n_315),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_334),
.A2(n_312),
.B1(n_319),
.B2(n_326),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_360),
.A2(n_336),
.B1(n_317),
.B2(n_324),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_333),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_361),
.B(n_365),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_360),
.B(n_311),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_362),
.B(n_364),
.Y(n_372)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_363),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_346),
.C(n_345),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_357),
.A2(n_334),
.B1(n_308),
.B2(n_306),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_366),
.B(n_368),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_344),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_367),
.A2(n_358),
.B(n_353),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_370),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_371),
.B(n_364),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_376),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_368),
.Y(n_376)
);

AOI21xp33_ASAP7_75t_L g377 ( 
.A1(n_374),
.A2(n_372),
.B(n_369),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_377),
.B(n_376),
.C(n_368),
.Y(n_379)
);

OAI21x1_ASAP7_75t_L g380 ( 
.A1(n_379),
.A2(n_378),
.B(n_362),
.Y(n_380)
);

OAI21xp33_ASAP7_75t_L g381 ( 
.A1(n_380),
.A2(n_351),
.B(n_358),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_337),
.Y(n_382)
);


endmodule