module real_aes_17850_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_360;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_578;
wire n_892;
wire n_372;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_1584;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g928 ( .A(n_0), .Y(n_928) );
AOI221x1_ASAP7_75t_SL g941 ( .A1(n_0), .A2(n_2), .B1(n_320), .B2(n_942), .C(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g860 ( .A(n_1), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_2), .A2(n_22), .B1(n_665), .B2(n_685), .Y(n_936) );
INVx1_ASAP7_75t_L g1043 ( .A(n_3), .Y(n_1043) );
INVx1_ASAP7_75t_L g1555 ( .A(n_4), .Y(n_1555) );
INVx1_ASAP7_75t_L g719 ( .A(n_5), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g759 ( .A1(n_5), .A2(n_760), .B(n_761), .C(n_768), .Y(n_759) );
XNOR2xp5_ASAP7_75t_L g313 ( .A(n_6), .B(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g680 ( .A(n_7), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_7), .A2(n_116), .B1(n_709), .B2(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g513 ( .A(n_8), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_8), .A2(n_133), .B1(n_606), .B2(n_610), .Y(n_605) );
INVx1_ASAP7_75t_L g965 ( .A(n_9), .Y(n_965) );
OAI211xp5_ASAP7_75t_L g1013 ( .A1(n_9), .A2(n_342), .B(n_422), .C(n_1014), .Y(n_1013) );
AOI21xp33_ASAP7_75t_L g935 ( .A1(n_10), .A2(n_682), .B(n_683), .Y(n_935) );
INVx1_ASAP7_75t_L g953 ( .A(n_10), .Y(n_953) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_11), .A2(n_250), .B1(n_709), .B2(n_1038), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_11), .A2(n_136), .B1(n_497), .B2(n_502), .C(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1123 ( .A(n_12), .Y(n_1123) );
INVx1_ASAP7_75t_L g297 ( .A(n_13), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_13), .B(n_307), .Y(n_385) );
AND2x2_ASAP7_75t_L g494 ( .A(n_13), .B(n_453), .Y(n_494) );
AND2x2_ASAP7_75t_L g511 ( .A(n_13), .B(n_243), .Y(n_511) );
INVx1_ASAP7_75t_L g1200 ( .A(n_14), .Y(n_1200) );
OAI221xp5_ASAP7_75t_L g520 ( .A1(n_15), .A2(n_266), .B1(n_521), .B2(n_525), .C(n_530), .Y(n_520) );
INVx1_ASAP7_75t_L g595 ( .A(n_15), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g1217 ( .A1(n_16), .A2(n_113), .B1(n_502), .B2(n_659), .C(n_661), .Y(n_1217) );
INVx1_ASAP7_75t_L g1241 ( .A(n_16), .Y(n_1241) );
INVx1_ASAP7_75t_L g1135 ( .A(n_17), .Y(n_1135) );
INVx1_ASAP7_75t_L g432 ( .A(n_18), .Y(n_432) );
INVx1_ASAP7_75t_L g336 ( .A(n_19), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_20), .A2(n_279), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
OAI211xp5_ASAP7_75t_L g1048 ( .A1(n_20), .A2(n_1049), .B(n_1050), .C(n_1054), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_21), .B(n_1273), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_21), .B(n_111), .Y(n_1275) );
INVx2_ASAP7_75t_L g1279 ( .A(n_21), .Y(n_1279) );
AOI221xp5_ASAP7_75t_L g948 ( .A1(n_22), .A2(n_195), .B1(n_942), .B2(n_949), .C(n_951), .Y(n_948) );
INVx1_ASAP7_75t_L g825 ( .A(n_23), .Y(n_825) );
INVx1_ASAP7_75t_L g1557 ( .A(n_24), .Y(n_1557) );
INVx1_ASAP7_75t_L g1172 ( .A(n_25), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g1290 ( .A1(n_26), .A2(n_188), .B1(n_1274), .B2(n_1280), .Y(n_1290) );
INVx1_ASAP7_75t_L g1040 ( .A(n_27), .Y(n_1040) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_27), .A2(n_177), .B1(n_1060), .B2(n_1061), .C(n_1062), .Y(n_1059) );
INVx1_ASAP7_75t_L g831 ( .A(n_28), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g418 ( .A1(n_29), .A2(n_419), .B(n_422), .C(n_426), .Y(n_418) );
INVx1_ASAP7_75t_L g475 ( .A(n_29), .Y(n_475) );
INVx1_ASAP7_75t_L g1176 ( .A(n_30), .Y(n_1176) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_31), .A2(n_80), .B1(n_664), .B2(n_665), .Y(n_1218) );
INVx1_ASAP7_75t_L g1247 ( .A(n_31), .Y(n_1247) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_32), .A2(n_224), .B1(n_1270), .B2(n_1277), .Y(n_1324) );
INVx1_ASAP7_75t_L g627 ( .A(n_33), .Y(n_627) );
INVx1_ASAP7_75t_L g988 ( .A(n_34), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_35), .A2(n_108), .B1(n_581), .B2(n_707), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_35), .A2(n_251), .B1(n_921), .B2(n_1058), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_36), .A2(n_246), .B1(n_749), .B2(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g762 ( .A(n_36), .Y(n_762) );
INVx1_ASAP7_75t_L g964 ( .A(n_37), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_38), .A2(n_239), .B1(n_686), .B2(n_1224), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1248 ( .A1(n_38), .A2(n_113), .B1(n_699), .B2(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1171 ( .A(n_39), .Y(n_1171) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_40), .A2(n_229), .B1(n_1270), .B2(n_1280), .Y(n_1297) );
AOI22xp5_ASAP7_75t_L g1313 ( .A1(n_41), .A2(n_117), .B1(n_1270), .B2(n_1277), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g966 ( .A1(n_42), .A2(n_179), .B1(n_967), .B2(n_968), .Y(n_966) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_42), .A2(n_179), .B1(n_1010), .B2(n_1012), .Y(n_1009) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_43), .A2(n_149), .B1(n_497), .B2(n_498), .C(n_502), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_43), .A2(n_87), .B1(n_578), .B2(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g1100 ( .A(n_44), .Y(n_1100) );
AOI22xp33_ASAP7_75t_SL g740 ( .A1(n_45), .A2(n_123), .B1(n_741), .B2(n_742), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_45), .A2(n_246), .B1(n_492), .B2(n_767), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g1289 ( .A1(n_46), .A2(n_103), .B1(n_1270), .B2(n_1277), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_47), .A2(n_183), .B1(n_504), .B2(n_508), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_47), .A2(n_110), .B1(n_320), .B2(n_587), .Y(n_586) );
OAI211xp5_ASAP7_75t_L g883 ( .A1(n_48), .A2(n_803), .B(n_884), .C(n_886), .Y(n_883) );
INVx1_ASAP7_75t_L g894 ( .A(n_48), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_49), .A2(n_269), .B1(n_414), .B2(n_809), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_49), .A2(n_135), .B1(n_477), .B2(n_897), .Y(n_896) );
OAI22xp5_ASAP7_75t_SL g916 ( .A1(n_50), .A2(n_196), .B1(n_549), .B2(n_562), .Y(n_916) );
INVx1_ASAP7_75t_L g920 ( .A(n_50), .Y(n_920) );
INVx1_ASAP7_75t_L g1151 ( .A(n_51), .Y(n_1151) );
INVx1_ASAP7_75t_L g325 ( .A(n_52), .Y(n_325) );
INVx1_ASAP7_75t_L g334 ( .A(n_52), .Y(n_334) );
INVx1_ASAP7_75t_L g747 ( .A(n_53), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_53), .A2(n_252), .B1(n_492), .B2(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_54), .A2(n_625), .B1(n_712), .B2(n_713), .Y(n_624) );
INVxp67_ASAP7_75t_L g713 ( .A(n_54), .Y(n_713) );
INVx1_ASAP7_75t_L g1074 ( .A(n_55), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1496 ( .A1(n_56), .A2(n_82), .B1(n_742), .B2(n_1497), .Y(n_1496) );
AOI221xp5_ASAP7_75t_L g1502 ( .A1(n_56), .A2(n_265), .B1(n_497), .B2(n_502), .C(n_765), .Y(n_1502) );
INVx1_ASAP7_75t_L g436 ( .A(n_57), .Y(n_436) );
OAI211xp5_ASAP7_75t_L g456 ( .A1(n_57), .A2(n_457), .B(n_461), .C(n_466), .Y(n_456) );
INVx1_ASAP7_75t_L g1559 ( .A(n_58), .Y(n_1559) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_59), .Y(n_652) );
INVx1_ASAP7_75t_L g1230 ( .A(n_60), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_61), .A2(n_715), .B1(n_716), .B2(n_775), .Y(n_714) );
INVxp67_ASAP7_75t_L g775 ( .A(n_61), .Y(n_775) );
INVx1_ASAP7_75t_L g290 ( .A(n_62), .Y(n_290) );
INVx1_ASAP7_75t_L g866 ( .A(n_63), .Y(n_866) );
INVx2_ASAP7_75t_L g356 ( .A(n_64), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_65), .A2(n_89), .B1(n_1277), .B2(n_1284), .Y(n_1298) );
OAI22xp33_ASAP7_75t_L g1202 ( .A1(n_66), .A2(n_167), .B1(n_809), .B2(n_882), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1209 ( .A1(n_66), .A2(n_167), .B1(n_970), .B2(n_1157), .Y(n_1209) );
INVx1_ASAP7_75t_L g838 ( .A(n_67), .Y(n_838) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_68), .A2(n_237), .B1(n_559), .B2(n_564), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_69), .A2(n_276), .B1(n_685), .B2(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g697 ( .A(n_69), .Y(n_697) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_70), .A2(n_74), .B1(n_299), .B2(n_795), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_70), .A2(n_74), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
INVx1_ASAP7_75t_L g557 ( .A(n_71), .Y(n_557) );
INVx1_ASAP7_75t_L g862 ( .A(n_72), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g1495 ( .A1(n_73), .A2(n_160), .B1(n_707), .B2(n_1494), .Y(n_1495) );
AOI22xp33_ASAP7_75t_L g1503 ( .A1(n_73), .A2(n_158), .B1(n_1504), .B2(n_1505), .Y(n_1503) );
INVx1_ASAP7_75t_L g1122 ( .A(n_75), .Y(n_1122) );
OAI22xp5_ASAP7_75t_L g1194 ( .A1(n_76), .A2(n_141), .B1(n_808), .B2(n_1195), .Y(n_1194) );
OAI22xp33_ASAP7_75t_L g1204 ( .A1(n_76), .A2(n_141), .B1(n_968), .B2(n_1205), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_77), .A2(n_112), .B1(n_661), .B2(n_930), .C(n_1222), .Y(n_1221) );
INVxp67_ASAP7_75t_SL g1234 ( .A(n_77), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_78), .A2(n_272), .B1(n_790), .B2(n_792), .Y(n_789) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_78), .A2(n_107), .B1(n_798), .B2(n_799), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g1294 ( .A1(n_79), .A2(n_140), .B1(n_1270), .B2(n_1277), .Y(n_1294) );
INVxp67_ASAP7_75t_SL g1235 ( .A(n_80), .Y(n_1235) );
OAI211xp5_ASAP7_75t_L g961 ( .A1(n_81), .A2(n_864), .B(n_962), .C(n_963), .Y(n_961) );
INVx1_ASAP7_75t_L g1016 ( .A(n_81), .Y(n_1016) );
INVx1_ASAP7_75t_L g1526 ( .A(n_82), .Y(n_1526) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_83), .Y(n_720) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_83), .A2(n_231), .B1(n_526), .B2(n_556), .C(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_84), .A2(n_116), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_84), .A2(n_211), .B1(n_699), .B2(n_702), .Y(n_698) );
INVx1_ASAP7_75t_L g1125 ( .A(n_85), .Y(n_1125) );
OAI211xp5_ASAP7_75t_L g1573 ( .A1(n_86), .A2(n_892), .B(n_962), .C(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1583 ( .A(n_86), .Y(n_1583) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_87), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_88), .A2(n_95), .B1(n_798), .B2(n_882), .Y(n_1148) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_88), .A2(n_119), .B1(n_299), .B2(n_450), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1577 ( .A1(n_90), .A2(n_199), .B1(n_477), .B2(n_1105), .Y(n_1577) );
OAI22xp33_ASAP7_75t_L g1584 ( .A1(n_90), .A2(n_199), .B1(n_438), .B2(n_440), .Y(n_1584) );
INVx1_ASAP7_75t_L g1073 ( .A(n_91), .Y(n_1073) );
INVx1_ASAP7_75t_L g1490 ( .A(n_92), .Y(n_1490) );
OAI211xp5_ASAP7_75t_L g1500 ( .A1(n_92), .A2(n_490), .B(n_1501), .C(n_1507), .Y(n_1500) );
OAI221xp5_ASAP7_75t_SL g646 ( .A1(n_93), .A2(n_96), .B1(n_647), .B2(n_649), .C(n_651), .Y(n_646) );
INVx1_ASAP7_75t_L g673 ( .A(n_93), .Y(n_673) );
INVx1_ASAP7_75t_L g933 ( .A(n_94), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_95), .A2(n_194), .B1(n_790), .B2(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g689 ( .A(n_96), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g725 ( .A(n_97), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g1302 ( .A1(n_98), .A2(n_137), .B1(n_1270), .B2(n_1277), .Y(n_1302) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_99), .B(n_778), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_100), .A2(n_958), .B1(n_959), .B2(n_1019), .Y(n_957) );
INVxp67_ASAP7_75t_SL g1019 ( .A(n_100), .Y(n_1019) );
AOI22xp5_ASAP7_75t_SL g1301 ( .A1(n_100), .A2(n_271), .B1(n_1280), .B2(n_1284), .Y(n_1301) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_101), .Y(n_1532) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_102), .Y(n_292) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_102), .B(n_290), .Y(n_1271) );
INVx1_ASAP7_75t_L g1260 ( .A(n_104), .Y(n_1260) );
INVx1_ASAP7_75t_L g1078 ( .A(n_105), .Y(n_1078) );
INVx1_ASAP7_75t_L g1136 ( .A(n_106), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_107), .A2(n_189), .B1(n_299), .B2(n_795), .Y(n_794) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_108), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g1312 ( .A1(n_109), .A2(n_121), .B1(n_1274), .B2(n_1280), .Y(n_1312) );
AOI221xp5_ASAP7_75t_L g536 ( .A1(n_110), .A2(n_176), .B1(n_500), .B2(n_537), .C(n_539), .Y(n_536) );
INVx1_ASAP7_75t_L g1273 ( .A(n_111), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_111), .B(n_1279), .Y(n_1281) );
INVx1_ASAP7_75t_L g1245 ( .A(n_112), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_114), .A2(n_275), .B1(n_1270), .B2(n_1274), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_115), .A2(n_251), .B1(n_581), .B2(n_1035), .Y(n_1034) );
AOI21xp33_ASAP7_75t_L g1064 ( .A1(n_115), .A2(n_539), .B(n_765), .Y(n_1064) );
XOR2xp5_ASAP7_75t_L g1542 ( .A(n_118), .B(n_1543), .Y(n_1542) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_119), .A2(n_194), .B1(n_808), .B2(n_809), .Y(n_1153) );
INVx1_ASAP7_75t_L g636 ( .A(n_120), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_122), .A2(n_265), .B1(n_742), .B2(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1517 ( .A(n_122), .Y(n_1517) );
AOI21xp33_ASAP7_75t_L g764 ( .A1(n_123), .A2(n_683), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g1082 ( .A(n_124), .Y(n_1082) );
INVx2_ASAP7_75t_L g355 ( .A(n_125), .Y(n_355) );
INVx1_ASAP7_75t_L g367 ( .A(n_125), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_125), .B(n_356), .Y(n_553) );
XNOR2xp5_ASAP7_75t_L g853 ( .A(n_126), .B(n_854), .Y(n_853) );
AOI22xp5_ASAP7_75t_L g1285 ( .A1(n_127), .A2(n_249), .B1(n_1270), .B2(n_1277), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1510 ( .A(n_128), .Y(n_1510) );
INVx1_ASAP7_75t_L g975 ( .A(n_129), .Y(n_975) );
INVx1_ASAP7_75t_L g341 ( .A(n_130), .Y(n_341) );
INVx1_ASAP7_75t_L g1178 ( .A(n_131), .Y(n_1178) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_132), .A2(n_219), .B1(n_610), .B2(n_635), .Y(n_1030) );
INVx1_ASAP7_75t_L g1052 ( .A(n_132), .Y(n_1052) );
INVx1_ASAP7_75t_L g516 ( .A(n_133), .Y(n_516) );
INVx1_ASAP7_75t_L g1575 ( .A(n_134), .Y(n_1575) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_135), .A2(n_198), .B1(n_798), .B2(n_882), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_136), .A2(n_201), .B1(n_579), .B2(n_749), .Y(n_1033) );
INVx1_ASAP7_75t_L g833 ( .A(n_138), .Y(n_833) );
INVx1_ASAP7_75t_L g1201 ( .A(n_139), .Y(n_1201) );
OAI211xp5_ASAP7_75t_L g1206 ( .A1(n_139), .A2(n_783), .B(n_864), .C(n_1207), .Y(n_1206) );
NOR2xp33_ASAP7_75t_L g1227 ( .A(n_142), .B(n_526), .Y(n_1227) );
INVxp67_ASAP7_75t_SL g1254 ( .A(n_142), .Y(n_1254) );
INVx1_ASAP7_75t_L g788 ( .A(n_143), .Y(n_788) );
OAI211xp5_ASAP7_75t_L g800 ( .A1(n_143), .A2(n_801), .B(n_803), .C(n_804), .Y(n_800) );
INVx1_ASAP7_75t_L g887 ( .A(n_144), .Y(n_887) );
XNOR2xp5_ASAP7_75t_L g1027 ( .A(n_145), .B(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1550 ( .A(n_146), .Y(n_1550) );
INVx1_ASAP7_75t_L g318 ( .A(n_147), .Y(n_318) );
INVx1_ASAP7_75t_L g730 ( .A(n_148), .Y(n_730) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_148), .A2(n_184), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_149), .A2(n_190), .B1(n_576), .B2(n_579), .Y(n_575) );
INVx1_ASAP7_75t_L g984 ( .A(n_150), .Y(n_984) );
OAI211xp5_ASAP7_75t_L g780 ( .A1(n_151), .A2(n_781), .B(n_783), .C(n_784), .Y(n_780) );
INVx1_ASAP7_75t_L g806 ( .A(n_151), .Y(n_806) );
INVx1_ASAP7_75t_L g905 ( .A(n_152), .Y(n_905) );
INVx1_ASAP7_75t_L g1551 ( .A(n_153), .Y(n_1551) );
INVx1_ASAP7_75t_L g370 ( .A(n_154), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_155), .A2(n_178), .B1(n_438), .B2(n_440), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_155), .A2(n_178), .B1(n_477), .B2(n_479), .Y(n_476) );
OAI211xp5_ASAP7_75t_L g1098 ( .A1(n_156), .A2(n_892), .B(n_962), .C(n_1099), .Y(n_1098) );
INVx1_ASAP7_75t_L g1112 ( .A(n_156), .Y(n_1112) );
INVx1_ASAP7_75t_L g841 ( .A(n_157), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g1492 ( .A1(n_158), .A2(n_162), .B1(n_707), .B2(n_709), .Y(n_1492) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_159), .Y(n_745) );
INVx1_ASAP7_75t_L g1515 ( .A(n_160), .Y(n_1515) );
INVx1_ASAP7_75t_L g1226 ( .A(n_161), .Y(n_1226) );
INVx1_ASAP7_75t_L g1521 ( .A(n_162), .Y(n_1521) );
INVx1_ASAP7_75t_L g736 ( .A(n_163), .Y(n_736) );
AOI21xp33_ASAP7_75t_L g769 ( .A1(n_163), .A2(n_500), .B(n_539), .Y(n_769) );
INVx1_ASAP7_75t_L g869 ( .A(n_164), .Y(n_869) );
INVx1_ASAP7_75t_L g1131 ( .A(n_165), .Y(n_1131) );
INVx1_ASAP7_75t_L g1181 ( .A(n_166), .Y(n_1181) );
AOI22xp5_ASAP7_75t_L g1292 ( .A1(n_168), .A2(n_261), .B1(n_1280), .B2(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1229 ( .A(n_169), .Y(n_1229) );
OAI322xp33_ASAP7_75t_L g1232 ( .A1(n_169), .A2(n_348), .A3(n_638), .B1(n_753), .B2(n_1233), .C1(n_1236), .C2(n_1242), .Y(n_1232) );
OAI22xp33_ASAP7_75t_L g1572 ( .A1(n_170), .A2(n_255), .B1(n_299), .B2(n_795), .Y(n_1572) );
OAI22xp5_ASAP7_75t_L g1579 ( .A1(n_170), .A2(n_255), .B1(n_1108), .B2(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g863 ( .A(n_171), .Y(n_863) );
BUFx3_ASAP7_75t_L g327 ( .A(n_172), .Y(n_327) );
INVx1_ASAP7_75t_L g987 ( .A(n_173), .Y(n_987) );
INVx1_ASAP7_75t_L g870 ( .A(n_174), .Y(n_870) );
INVx1_ASAP7_75t_L g1214 ( .A(n_175), .Y(n_1214) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_176), .A2(n_183), .B1(n_581), .B2(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g1041 ( .A(n_177), .Y(n_1041) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_180), .Y(n_304) );
INVx1_ASAP7_75t_L g630 ( .A(n_181), .Y(n_630) );
INVx1_ASAP7_75t_L g823 ( .A(n_182), .Y(n_823) );
INVx1_ASAP7_75t_L g728 ( .A(n_184), .Y(n_728) );
INVx1_ASAP7_75t_L g1086 ( .A(n_185), .Y(n_1086) );
INVx1_ASAP7_75t_L g372 ( .A(n_186), .Y(n_372) );
INVx1_ASAP7_75t_L g358 ( .A(n_187), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_189), .A2(n_272), .B1(n_808), .B2(n_809), .Y(n_807) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_190), .Y(n_533) );
INVx1_ASAP7_75t_L g888 ( .A(n_191), .Y(n_888) );
OAI211xp5_ASAP7_75t_SL g891 ( .A1(n_191), .A2(n_783), .B(n_892), .C(n_893), .Y(n_891) );
INVx1_ASAP7_75t_L g1080 ( .A(n_192), .Y(n_1080) );
OAI211xp5_ASAP7_75t_L g1149 ( .A1(n_193), .A2(n_801), .B(n_803), .C(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1161 ( .A(n_193), .Y(n_1161) );
AOI21xp33_ASAP7_75t_L g929 ( .A1(n_195), .A2(n_662), .B(n_930), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_196), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1251 ( .A(n_197), .Y(n_1251) );
OAI22xp33_ASAP7_75t_L g899 ( .A1(n_198), .A2(n_269), .B1(n_299), .B2(n_450), .Y(n_899) );
XOR2x2_ASAP7_75t_L g486 ( .A(n_200), .B(n_487), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_201), .A2(n_250), .B1(n_686), .B2(n_921), .Y(n_1065) );
INVx1_ASAP7_75t_L g1077 ( .A(n_202), .Y(n_1077) );
INVx1_ASAP7_75t_L g1103 ( .A(n_203), .Y(n_1103) );
OAI211xp5_ASAP7_75t_SL g1110 ( .A1(n_203), .A2(n_803), .B(n_946), .C(n_1111), .Y(n_1110) );
OAI222xp33_ASAP7_75t_L g907 ( .A1(n_204), .A2(n_244), .B1(n_254), .B2(n_564), .C1(n_908), .C2(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g1219 ( .A(n_205), .Y(n_1219) );
XOR2xp5_ASAP7_75t_L g1166 ( .A(n_206), .B(n_1167), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_206), .A2(n_212), .B1(n_1274), .B2(n_1280), .Y(n_1323) );
AOI22xp5_ASAP7_75t_L g1283 ( .A1(n_207), .A2(n_278), .B1(n_1280), .B2(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1533 ( .A(n_207), .Y(n_1533) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_207), .A2(n_1538), .B1(n_1541), .B2(n_1585), .Y(n_1537) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_208), .A2(n_277), .B1(n_665), .B2(n_685), .Y(n_931) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_208), .Y(n_952) );
INVx1_ASAP7_75t_L g1174 ( .A(n_209), .Y(n_1174) );
INVx1_ASAP7_75t_L g1487 ( .A(n_210), .Y(n_1487) );
OAI222xp33_ASAP7_75t_L g1513 ( .A1(n_210), .A2(n_274), .B1(n_525), .B2(n_938), .C1(n_1514), .C2(n_1520), .Y(n_1513) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_211), .A2(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g1129 ( .A(n_213), .Y(n_1129) );
INVx1_ASAP7_75t_L g983 ( .A(n_214), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_215), .Y(n_1512) );
INVx1_ASAP7_75t_L g1576 ( .A(n_216), .Y(n_1576) );
OAI211xp5_ASAP7_75t_L g1581 ( .A1(n_216), .A2(n_422), .B(n_946), .C(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g360 ( .A(n_217), .Y(n_360) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
INVx1_ASAP7_75t_L g1051 ( .A(n_219), .Y(n_1051) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_220), .A2(n_236), .B1(n_411), .B2(n_414), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g449 ( .A1(n_220), .A2(n_236), .B1(n_299), .B2(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g978 ( .A(n_221), .Y(n_978) );
INVx1_ASAP7_75t_L g994 ( .A(n_222), .Y(n_994) );
INVx1_ASAP7_75t_L g1085 ( .A(n_223), .Y(n_1085) );
INVx1_ASAP7_75t_L g1562 ( .A(n_225), .Y(n_1562) );
INVx1_ASAP7_75t_L g867 ( .A(n_226), .Y(n_867) );
INVx1_ASAP7_75t_L g724 ( .A(n_227), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_228), .A2(n_238), .B1(n_659), .B2(n_661), .C(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g696 ( .A(n_228), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g969 ( .A1(n_230), .A2(n_245), .B1(n_970), .B2(n_971), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g1017 ( .A1(n_230), .A2(n_245), .B1(n_809), .B2(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g723 ( .A(n_231), .Y(n_723) );
INVx1_ASAP7_75t_L g1132 ( .A(n_232), .Y(n_1132) );
CKINVDCx5p33_ASAP7_75t_R g914 ( .A(n_233), .Y(n_914) );
INVx1_ASAP7_75t_L g328 ( .A(n_234), .Y(n_328) );
INVx1_ASAP7_75t_L g814 ( .A(n_235), .Y(n_814) );
OAI211xp5_ASAP7_75t_L g489 ( .A1(n_237), .A2(n_490), .B(n_495), .C(n_512), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_238), .A2(n_276), .B1(n_706), .B2(n_707), .Y(n_705) );
INVxp67_ASAP7_75t_SL g1237 ( .A(n_239), .Y(n_1237) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_240), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_241), .A2(n_256), .B1(n_477), .B2(n_1105), .Y(n_1104) );
OAI22xp33_ASAP7_75t_L g1113 ( .A1(n_241), .A2(n_256), .B1(n_438), .B2(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1554 ( .A(n_242), .Y(n_1554) );
BUFx3_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
INVx1_ASAP7_75t_L g453 ( .A(n_243), .Y(n_453) );
INVx1_ASAP7_75t_L g1152 ( .A(n_247), .Y(n_1152) );
OAI211xp5_ASAP7_75t_L g1159 ( .A1(n_247), .A2(n_892), .B(n_962), .C(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g993 ( .A(n_248), .Y(n_993) );
INVx1_ASAP7_75t_L g739 ( .A(n_252), .Y(n_739) );
INVx1_ASAP7_75t_L g353 ( .A(n_253), .Y(n_353) );
INVx1_ASAP7_75t_L g366 ( .A(n_253), .Y(n_366) );
INVx2_ASAP7_75t_L g384 ( .A(n_253), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_254), .A2(n_259), .B1(n_758), .B2(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g1183 ( .A(n_257), .Y(n_1183) );
OAI211xp5_ASAP7_75t_L g1197 ( .A1(n_258), .A2(n_803), .B(n_1198), .C(n_1199), .Y(n_1197) );
INVx1_ASAP7_75t_L g1208 ( .A(n_258), .Y(n_1208) );
INVx1_ASAP7_75t_L g915 ( .A(n_259), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1276 ( .A1(n_260), .A2(n_262), .B1(n_1277), .B2(n_1280), .Y(n_1276) );
INVx1_ASAP7_75t_L g818 ( .A(n_263), .Y(n_818) );
INVx1_ASAP7_75t_L g1179 ( .A(n_264), .Y(n_1179) );
INVx1_ASAP7_75t_L g600 ( .A(n_266), .Y(n_600) );
XNOR2xp5_ASAP7_75t_L g1068 ( .A(n_267), .B(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g785 ( .A(n_268), .Y(n_785) );
INVx1_ASAP7_75t_L g1561 ( .A(n_270), .Y(n_1561) );
INVx1_ASAP7_75t_L g859 ( .A(n_273), .Y(n_859) );
INVx1_ASAP7_75t_L g1486 ( .A(n_274), .Y(n_1486) );
XOR2x2_ASAP7_75t_L g1117 ( .A(n_275), .B(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g944 ( .A(n_277), .Y(n_944) );
OAI21xp33_ASAP7_75t_L g1528 ( .A1(n_280), .A2(n_1529), .B(n_1530), .Y(n_1528) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_308), .B(n_1264), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx4f_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_293), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g1536 ( .A(n_287), .B(n_296), .Y(n_1536) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g1540 ( .A(n_289), .B(n_292), .Y(n_1540) );
INVx1_ASAP7_75t_L g1587 ( .A(n_289), .Y(n_1587) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g1589 ( .A(n_292), .B(n_1587), .Y(n_1589) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g483 ( .A(n_296), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x4_ASAP7_75t_L g406 ( .A(n_297), .B(n_307), .Y(n_406) );
AND2x4_ASAP7_75t_L g540 ( .A(n_297), .B(n_306), .Y(n_540) );
INVx1_ASAP7_75t_L g967 ( .A(n_298), .Y(n_967) );
INVx1_ASAP7_75t_L g1205 ( .A(n_298), .Y(n_1205) );
AND2x4_ASAP7_75t_SL g1535 ( .A(n_298), .B(n_1536), .Y(n_1535) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_300), .B(n_305), .Y(n_299) );
BUFx4f_ASAP7_75t_L g375 ( .A(n_300), .Y(n_375) );
OR2x6_ASAP7_75t_L g478 ( .A(n_300), .B(n_452), .Y(n_478) );
INVx1_ASAP7_75t_L g1146 ( .A(n_300), .Y(n_1146) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g401 ( .A(n_301), .Y(n_401) );
BUFx4f_ASAP7_75t_L g817 ( .A(n_301), .Y(n_817) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx2_ASAP7_75t_L g380 ( .A(n_303), .Y(n_380) );
INVx2_ASAP7_75t_L g391 ( .A(n_303), .Y(n_391) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_303), .B(n_304), .Y(n_395) );
AND2x2_ASAP7_75t_L g454 ( .A(n_303), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g465 ( .A(n_303), .B(n_304), .Y(n_465) );
INVx1_ASAP7_75t_L g474 ( .A(n_303), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_304), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g390 ( .A(n_304), .B(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g455 ( .A(n_304), .Y(n_455) );
BUFx2_ASAP7_75t_L g469 ( .A(n_304), .Y(n_469) );
AND2x2_ASAP7_75t_L g493 ( .A(n_304), .B(n_380), .Y(n_493) );
INVx1_ASAP7_75t_L g507 ( .A(n_304), .Y(n_507) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g463 ( .A(n_306), .Y(n_463) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g468 ( .A(n_307), .Y(n_468) );
AND2x4_ASAP7_75t_L g472 ( .A(n_307), .B(n_473), .Y(n_472) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_1021), .B1(n_1022), .B2(n_1262), .Y(n_308) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_620), .Y(n_309) );
XNOR2xp5_ASAP7_75t_L g1263 ( .A(n_310), .B(n_620), .Y(n_1263) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_486), .B1(n_618), .B2(n_619), .Y(n_310) );
INVx1_ASAP7_75t_L g618 ( .A(n_311), .Y(n_618) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_409), .C(n_448), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_373), .Y(n_315) );
OAI33xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_335), .A3(n_348), .B1(n_357), .B2(n_361), .B3(n_368), .Y(n_316) );
OAI22xp33_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_319), .B1(n_328), .B2(n_329), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_318), .A2(n_370), .B1(n_387), .B2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g876 ( .A(n_320), .Y(n_876) );
INVx8_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
INVx5_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_SL g874 ( .A(n_322), .Y(n_874) );
INVx3_ASAP7_75t_L g1128 ( .A(n_322), .Y(n_1128) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_323), .Y(n_417) );
BUFx8_ASAP7_75t_L g613 ( .A(n_323), .Y(n_613) );
INVx2_ASAP7_75t_L g641 ( .A(n_323), .Y(n_641) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVxp67_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g340 ( .A(n_325), .Y(n_340) );
AND2x4_ASAP7_75t_L g566 ( .A(n_326), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_327), .B(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g339 ( .A(n_327), .B(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_327), .Y(n_347) );
AND2x4_ASAP7_75t_L g424 ( .A(n_327), .B(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_328), .A2(n_372), .B1(n_400), .B2(n_402), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_329), .A2(n_695), .B1(n_696), .B2(n_697), .C(n_698), .Y(n_694) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g877 ( .A(n_331), .Y(n_877) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g371 ( .A(n_332), .Y(n_371) );
OR2x6_ASAP7_75t_L g442 ( .A(n_332), .B(n_364), .Y(n_442) );
BUFx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g551 ( .A(n_333), .Y(n_551) );
INVx1_ASAP7_75t_L g346 ( .A(n_334), .Y(n_346) );
INVx2_ASAP7_75t_L g425 ( .A(n_334), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B1(n_341), .B2(n_342), .Y(n_335) );
OAI22xp33_ASAP7_75t_L g374 ( .A1(n_336), .A2(n_358), .B1(n_375), .B2(n_376), .Y(n_374) );
BUFx4f_ASAP7_75t_SL g945 ( .A(n_337), .Y(n_945) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_SL g607 ( .A(n_338), .Y(n_607) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g359 ( .A(n_339), .Y(n_359) );
OR2x4_ASAP7_75t_L g413 ( .A(n_339), .B(n_364), .Y(n_413) );
OR2x4_ASAP7_75t_L g439 ( .A(n_339), .B(n_416), .Y(n_439) );
BUFx4f_ASAP7_75t_L g850 ( .A(n_339), .Y(n_850) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_339), .Y(n_1240) );
INVx1_ASAP7_75t_L g567 ( .A(n_340), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_341), .A2(n_360), .B1(n_397), .B2(n_398), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_342), .A2(n_358), .B1(n_359), .B2(n_360), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_342), .A2(n_607), .B1(n_814), .B2(n_831), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_342), .A2(n_976), .B1(n_993), .B2(n_994), .Y(n_992) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_344), .Y(n_851) );
HB1xp67_ASAP7_75t_L g1552 ( .A(n_344), .Y(n_1552) );
HB1xp67_ASAP7_75t_L g1563 ( .A(n_344), .Y(n_1563) );
BUFx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g421 ( .A(n_345), .Y(n_421) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_345), .Y(n_563) );
NAND2x1p5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
BUFx2_ASAP7_75t_L g435 ( .A(n_346), .Y(n_435) );
BUFx2_ASAP7_75t_L g431 ( .A(n_347), .Y(n_431) );
AND2x4_ASAP7_75t_L g584 ( .A(n_347), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g598 ( .A(n_347), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_348), .A2(n_734), .B1(n_743), .B2(n_753), .Y(n_733) );
OAI33xp33_ASAP7_75t_L g973 ( .A1(n_348), .A2(n_974), .A3(n_982), .B1(n_986), .B2(n_989), .B3(n_992), .Y(n_973) );
OAI33xp33_ASAP7_75t_L g1120 ( .A1(n_348), .A2(n_753), .A3(n_1121), .B1(n_1124), .B2(n_1130), .B3(n_1133), .Y(n_1120) );
OAI33xp33_ASAP7_75t_L g1169 ( .A1(n_348), .A2(n_989), .A3(n_1170), .B1(n_1173), .B2(n_1177), .B3(n_1180), .Y(n_1169) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx4f_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx4f_ASAP7_75t_L g703 ( .A(n_350), .Y(n_703) );
BUFx8_ASAP7_75t_L g1548 ( .A(n_350), .Y(n_1548) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g408 ( .A(n_351), .Y(n_408) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_351), .Y(n_447) );
OR2x2_ASAP7_75t_L g552 ( .A(n_351), .B(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g485 ( .A(n_352), .Y(n_485) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp33_ASAP7_75t_SL g354 ( .A(n_355), .B(n_356), .Y(n_354) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_355), .Y(n_445) );
INVx1_ASAP7_75t_L g569 ( .A(n_355), .Y(n_569) );
AND3x4_ASAP7_75t_L g574 ( .A(n_355), .B(n_430), .C(n_545), .Y(n_574) );
INVx3_ASAP7_75t_L g364 ( .A(n_356), .Y(n_364) );
BUFx3_ASAP7_75t_L g430 ( .A(n_356), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g1072 ( .A1(n_359), .A2(n_1073), .B1(n_1074), .B2(n_1075), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1549 ( .A1(n_359), .A2(n_1550), .B1(n_1551), .B2(n_1552), .Y(n_1549) );
OAI22xp33_ASAP7_75t_L g1560 ( .A1(n_359), .A2(n_1561), .B1(n_1562), .B2(n_1563), .Y(n_1560) );
OAI33xp33_ASAP7_75t_L g1071 ( .A1(n_361), .A2(n_703), .A3(n_1072), .B1(n_1076), .B2(n_1079), .B3(n_1084), .Y(n_1071) );
OAI33xp33_ASAP7_75t_L g1547 ( .A1(n_361), .A2(n_1548), .A3(n_1549), .B1(n_1553), .B2(n_1556), .B3(n_1560), .Y(n_1547) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_362), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_362), .B(n_705), .C(n_708), .Y(n_704) );
INVx2_ASAP7_75t_L g753 ( .A(n_362), .Y(n_753) );
INVx2_ASAP7_75t_L g878 ( .A(n_362), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g940 ( .A1(n_362), .A2(n_616), .B1(n_941), .B2(n_948), .C(n_955), .Y(n_940) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g991 ( .A(n_363), .Y(n_991) );
NAND3x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .C(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g416 ( .A(n_364), .Y(n_416) );
AND2x4_ASAP7_75t_L g423 ( .A(n_364), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g568 ( .A(n_364), .B(n_569), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_364), .B(n_367), .Y(n_590) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g555 ( .A(n_366), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_370), .B1(n_371), .B2(n_372), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g1233 ( .A1(n_369), .A2(n_737), .B1(n_1234), .B2(n_1235), .Y(n_1233) );
INVx1_ASAP7_75t_L g1494 ( .A(n_369), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1553 ( .A1(n_369), .A2(n_737), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_371), .A2(n_823), .B1(n_838), .B2(n_845), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_371), .A2(n_862), .B1(n_869), .B2(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g1556 ( .A1(n_371), .A2(n_1557), .B1(n_1558), .B2(n_1559), .Y(n_1556) );
OAI33xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_381), .A3(n_386), .B1(n_396), .B2(n_399), .B3(n_404), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_376), .A2(n_1550), .B1(n_1561), .B2(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_377), .Y(n_403) );
INVx2_ASAP7_75t_SL g821 ( .A(n_377), .Y(n_821) );
INVx1_ASAP7_75t_L g840 ( .A(n_377), .Y(n_840) );
INVx4_ASAP7_75t_L g1002 ( .A(n_377), .Y(n_1002) );
INVx2_ASAP7_75t_L g1525 ( .A(n_377), .Y(n_1525) );
INVx8_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g481 ( .A(n_378), .B(n_468), .Y(n_481) );
BUFx2_ASAP7_75t_L g534 ( .A(n_378), .Y(n_534) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI33xp33_ASAP7_75t_L g812 ( .A1(n_381), .A2(n_813), .A3(n_822), .B1(n_827), .B2(n_834), .B3(n_837), .Y(n_812) );
OAI33xp33_ASAP7_75t_L g995 ( .A1(n_381), .A2(n_834), .A3(n_996), .B1(n_1003), .B2(n_1006), .B3(n_1007), .Y(n_995) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx4_ASAP7_75t_L g857 ( .A(n_382), .Y(n_857) );
INVx2_ASAP7_75t_L g1089 ( .A(n_382), .Y(n_1089) );
INVx2_ASAP7_75t_L g1138 ( .A(n_382), .Y(n_1138) );
AND2x4_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
OR2x6_ASAP7_75t_L g589 ( .A(n_383), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g692 ( .A(n_383), .Y(n_692) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g545 ( .A(n_384), .Y(n_545) );
INVx4_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g397 ( .A(n_388), .Y(n_397) );
INVx2_ASAP7_75t_L g824 ( .A(n_388), .Y(n_824) );
INVx2_ASAP7_75t_L g1516 ( .A(n_388), .Y(n_1516) );
INVx4_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g830 ( .A(n_390), .Y(n_830) );
INVx2_ASAP7_75t_L g1005 ( .A(n_390), .Y(n_1005) );
AND2x2_ASAP7_75t_L g506 ( .A(n_391), .B(n_507), .Y(n_506) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_391), .Y(n_671) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_392), .A2(n_680), .B(n_681), .C(n_684), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_392), .A2(n_828), .B1(n_866), .B2(n_867), .Y(n_865) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_392), .A2(n_1077), .B1(n_1080), .B2(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1567 ( .A1(n_392), .A2(n_1092), .B1(n_1554), .B2(n_1557), .Y(n_1567) );
INVx5_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_SL g398 ( .A(n_394), .Y(n_398) );
BUFx3_ASAP7_75t_L g763 ( .A(n_394), .Y(n_763) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_395), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g1568 ( .A1(n_397), .A2(n_398), .B1(n_1551), .B2(n_1562), .Y(n_1568) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_398), .A2(n_1074), .B1(n_1086), .B2(n_1092), .Y(n_1094) );
OAI221xp5_ASAP7_75t_L g1514 ( .A1(n_398), .A2(n_1515), .B1(n_1516), .B2(n_1517), .C(n_1518), .Y(n_1514) );
BUFx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g532 ( .A(n_401), .Y(n_532) );
BUFx6f_ASAP7_75t_L g1522 ( .A(n_401), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_402), .A2(n_997), .B1(n_1073), .B2(n_1085), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_402), .A2(n_999), .B1(n_1078), .B2(n_1082), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g1569 ( .A1(n_402), .A2(n_1555), .B1(n_1559), .B2(n_1570), .Y(n_1569) );
INVx6_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI33xp33_ASAP7_75t_L g1087 ( .A1(n_404), .A2(n_1088), .A3(n_1090), .B1(n_1091), .B2(n_1094), .B3(n_1095), .Y(n_1087) );
OAI33xp33_ASAP7_75t_L g1137 ( .A1(n_404), .A2(n_1138), .A3(n_1139), .B1(n_1140), .B2(n_1141), .B3(n_1142), .Y(n_1137) );
OAI33xp33_ASAP7_75t_L g1564 ( .A1(n_404), .A2(n_1088), .A3(n_1565), .B1(n_1567), .B2(n_1568), .B3(n_1569), .Y(n_1564) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx1_ASAP7_75t_SL g502 ( .A(n_406), .Y(n_502) );
INVx4_ASAP7_75t_L g683 ( .A(n_406), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_406), .B(n_407), .Y(n_836) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI31xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_418), .A3(n_437), .B(n_443), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g729 ( .A(n_413), .Y(n_729) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_413), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1108 ( .A(n_413), .Y(n_1108) );
INVx1_ASAP7_75t_L g1196 ( .A(n_413), .Y(n_1196) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_415), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g808 ( .A(n_415), .Y(n_808) );
INVx2_ASAP7_75t_L g1012 ( .A(n_415), .Y(n_1012) );
INVx1_ASAP7_75t_L g1109 ( .A(n_415), .Y(n_1109) );
INVx1_ASAP7_75t_L g1580 ( .A(n_415), .Y(n_1580) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_417), .Y(n_581) );
INVx2_ASAP7_75t_L g695 ( .A(n_417), .Y(n_695) );
INVx1_ASAP7_75t_L g1081 ( .A(n_417), .Y(n_1081) );
BUFx6f_ASAP7_75t_L g1244 ( .A(n_417), .Y(n_1244) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_SL g885 ( .A(n_420), .Y(n_885) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND4xp25_ASAP7_75t_L g717 ( .A(n_422), .B(n_718), .C(n_722), .D(n_727), .Y(n_717) );
CKINVDCx8_ASAP7_75t_R g422 ( .A(n_423), .Y(n_422) );
CKINVDCx8_ASAP7_75t_R g803 ( .A(n_423), .Y(n_803) );
BUFx2_ASAP7_75t_L g579 ( .A(n_424), .Y(n_579) );
INVx2_ASAP7_75t_L g593 ( .A(n_424), .Y(n_593) );
BUFx2_ASAP7_75t_L g617 ( .A(n_424), .Y(n_617) );
BUFx2_ASAP7_75t_L g702 ( .A(n_424), .Y(n_702) );
BUFx2_ASAP7_75t_L g726 ( .A(n_424), .Y(n_726) );
BUFx2_ASAP7_75t_L g1038 ( .A(n_424), .Y(n_1038) );
INVx1_ASAP7_75t_L g585 ( .A(n_425), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_432), .B1(n_433), .B2(n_436), .Y(n_426) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_427), .A2(n_433), .B1(n_723), .B2(n_724), .C1(n_725), .C2(n_726), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g1582 ( .A1(n_427), .A2(n_433), .B1(n_1575), .B2(n_1583), .Y(n_1582) );
BUFx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_428), .Y(n_1015) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x4_ASAP7_75t_L g434 ( .A(n_429), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g805 ( .A(n_429), .B(n_431), .Y(n_805) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_432), .A2(n_467), .B1(n_470), .B2(n_475), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_433), .A2(n_964), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_433), .A2(n_1015), .B1(n_1100), .B2(n_1112), .Y(n_1111) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_434), .A2(n_785), .B1(n_805), .B2(n_806), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_434), .A2(n_805), .B1(n_887), .B2(n_888), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_434), .A2(n_805), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_434), .A2(n_805), .B1(n_1200), .B2(n_1201), .Y(n_1199) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g731 ( .A(n_439), .Y(n_731) );
BUFx2_ASAP7_75t_L g799 ( .A(n_439), .Y(n_799) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g721 ( .A(n_442), .Y(n_721) );
BUFx3_ASAP7_75t_L g809 ( .A(n_442), .Y(n_809) );
INVx1_ASAP7_75t_L g1115 ( .A(n_442), .Y(n_1115) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_446), .Y(n_443) );
AND2x4_ASAP7_75t_L g732 ( .A(n_444), .B(n_446), .Y(n_732) );
AND2x2_ASAP7_75t_SL g810 ( .A(n_444), .B(n_446), .Y(n_810) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OAI31xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_456), .A3(n_476), .B(n_482), .Y(n_448) );
CKINVDCx16_ASAP7_75t_R g450 ( .A(n_451), .Y(n_450) );
INVx4_ASAP7_75t_L g795 ( .A(n_451), .Y(n_795) );
INVx3_ASAP7_75t_SL g968 ( .A(n_451), .Y(n_968) );
AND2x4_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g501 ( .A(n_454), .Y(n_501) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_454), .Y(n_519) );
BUFx3_ASAP7_75t_L g930 ( .A(n_454), .Y(n_930) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx4_ASAP7_75t_L g782 ( .A(n_460), .Y(n_782) );
BUFx4f_ASAP7_75t_L g826 ( .A(n_460), .Y(n_826) );
BUFx4f_ASAP7_75t_L g864 ( .A(n_460), .Y(n_864) );
BUFx6f_ASAP7_75t_L g1191 ( .A(n_460), .Y(n_1191) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g783 ( .A(n_462), .Y(n_783) );
INVx1_ASAP7_75t_L g962 ( .A(n_462), .Y(n_962) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
BUFx3_ASAP7_75t_L g497 ( .A(n_464), .Y(n_497) );
AND2x6_ASAP7_75t_L g510 ( .A(n_464), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_SL g524 ( .A(n_464), .B(n_494), .Y(n_524) );
INVx1_ASAP7_75t_L g538 ( .A(n_464), .Y(n_538) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_464), .Y(n_661) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g676 ( .A(n_465), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_467), .A2(n_1100), .B1(n_1101), .B2(n_1103), .Y(n_1099) );
AND2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
AND2x4_ASAP7_75t_L g787 ( .A(n_468), .B(n_469), .Y(n_787) );
INVx1_ASAP7_75t_L g528 ( .A(n_469), .Y(n_528) );
BUFx2_ASAP7_75t_L g925 ( .A(n_469), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_470), .A2(n_785), .B1(n_786), .B2(n_788), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_470), .A2(n_786), .B1(n_1200), .B2(n_1208), .Y(n_1207) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx3_ASAP7_75t_L g895 ( .A(n_472), .Y(n_895) );
INVx2_ASAP7_75t_L g1102 ( .A(n_472), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1574 ( .A1(n_472), .A2(n_787), .B1(n_1575), .B2(n_1576), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_473), .B(n_511), .Y(n_561) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g791 ( .A(n_478), .Y(n_791) );
HB1xp67_ASAP7_75t_L g970 ( .A(n_478), .Y(n_970) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g971 ( .A(n_480), .Y(n_971) );
INVx2_ASAP7_75t_L g1105 ( .A(n_480), .Y(n_1105) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g793 ( .A(n_481), .Y(n_793) );
BUFx2_ASAP7_75t_L g898 ( .A(n_481), .Y(n_898) );
OAI31xp33_ASAP7_75t_L g779 ( .A1(n_482), .A2(n_780), .A3(n_789), .B(n_794), .Y(n_779) );
OAI31xp33_ASAP7_75t_L g1096 ( .A1(n_482), .A2(n_1097), .A3(n_1098), .B(n_1104), .Y(n_1096) );
OAI31xp33_ASAP7_75t_SL g1203 ( .A1(n_482), .A2(n_1204), .A3(n_1206), .B(n_1209), .Y(n_1203) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx2_ASAP7_75t_SL g900 ( .A(n_483), .Y(n_900) );
OAI31xp33_ASAP7_75t_L g960 ( .A1(n_483), .A2(n_961), .A3(n_966), .B(n_969), .Y(n_960) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g560 ( .A(n_485), .B(n_561), .Y(n_560) );
INVxp67_ASAP7_75t_L g570 ( .A(n_485), .Y(n_570) );
INVx1_ASAP7_75t_L g634 ( .A(n_485), .Y(n_634) );
INVx1_ASAP7_75t_L g619 ( .A(n_486), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_488), .B(n_546), .C(n_571), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_520), .B(n_541), .Y(n_488) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
INVx3_ASAP7_75t_L g1049 ( .A(n_491), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_491), .A2(n_518), .B1(n_1229), .B2(n_1230), .Y(n_1228) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_492), .Y(n_1058) );
INVx1_ASAP7_75t_L g1506 ( .A(n_492), .Y(n_1506) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g509 ( .A(n_493), .Y(n_509) );
BUFx3_ASAP7_75t_L g665 ( .A(n_493), .Y(n_665) );
BUFx3_ASAP7_75t_L g686 ( .A(n_493), .Y(n_686) );
AND2x2_ASAP7_75t_L g515 ( .A(n_494), .B(n_506), .Y(n_515) );
AND2x4_ASAP7_75t_L g518 ( .A(n_494), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g644 ( .A(n_494), .B(n_519), .Y(n_644) );
AND2x2_ASAP7_75t_L g688 ( .A(n_494), .B(n_508), .Y(n_688) );
AOI21xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_503), .B(n_510), .Y(n_495) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g765 ( .A(n_501), .Y(n_765) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g664 ( .A(n_505), .Y(n_664) );
INVx2_ASAP7_75t_SL g668 ( .A(n_505), .Y(n_668) );
INVx1_ASAP7_75t_L g685 ( .A(n_505), .Y(n_685) );
INVx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_506), .B(n_511), .Y(n_556) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_506), .Y(n_767) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI211xp5_ASAP7_75t_SL g771 ( .A1(n_510), .A2(n_690), .B(n_724), .C(n_772), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g1054 ( .A1(n_510), .A2(n_1055), .B(n_1057), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_510), .A2(n_690), .B1(n_1217), .B2(n_1218), .C(n_1219), .Y(n_1216) );
AOI21xp5_ASAP7_75t_L g1501 ( .A1(n_510), .A2(n_1502), .B(n_1503), .Y(n_1501) );
INVx1_ASAP7_75t_L g529 ( .A(n_511), .Y(n_529) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_511), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B1(n_516), .B2(n_517), .Y(n_512) );
INVx1_ASAP7_75t_L g757 ( .A(n_514), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_514), .A2(n_1051), .B1(n_1052), .B2(n_1053), .Y(n_1050) );
AOI221xp5_ASAP7_75t_SL g1220 ( .A1(n_514), .A2(n_1221), .B1(n_1223), .B2(n_1226), .C(n_1227), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x4_ASAP7_75t_L g633 ( .A(n_515), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g1509 ( .A(n_515), .Y(n_1509) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g760 ( .A(n_518), .Y(n_760) );
BUFx6f_ASAP7_75t_L g1053 ( .A(n_518), .Y(n_1053) );
HB1xp67_ASAP7_75t_L g1511 ( .A(n_518), .Y(n_1511) );
INVx1_ASAP7_75t_L g660 ( .A(n_519), .Y(n_660) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_519), .Y(n_682) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g938 ( .A(n_522), .Y(n_938) );
INVx2_ASAP7_75t_L g1060 ( .A(n_522), .Y(n_1060) );
INVx4_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx3_ASAP7_75t_L g690 ( .A(n_524), .Y(n_690) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g1061 ( .A(n_527), .Y(n_1061) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g672 ( .A(n_528), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_533), .B1(n_534), .B2(n_535), .C(n_536), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g662 ( .A(n_540), .Y(n_662) );
INVx1_ASAP7_75t_L g1222 ( .A(n_540), .Y(n_1222) );
INVx2_ASAP7_75t_L g1519 ( .A(n_540), .Y(n_1519) );
OAI21xp5_ASAP7_75t_SL g1047 ( .A1(n_541), .A2(n_1048), .B(n_1059), .Y(n_1047) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI21xp33_ASAP7_75t_L g754 ( .A1(n_542), .A2(n_755), .B(n_771), .Y(n_754) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g939 ( .A(n_543), .Y(n_939) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_544), .Y(n_1231) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_SL g1527 ( .A(n_545), .Y(n_1527) );
AOI21xp33_ASAP7_75t_SL g546 ( .A1(n_547), .A2(n_557), .B(n_558), .Y(n_546) );
AOI21xp33_ASAP7_75t_L g1042 ( .A1(n_547), .A2(n_1043), .B(n_1044), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g1250 ( .A1(n_547), .A2(n_1251), .B(n_1252), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_547), .B(n_1532), .Y(n_1531) );
INVx8_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_549), .B(n_554), .Y(n_548) );
INVx1_ASAP7_75t_L g653 ( .A(n_549), .Y(n_653) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_551), .Y(n_738) );
OR2x2_ASAP7_75t_L g562 ( .A(n_552), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g609 ( .A(n_552), .Y(n_609) );
INVx1_ASAP7_75t_L g612 ( .A(n_552), .Y(n_612) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
AND2x4_ASAP7_75t_L g599 ( .A(n_555), .B(n_568), .Y(n_599) );
INVx2_ASAP7_75t_L g1213 ( .A(n_559), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1529 ( .A(n_559), .Y(n_1529) );
AND2x4_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
AND2x4_ASAP7_75t_L g1045 ( .A(n_560), .B(n_562), .Y(n_1045) );
INVx1_ASAP7_75t_L g774 ( .A(n_561), .Y(n_774) );
INVx2_ASAP7_75t_L g655 ( .A(n_562), .Y(n_655) );
INVx3_ASAP7_75t_L g802 ( .A(n_563), .Y(n_802) );
INVx4_ASAP7_75t_L g947 ( .A(n_563), .Y(n_947) );
BUFx6f_ASAP7_75t_L g981 ( .A(n_563), .Y(n_981) );
INVx3_ASAP7_75t_L g628 ( .A(n_564), .Y(n_628) );
INVx5_ASAP7_75t_L g1256 ( .A(n_564), .Y(n_1256) );
OR2x6_ASAP7_75t_L g564 ( .A(n_565), .B(n_570), .Y(n_564) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_565), .B(n_570), .Y(n_1046) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
BUFx3_ASAP7_75t_L g578 ( .A(n_566), .Y(n_578) );
BUFx3_ASAP7_75t_L g701 ( .A(n_566), .Y(n_701) );
INVx8_ASAP7_75t_L g710 ( .A(n_566), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_605), .C(n_614), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_573), .B(n_594), .Y(n_572) );
AOI33xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .A3(n_580), .B1(n_586), .B2(n_588), .B3(n_591), .Y(n_573) );
BUFx3_ASAP7_75t_L g955 ( .A(n_574), .Y(n_955) );
AOI33xp33_ASAP7_75t_L g1032 ( .A1(n_574), .A2(n_588), .A3(n_1033), .B1(n_1034), .B2(n_1036), .B3(n_1037), .Y(n_1032) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
BUFx3_ASAP7_75t_L g741 ( .A(n_578), .Y(n_741) );
INVx1_ASAP7_75t_L g750 ( .A(n_578), .Y(n_750) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_R g1035 ( .A(n_583), .Y(n_1035) );
INVx5_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx3_ASAP7_75t_L g587 ( .A(n_584), .Y(n_587) );
BUFx12f_ASAP7_75t_L g707 ( .A(n_584), .Y(n_707) );
BUFx3_ASAP7_75t_L g942 ( .A(n_584), .Y(n_942) );
INVx1_ASAP7_75t_L g604 ( .A(n_585), .Y(n_604) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g711 ( .A(n_593), .Y(n_711) );
INVx1_ASAP7_75t_L g742 ( .A(n_593), .Y(n_742) );
INVx2_ASAP7_75t_L g1249 ( .A(n_593), .Y(n_1249) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_600), .B2(n_601), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_596), .A2(n_601), .B1(n_1040), .B2(n_1041), .Y(n_1039) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
AND2x4_ASAP7_75t_SL g648 ( .A(n_597), .B(n_599), .Y(n_648) );
NAND2x1_ASAP7_75t_L g913 ( .A(n_597), .B(n_599), .Y(n_913) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g601 ( .A(n_599), .B(n_602), .Y(n_601) );
AND2x4_ASAP7_75t_L g616 ( .A(n_599), .B(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_SL g650 ( .A(n_599), .B(n_602), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g911 ( .A1(n_601), .A2(n_912), .B1(n_914), .B2(n_915), .C(n_916), .Y(n_911) );
AOI221xp5_ASAP7_75t_L g1253 ( .A1(n_601), .A2(n_616), .B1(n_648), .B2(n_1219), .C(n_1254), .Y(n_1253) );
HB1xp67_ASAP7_75t_L g1488 ( .A(n_601), .Y(n_1488) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
OR2x6_ASAP7_75t_L g635 ( .A(n_607), .B(n_608), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_607), .A2(n_851), .B1(n_859), .B2(n_866), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g879 ( .A1(n_607), .A2(n_801), .B1(n_860), .B2(n_867), .Y(n_879) );
INVx2_ASAP7_75t_SL g977 ( .A(n_607), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g1170 ( .A1(n_607), .A2(n_954), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
OAI22xp33_ASAP7_75t_L g1180 ( .A1(n_607), .A2(n_1181), .B1(n_1182), .B2(n_1183), .Y(n_1180) );
INVxp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g639 ( .A(n_609), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1530 ( .A1(n_611), .A2(n_1258), .B1(n_1510), .B2(n_1512), .Y(n_1530) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x4_ASAP7_75t_L g1258 ( .A(n_612), .B(n_1259), .Y(n_1258) );
INVx3_ASAP7_75t_L g845 ( .A(n_613), .Y(n_845) );
INVx3_ASAP7_75t_L g847 ( .A(n_613), .Y(n_847) );
INVx2_ASAP7_75t_SL g950 ( .A(n_613), .Y(n_950) );
NOR3xp33_ASAP7_75t_L g1029 ( .A(n_614), .B(n_1030), .C(n_1031), .Y(n_1029) );
INVx2_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_615), .A2(n_694), .B(n_703), .C(n_704), .Y(n_693) );
AND4x1_ASAP7_75t_L g1484 ( .A(n_615), .B(n_1485), .C(n_1489), .D(n_1491), .Y(n_1484) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
XOR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_903), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_623), .B1(n_776), .B2(n_902), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
XOR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_714), .Y(n_623) );
INVx1_ASAP7_75t_L g712 ( .A(n_625), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .C(n_645), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_627), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_631), .B1(n_636), .B2(n_637), .Y(n_629) );
INVxp67_ASAP7_75t_L g908 ( .A(n_631), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_L g643 ( .A(n_634), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g909 ( .A(n_637), .Y(n_909) );
NAND2x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g706 ( .A(n_641), .Y(n_706) );
BUFx2_ASAP7_75t_L g744 ( .A(n_641), .Y(n_744) );
BUFx2_ASAP7_75t_L g1175 ( .A(n_641), .Y(n_1175) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NOR3xp33_ASAP7_75t_SL g645 ( .A(n_646), .B(n_656), .C(n_693), .Y(n_645) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_654), .B2(n_655), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_652), .B(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_654), .A2(n_670), .B1(n_672), .B2(n_673), .C(n_674), .Y(n_669) );
AOI31xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_679), .A3(n_687), .B(n_691), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_663), .B(n_666), .Y(n_657) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_669), .B(n_677), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_670), .A2(n_914), .B1(n_925), .B2(n_926), .Y(n_924) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
A2O1A1Ixp33_ASAP7_75t_L g919 ( .A1(n_678), .A2(n_920), .B(n_921), .C(n_922), .Y(n_919) );
INVx2_ASAP7_75t_L g758 ( .A(n_688), .Y(n_758) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI33xp33_ASAP7_75t_L g842 ( .A1(n_703), .A2(n_753), .A3(n_843), .B1(n_844), .B2(n_846), .B3(n_848), .Y(n_842) );
OAI33xp33_ASAP7_75t_L g871 ( .A1(n_703), .A2(n_872), .A3(n_873), .B1(n_875), .B2(n_878), .B3(n_879), .Y(n_871) );
INVx1_ASAP7_75t_L g735 ( .A(n_706), .Y(n_735) );
INVx1_ASAP7_75t_L g1558 ( .A(n_706), .Y(n_1558) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g1259 ( .A(n_710), .Y(n_1259) );
INVx8_ASAP7_75t_L g1498 ( .A(n_710), .Y(n_1498) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_732), .B(n_733), .C(n_754), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_725), .B(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g752 ( .A(n_726), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_729), .B1(n_730), .B2(n_731), .Y(n_727) );
INVx2_ASAP7_75t_L g798 ( .A(n_729), .Y(n_798) );
INVx2_ASAP7_75t_L g882 ( .A(n_731), .Y(n_882) );
INVx1_ASAP7_75t_L g1018 ( .A(n_731), .Y(n_1018) );
OAI31xp33_ASAP7_75t_L g880 ( .A1(n_732), .A2(n_881), .A3(n_883), .B(n_889), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_737), .B2(n_739), .C(n_740), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g1130 ( .A1(n_735), .A2(n_979), .B1(n_1131), .B2(n_1132), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_737), .A2(n_874), .B1(n_1077), .B2(n_1078), .Y(n_1076) );
CKINVDCx8_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
INVx3_ASAP7_75t_L g746 ( .A(n_738), .Y(n_746) );
INVx3_ASAP7_75t_L g985 ( .A(n_738), .Y(n_985) );
INVx3_ASAP7_75t_L g1083 ( .A(n_738), .Y(n_1083) );
INVx1_ASAP7_75t_L g1246 ( .A(n_738), .Y(n_1246) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_747), .C(n_748), .Y(n_743) );
OAI211xp5_ASAP7_75t_SL g768 ( .A1(n_745), .A2(n_763), .B(n_769), .C(n_770), .Y(n_768) );
OAI22xp5_ASAP7_75t_L g846 ( .A1(n_746), .A2(n_825), .B1(n_841), .B2(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_756), .B(n_759), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B(n_764), .C(n_766), .Y(n_761) );
BUFx2_ASAP7_75t_L g892 ( .A(n_763), .Y(n_892) );
BUFx6f_ASAP7_75t_L g921 ( .A(n_767), .Y(n_921) );
INVx3_ASAP7_75t_L g1225 ( .A(n_767), .Y(n_1225) );
INVx1_ASAP7_75t_L g902 ( .A(n_776), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_852), .B1(n_853), .B2(n_901), .Y(n_776) );
INVx1_ASAP7_75t_L g901 ( .A(n_777), .Y(n_901) );
NAND3xp33_ASAP7_75t_SL g778 ( .A(n_779), .B(n_796), .C(n_811), .Y(n_778) );
OAI211xp5_ASAP7_75t_L g927 ( .A1(n_781), .A2(n_928), .B(n_929), .C(n_931), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g1142 ( .A1(n_781), .A2(n_1129), .B1(n_1132), .B2(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g832 ( .A(n_782), .Y(n_832) );
INVx1_ASAP7_75t_L g923 ( .A(n_782), .Y(n_923) );
INVx2_ASAP7_75t_L g934 ( .A(n_782), .Y(n_934) );
INVx2_ASAP7_75t_L g1188 ( .A(n_782), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_786), .A2(n_887), .B1(n_894), .B2(n_895), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_786), .A2(n_895), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_786), .A2(n_895), .B1(n_1151), .B2(n_1161), .Y(n_1160) );
BUFx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OAI31xp33_ASAP7_75t_SL g796 ( .A1(n_797), .A2(n_800), .A3(n_807), .B(n_810), .Y(n_796) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_801), .A2(n_945), .B1(n_1085), .B2(n_1086), .Y(n_1084) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g954 ( .A(n_802), .Y(n_954) );
OAI31xp33_ASAP7_75t_L g1008 ( .A1(n_810), .A2(n_1009), .A3(n_1013), .B(n_1017), .Y(n_1008) );
OAI31xp33_ASAP7_75t_L g1106 ( .A1(n_810), .A2(n_1107), .A3(n_1110), .B(n_1113), .Y(n_1106) );
OAI31xp33_ASAP7_75t_SL g1147 ( .A1(n_810), .A2(n_1148), .A3(n_1149), .B(n_1153), .Y(n_1147) );
OAI31xp33_ASAP7_75t_L g1193 ( .A1(n_810), .A2(n_1194), .A3(n_1197), .B(n_1202), .Y(n_1193) );
OAI31xp33_ASAP7_75t_L g1578 ( .A1(n_810), .A2(n_1579), .A3(n_1581), .B(n_1584), .Y(n_1578) );
NOR2xp33_ASAP7_75t_SL g811 ( .A(n_812), .B(n_842), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B1(n_818), .B2(n_819), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_815), .A2(n_838), .B1(n_839), .B2(n_841), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_815), .A2(n_819), .B1(n_859), .B2(n_860), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_815), .A2(n_839), .B1(n_869), .B2(n_870), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_815), .A2(n_819), .B1(n_1122), .B2(n_1135), .Y(n_1139) );
OAI22xp33_ASAP7_75t_L g1185 ( .A1(n_815), .A2(n_839), .B1(n_1171), .B2(n_1181), .Y(n_1185) );
OAI22xp33_ASAP7_75t_L g1192 ( .A1(n_815), .A2(n_839), .B1(n_1176), .B2(n_1179), .Y(n_1192) );
INVx2_ASAP7_75t_SL g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g1566 ( .A(n_816), .Y(n_1566) );
INVx2_ASAP7_75t_L g1570 ( .A(n_816), .Y(n_1570) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx3_ASAP7_75t_L g999 ( .A(n_817), .Y(n_999) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_818), .A2(n_833), .B1(n_849), .B2(n_851), .Y(n_848) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_819), .A2(n_828), .B1(n_1123), .B2(n_1136), .Y(n_1141) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_824), .B1(n_825), .B2(n_826), .Y(n_822) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_824), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g1140 ( .A1(n_824), .A2(n_864), .B1(n_1125), .B2(n_1131), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_826), .A2(n_983), .B1(n_987), .B2(n_1004), .Y(n_1003) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_826), .A2(n_978), .B1(n_994), .B2(n_1004), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_828), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_827) );
INVx3_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
OAI211xp5_ASAP7_75t_SL g1062 ( .A1(n_832), .A2(n_1063), .B(n_1064), .C(n_1065), .Y(n_1062) );
OAI33xp33_ASAP7_75t_L g1184 ( .A1(n_834), .A2(n_1088), .A3(n_1185), .B1(n_1186), .B2(n_1189), .B3(n_1192), .Y(n_1184) );
INVx2_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OAI33xp33_ASAP7_75t_L g856 ( .A1(n_836), .A2(n_857), .A3(n_858), .B1(n_861), .B2(n_865), .B3(n_868), .Y(n_856) );
BUFx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_847), .A2(n_985), .B1(n_987), .B2(n_988), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g1121 ( .A1(n_849), .A2(n_851), .B1(n_1122), .B2(n_1123), .Y(n_1121) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_850), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_951) );
HB1xp67_ASAP7_75t_L g1134 ( .A(n_850), .Y(n_1134) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_851), .A2(n_1237), .B1(n_1238), .B2(n_1241), .Y(n_1236) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_880), .C(n_890), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_871), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_863), .A2(n_870), .B1(n_876), .B2(n_877), .Y(n_875) );
OAI22xp5_ASAP7_75t_L g982 ( .A1(n_876), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
OAI22xp33_ASAP7_75t_SL g1124 ( .A1(n_877), .A2(n_1125), .B1(n_1126), .B2(n_1129), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
OAI31xp33_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_896), .A3(n_899), .B(n_900), .Y(n_890) );
HB1xp67_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_SL g1158 ( .A(n_898), .Y(n_1158) );
OAI31xp33_ASAP7_75t_L g1154 ( .A1(n_900), .A2(n_1155), .A3(n_1156), .B(n_1159), .Y(n_1154) );
OAI31xp33_ASAP7_75t_L g1571 ( .A1(n_900), .A2(n_1572), .A3(n_1573), .B(n_1577), .Y(n_1571) );
AO22x2_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_956), .B1(n_957), .B2(n_1020), .Y(n_903) );
INVx1_ASAP7_75t_SL g1020 ( .A(n_904), .Y(n_1020) );
XNOR2x1_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
NOR2x1_ASAP7_75t_L g906 ( .A(n_907), .B(n_910), .Y(n_906) );
NAND3xp33_ASAP7_75t_SL g910 ( .A(n_911), .B(n_917), .C(n_940), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_912), .A2(n_1486), .B1(n_1487), .B2(n_1488), .Y(n_1485) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
OAI21xp5_ASAP7_75t_L g917 ( .A1(n_918), .A2(n_937), .B(n_939), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_927), .C(n_932), .Y(n_918) );
HB1xp67_ASAP7_75t_L g1504 ( .A(n_921), .Y(n_1504) );
NAND2xp5_ASAP7_75t_SL g922 ( .A(n_923), .B(n_924), .Y(n_922) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_930), .Y(n_1056) );
OAI211xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B(n_935), .C(n_936), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_933), .A2(n_944), .B1(n_945), .B2(n_946), .Y(n_943) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g1198 ( .A(n_947), .Y(n_1198) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_950), .A2(n_985), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AOI33xp33_ASAP7_75t_L g1491 ( .A1(n_955), .A2(n_990), .A3(n_1492), .B1(n_1493), .B2(n_1495), .B3(n_1496), .Y(n_1491) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_972), .C(n_1008), .Y(n_959) );
NOR2xp33_ASAP7_75t_SL g972 ( .A(n_973), .B(n_995), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g974 ( .A1(n_975), .A2(n_976), .B1(n_978), .B2(n_979), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g996 ( .A1(n_975), .A2(n_993), .B1(n_997), .B2(n_1000), .Y(n_996) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVx2_ASAP7_75t_SL g979 ( .A(n_980), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
HB1xp67_ASAP7_75t_L g1075 ( .A(n_981), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_981), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_984), .A2(n_988), .B1(n_997), .B2(n_1000), .Y(n_1007) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
BUFx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx2_ASAP7_75t_SL g998 ( .A(n_999), .Y(n_998) );
INVx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
OAI22xp33_ASAP7_75t_SL g1189 ( .A1(n_1004), .A2(n_1172), .B1(n_1183), .B2(n_1190), .Y(n_1189) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1093 ( .A(n_1005), .Y(n_1093) );
INVx2_ASAP7_75t_L g1187 ( .A(n_1005), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1010 ( .A(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1024), .B1(n_1164), .B2(n_1261), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_1025), .A2(n_1026), .B1(n_1066), .B2(n_1163), .Y(n_1024) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
AND3x1_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1042), .C(n_1047), .Y(n_1028) );
NAND2xp5_ASAP7_75t_SL g1031 ( .A(n_1032), .B(n_1039), .Y(n_1031) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1066), .Y(n_1163) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1116), .B1(n_1117), .B2(n_1162), .Y(n_1066) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1067), .Y(n_1162) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
AND3x1_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1096), .C(n_1106), .Y(n_1069) );
NOR2xp33_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1087), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1083), .A2(n_1134), .B1(n_1135), .B2(n_1136), .Y(n_1133) );
OAI22xp5_ASAP7_75t_L g1173 ( .A1(n_1083), .A2(n_1174), .B1(n_1175), .B2(n_1176), .Y(n_1173) );
BUFx6f_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx4_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx2_ASAP7_75t_SL g1116 ( .A(n_1117), .Y(n_1116) );
NAND3xp33_ASAP7_75t_L g1118 ( .A(n_1119), .B(n_1147), .C(n_1154), .Y(n_1118) );
NOR2xp33_ASAP7_75t_SL g1119 ( .A(n_1120), .B(n_1137), .Y(n_1119) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1164), .Y(n_1261) );
HB1xp67_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
XNOR2xp5_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1210), .Y(n_1165) );
NAND3xp33_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1193), .C(n_1203), .Y(n_1167) );
NOR2xp33_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1184), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_1174), .A2(n_1178), .B1(n_1187), .B2(n_1188), .Y(n_1186) );
HB1xp67_ASAP7_75t_L g1190 ( .A(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
XNOR2xp5_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1260), .Y(n_1210) );
NAND2xp5_ASAP7_75t_SL g1211 ( .A(n_1212), .B(n_1250), .Y(n_1211) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1213), .A2(n_1214), .B1(n_1215), .B2(n_1231), .C(n_1232), .Y(n_1212) );
NAND3xp33_ASAP7_75t_L g1215 ( .A(n_1216), .B(n_1220), .C(n_1228), .Y(n_1215) );
INVx2_ASAP7_75t_SL g1224 ( .A(n_1225), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1257 ( .A(n_1226), .B(n_1258), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1255 ( .A(n_1230), .B(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1239 ( .A(n_1240), .Y(n_1239) );
OAI221xp5_ASAP7_75t_L g1242 ( .A1(n_1243), .A2(n_1245), .B1(n_1246), .B2(n_1247), .C(n_1248), .Y(n_1242) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
NAND3xp33_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1255), .C(n_1257), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1256), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OAI221xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1478), .B1(n_1481), .B2(n_1534), .C(n_1537), .Y(n_1264) );
AOI21xp5_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1369), .B(n_1390), .Y(n_1265) );
OAI211xp5_ASAP7_75t_L g1266 ( .A1(n_1267), .A2(n_1286), .B(n_1317), .C(n_1355), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1282), .Y(n_1267) );
INVx3_ASAP7_75t_L g1326 ( .A(n_1268), .Y(n_1326) );
INVx3_ASAP7_75t_L g1366 ( .A(n_1268), .Y(n_1366) );
NOR2xp33_ASAP7_75t_L g1368 ( .A(n_1268), .B(n_1343), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1268), .B(n_1389), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1268), .B(n_1411), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1268), .B(n_1282), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1268), .B(n_1335), .Y(n_1435) );
AND2x4_ASAP7_75t_SL g1268 ( .A(n_1269), .B(n_1276), .Y(n_1268) );
AND2x6_ASAP7_75t_L g1270 ( .A(n_1271), .B(n_1272), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1274 ( .A(n_1271), .B(n_1275), .Y(n_1274) );
AND2x4_ASAP7_75t_L g1277 ( .A(n_1271), .B(n_1278), .Y(n_1277) );
AND2x6_ASAP7_75t_L g1280 ( .A(n_1271), .B(n_1281), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1271), .B(n_1275), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1271), .B(n_1275), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1273), .B(n_1279), .Y(n_1278) );
INVx2_ASAP7_75t_L g1480 ( .A(n_1280), .Y(n_1480) );
OAI21xp5_ASAP7_75t_L g1586 ( .A1(n_1281), .A2(n_1587), .B(n_1588), .Y(n_1586) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1282), .B(n_1311), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1282), .B(n_1366), .Y(n_1365) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1282), .B(n_1310), .Y(n_1374) );
OR2x2_ASAP7_75t_L g1382 ( .A(n_1282), .B(n_1311), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1282), .B(n_1397), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1283), .B(n_1285), .Y(n_1282) );
AND2x4_ASAP7_75t_L g1330 ( .A(n_1283), .B(n_1285), .Y(n_1330) );
AOI211xp5_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1295), .B(n_1303), .C(n_1308), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1287), .B(n_1347), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1287), .B(n_1342), .Y(n_1412) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1287), .B(n_1307), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1291), .Y(n_1287) );
INVx3_ASAP7_75t_L g1306 ( .A(n_1288), .Y(n_1306) );
INVx2_ASAP7_75t_L g1339 ( .A(n_1288), .Y(n_1339) );
NOR2xp33_ASAP7_75t_L g1373 ( .A(n_1288), .B(n_1291), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1288), .B(n_1423), .Y(n_1422) );
OR2x2_ASAP7_75t_L g1438 ( .A(n_1288), .B(n_1310), .Y(n_1438) );
NOR2xp33_ASAP7_75t_L g1458 ( .A(n_1288), .B(n_1459), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1290), .Y(n_1288) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1291), .B(n_1334), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1291), .B(n_1316), .Y(n_1340) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_1291), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1291), .B(n_1350), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1291), .B(n_1357), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1291), .B(n_1347), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1294), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1292), .B(n_1294), .Y(n_1319) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1295), .Y(n_1342) );
NOR2xp33_ASAP7_75t_L g1442 ( .A(n_1295), .B(n_1306), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1299), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1296), .B(n_1299), .Y(n_1307) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1296), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1296), .B(n_1300), .Y(n_1347) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1296), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1297), .B(n_1298), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1299), .B(n_1316), .Y(n_1315) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1299), .Y(n_1334) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1300), .Y(n_1350) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1302), .Y(n_1300) );
INVxp67_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1307), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1305), .B(n_1333), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1305), .B(n_1335), .Y(n_1352) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
NAND2xp5_ASAP7_75t_L g1309 ( .A(n_1306), .B(n_1310), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1306), .B(n_1307), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1306), .B(n_1362), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1306), .B(n_1402), .Y(n_1424) );
OAI21xp33_ASAP7_75t_L g1427 ( .A1(n_1306), .A2(n_1418), .B(n_1428), .Y(n_1427) );
NOR2xp33_ASAP7_75t_L g1446 ( .A(n_1306), .B(n_1447), .Y(n_1446) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1306), .B(n_1462), .Y(n_1461) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1307), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1307), .B(n_1373), .Y(n_1409) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1314), .Y(n_1308) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1309), .Y(n_1477) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1310), .B(n_1330), .Y(n_1329) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1311), .Y(n_1344) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1311), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
NOR3xp33_ASAP7_75t_L g1437 ( .A(n_1314), .B(n_1366), .C(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1315), .B(n_1351), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1315), .B(n_1435), .Y(n_1434) );
OAI32xp33_ASAP7_75t_L g1317 ( .A1(n_1318), .A2(n_1321), .A3(n_1325), .B1(n_1327), .B2(n_1353), .Y(n_1317) );
AOI332xp33_ASAP7_75t_L g1443 ( .A1(n_1318), .A2(n_1326), .A3(n_1383), .B1(n_1389), .B2(n_1411), .B3(n_1444), .C1(n_1446), .C2(n_1448), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1319), .B(n_1320), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1319), .B(n_1342), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1418 ( .A(n_1319), .B(n_1387), .Y(n_1418) );
AOI22xp5_ASAP7_75t_SL g1328 ( .A1(n_1320), .A2(n_1329), .B1(n_1331), .B2(n_1335), .Y(n_1328) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1321), .Y(n_1354) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1321), .B(n_1326), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_1321), .A2(n_1322), .B1(n_1457), .B2(n_1465), .Y(n_1456) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
AOI211xp5_ASAP7_75t_L g1371 ( .A1(n_1322), .A2(n_1372), .B(n_1374), .C(n_1375), .Y(n_1371) );
O2A1O1Ixp33_ASAP7_75t_SL g1413 ( .A1(n_1322), .A2(n_1414), .B(n_1415), .C(n_1416), .Y(n_1413) );
O2A1O1Ixp33_ASAP7_75t_L g1420 ( .A1(n_1322), .A2(n_1421), .B(n_1431), .C(n_1439), .Y(n_1420) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1322), .Y(n_1449) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1324), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1325), .B(n_1354), .Y(n_1353) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g1369 ( .A1(n_1326), .A2(n_1370), .B1(n_1371), .B2(n_1378), .C(n_1379), .Y(n_1369) );
AOI22xp5_ASAP7_75t_L g1454 ( .A1(n_1326), .A2(n_1455), .B1(n_1456), .B2(n_1469), .Y(n_1454) );
INVxp67_ASAP7_75t_SL g1370 ( .A(n_1327), .Y(n_1370) );
NAND4xp25_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1336), .C(n_1345), .D(n_1348), .Y(n_1327) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1329), .B(n_1346), .Y(n_1345) );
NAND2xp5_ASAP7_75t_SL g1359 ( .A(n_1329), .B(n_1339), .Y(n_1359) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1329), .Y(n_1414) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1330), .Y(n_1389) );
CKINVDCx6p67_ASAP7_75t_R g1394 ( .A(n_1330), .Y(n_1394) );
NOR2xp33_ASAP7_75t_L g1448 ( .A(n_1330), .B(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
AOI21xp33_ASAP7_75t_L g1463 ( .A1(n_1332), .A2(n_1338), .B(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1333), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1334), .B(n_1351), .Y(n_1362) );
CKINVDCx14_ASAP7_75t_R g1464 ( .A(n_1335), .Y(n_1464) );
OAI21xp5_ASAP7_75t_L g1336 ( .A1(n_1337), .A2(n_1341), .B(n_1343), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_1337), .A2(n_1426), .B1(n_1427), .B2(n_1429), .Y(n_1425) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1340), .Y(n_1338) );
INVx2_ASAP7_75t_L g1397 ( .A(n_1339), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1339), .B(n_1445), .Y(n_1444) );
NAND2xp5_ASAP7_75t_SL g1453 ( .A(n_1339), .B(n_1342), .Y(n_1453) );
CKINVDCx14_ASAP7_75t_R g1403 ( .A(n_1340), .Y(n_1403) );
CKINVDCx5p33_ASAP7_75t_R g1433 ( .A(n_1341), .Y(n_1433) );
OAI21xp5_ASAP7_75t_L g1348 ( .A1(n_1342), .A2(n_1349), .B(n_1352), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1342), .B(n_1373), .Y(n_1372) );
OAI21xp5_ASAP7_75t_L g1416 ( .A1(n_1342), .A2(n_1352), .B(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1343), .Y(n_1377) );
OAI21xp33_ASAP7_75t_L g1450 ( .A1(n_1343), .A2(n_1388), .B(n_1451), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1343), .B(n_1468), .Y(n_1467) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
OAI21xp5_ASAP7_75t_SL g1408 ( .A1(n_1344), .A2(n_1409), .B(n_1410), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1346), .B(n_1377), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1347), .B(n_1351), .Y(n_1402) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1347), .Y(n_1459) );
INVx1_ASAP7_75t_L g1428 ( .A(n_1349), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1350), .B(n_1351), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1351), .B(n_1387), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1351), .B(n_1442), .Y(n_1441) );
OR2x2_ASAP7_75t_L g1452 ( .A(n_1351), .B(n_1453), .Y(n_1452) );
A2O1A1Ixp33_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1358), .B(n_1360), .C(n_1363), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1357), .B(n_1373), .Y(n_1415) );
INVxp67_ASAP7_75t_L g1358 ( .A(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1367), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
OR2x2_ASAP7_75t_L g1381 ( .A(n_1366), .B(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
NOR2xp33_ASAP7_75t_L g1406 ( .A(n_1374), .B(n_1407), .Y(n_1406) );
A2O1A1Ixp33_ASAP7_75t_L g1421 ( .A1(n_1374), .A2(n_1422), .B(n_1424), .C(n_1425), .Y(n_1421) );
INVx2_ASAP7_75t_SL g1462 ( .A(n_1374), .Y(n_1462) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
AOI211xp5_ASAP7_75t_L g1391 ( .A1(n_1378), .A2(n_1392), .B(n_1413), .C(n_1419), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1379 ( .A1(n_1380), .A2(n_1383), .B1(n_1385), .B2(n_1388), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1419 ( .A(n_1381), .B(n_1386), .Y(n_1419) );
OAI211xp5_ASAP7_75t_SL g1439 ( .A1(n_1381), .A2(n_1440), .B(n_1443), .C(n_1450), .Y(n_1439) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1382), .Y(n_1445) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1460 ( .A(n_1387), .B(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1388), .Y(n_1432) );
A2O1A1Ixp33_ASAP7_75t_L g1469 ( .A1(n_1389), .A2(n_1412), .B(n_1470), .C(n_1471), .Y(n_1469) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_1389), .A2(n_1462), .B1(n_1472), .B2(n_1473), .C(n_1476), .Y(n_1471) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_1391), .B(n_1420), .C(n_1454), .Y(n_1390) );
OAI211xp5_ASAP7_75t_L g1392 ( .A1(n_1393), .A2(n_1395), .B(n_1399), .C(n_1408), .Y(n_1392) );
CKINVDCx6p67_ASAP7_75t_R g1393 ( .A(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
AOI211xp5_ASAP7_75t_L g1465 ( .A1(n_1396), .A2(n_1411), .B(n_1466), .C(n_1467), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1398), .Y(n_1396) );
NOR2xp33_ASAP7_75t_L g1466 ( .A(n_1397), .B(n_1447), .Y(n_1466) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1398), .Y(n_1407) );
AOI21xp5_ASAP7_75t_L g1399 ( .A1(n_1400), .A2(n_1404), .B(n_1406), .Y(n_1399) );
NAND2xp5_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1403), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1402), .B(n_1477), .Y(n_1476) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1412), .Y(n_1410) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1424), .Y(n_1472) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
OAI211xp5_ASAP7_75t_L g1431 ( .A1(n_1432), .A2(n_1433), .B(n_1434), .C(n_1436), .Y(n_1431) );
INVxp67_ASAP7_75t_SL g1436 ( .A(n_1437), .Y(n_1436) );
NAND2xp5_ASAP7_75t_SL g1473 ( .A(n_1440), .B(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
AOI211xp5_ASAP7_75t_L g1457 ( .A1(n_1445), .A2(n_1458), .B(n_1460), .C(n_1463), .Y(n_1457) );
INVxp67_ASAP7_75t_L g1455 ( .A(n_1448), .Y(n_1455) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1467), .Y(n_1470) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
CKINVDCx20_ASAP7_75t_R g1478 ( .A(n_1479), .Y(n_1478) );
CKINVDCx20_ASAP7_75t_R g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
XOR2x2_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1533), .Y(n_1482) );
NAND3x1_ASAP7_75t_SL g1483 ( .A(n_1484), .B(n_1499), .C(n_1531), .Y(n_1483) );
BUFx2_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
O2A1O1Ixp5_ASAP7_75t_L g1499 ( .A1(n_1500), .A2(n_1513), .B(n_1527), .C(n_1528), .Y(n_1499) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1506), .Y(n_1505) );
AOI22xp33_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1510), .B1(n_1511), .B2(n_1512), .Y(n_1507) );
INVx2_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1519), .Y(n_1518) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_1521), .A2(n_1522), .B1(n_1523), .B2(n_1526), .Y(n_1520) );
BUFx2_ASAP7_75t_L g1523 ( .A(n_1524), .Y(n_1523) );
BUFx6f_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
INVx2_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
HB1xp67_ASAP7_75t_SL g1538 ( .A(n_1539), .Y(n_1538) );
BUFx3_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVxp33_ASAP7_75t_SL g1541 ( .A(n_1542), .Y(n_1541) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1544), .Y(n_1543) );
HB1xp67_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
AND3x1_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1571), .C(n_1578), .Y(n_1545) );
NOR2xp33_ASAP7_75t_L g1546 ( .A(n_1547), .B(n_1564), .Y(n_1546) );
HB1xp67_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
endmodule