module real_jpeg_29067_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_300, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_300;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_286;
wire n_292;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_293;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_167;
wire n_202;
wire n_216;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_72),
.B1(n_73),
.B2(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_0),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_97),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_0),
.A2(n_32),
.B1(n_35),
.B2(n_97),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_97),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_1),
.A2(n_32),
.B1(n_35),
.B2(n_53),
.Y(n_225)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_2),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_3),
.B(n_26),
.Y(n_132)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_3),
.A2(n_25),
.B(n_26),
.C(n_132),
.D(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_3),
.B(n_48),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_3),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_3),
.A2(n_83),
.B(n_149),
.Y(n_169)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_3),
.A2(n_44),
.B(n_47),
.C(n_182),
.D(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_3),
.B(n_44),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_3),
.B(n_68),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_3),
.A2(n_70),
.B(n_73),
.C(n_227),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_72),
.B1(n_73),
.B2(n_164),
.Y(n_232)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_40),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_5),
.A2(n_32),
.B1(n_35),
.B2(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_8),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_75),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_75),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_75),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_144),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_9),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_9),
.A2(n_32),
.B1(n_35),
.B2(n_144),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_144),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_9),
.A2(n_72),
.B1(n_73),
.B2(n_144),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_10),
.A2(n_72),
.B1(n_73),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_10),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_32),
.B1(n_35),
.B2(n_119),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_119),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_119),
.Y(n_238)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_11),
.B(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_11),
.A2(n_29),
.B1(n_32),
.B2(n_35),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_32),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_37),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_13),
.A2(n_46),
.B1(n_72),
.B2(n_73),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_46),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_13),
.A2(n_32),
.B1(n_35),
.B2(n_46),
.Y(n_209)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

XNOR2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_121),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_80),
.B2(n_81),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_54),
.B1(n_55),
.B2(n_79),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_23),
.A2(n_24),
.B(n_41),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_38),
.Y(n_24)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_25),
.A2(n_31),
.B1(n_36),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_25),
.B(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_25),
.A2(n_31),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_26),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AOI32xp33_ASAP7_75t_L g192 ( 
.A1(n_26),
.A2(n_45),
.A3(n_182),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_27),
.A2(n_29),
.A3(n_35),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_27),
.B(n_50),
.Y(n_194)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_32),
.B(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_35),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_43),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_45),
.B1(n_69),
.B2(n_70),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_44),
.A2(n_69),
.B(n_164),
.Y(n_227)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_47),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_47),
.A2(n_48),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_50),
.Y(n_193)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_78),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_61),
.A2(n_62),
.B1(n_92),
.B2(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_61),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_61),
.A2(n_62),
.B1(n_111),
.B2(n_241),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_62),
.B(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_143),
.B(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_62),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_62),
.A2(n_145),
.B(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_66),
.A2(n_117),
.B(n_120),
.Y(n_116)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_67),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_67),
.A2(n_68),
.B1(n_118),
.B2(n_255),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_68),
.B(n_96),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_76),
.B(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_76),
.A2(n_95),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_88),
.B(n_93),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_93),
.B1(n_94),
.B2(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_82),
.A2(n_89),
.B1(n_90),
.B2(n_102),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_83),
.A2(n_85),
.B1(n_87),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_83),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_83),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_83),
.B(n_151),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_83),
.A2(n_191),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_83),
.A2(n_85),
.B1(n_109),
.B2(n_259),
.Y(n_258)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_84),
.A2(n_156),
.B(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_86),
.B(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_86),
.A2(n_167),
.B(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_SL g210 ( 
.A(n_86),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_86),
.A2(n_157),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_101),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_105),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_104),
.Y(n_287)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_105),
.B(n_287),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_112),
.C(n_116),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_106),
.A2(n_107),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_108),
.B(n_110),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_112),
.B(n_116),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_113),
.A2(n_251),
.B(n_252),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_114),
.A2(n_115),
.B(n_202),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_115),
.B(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_115),
.A2(n_201),
.B(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_120),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI321xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_279),
.A3(n_288),
.B1(n_293),
.B2(n_298),
.C(n_300),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_243),
.C(n_275),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_217),
.B(n_242),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_196),
.B(n_216),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_177),
.B(n_195),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_152),
.B(n_176),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_130),
.B(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_134),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_135),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_136),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_147),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_142),
.C(n_147),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_148),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_161),
.B(n_175),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_154),
.B(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_168),
.B(n_174),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_165),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_188),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_184),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_192),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_192),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_211),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_212),
.C(n_213),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_205),
.C(n_208),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_201),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_208),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_219),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_221),
.B(n_222),
.C(n_230),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_225),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_236),
.C(n_239),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_244),
.A2(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_262),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_245),
.B(n_262),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_257),
.C(n_261),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_249),
.C(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_256),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_271),
.C(n_274),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_268),
.C(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_277),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_289),
.A2(n_294),
.B(n_297),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);


endmodule