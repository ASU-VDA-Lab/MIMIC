module fake_netlist_1_8546_n_908 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_908);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_908;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_384;
wire n_476;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_624;
wire n_255;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_565;
wire n_207;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_212;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g108 ( .A(n_44), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_3), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_41), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_58), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_107), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_65), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_56), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_48), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_75), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_29), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_1), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_91), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_5), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_43), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_14), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_11), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_31), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_55), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_84), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_18), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_86), .Y(n_130) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_16), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_92), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_0), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_42), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_64), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_76), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_12), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_95), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_71), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_0), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_6), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_8), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_50), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_24), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_106), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_94), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_54), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_32), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_17), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_37), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_82), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
INVx5_ASAP7_75t_L g153 ( .A(n_115), .Y(n_153) );
NOR2x1_ASAP7_75t_L g154 ( .A(n_113), .B(n_1), .Y(n_154) );
BUFx12f_ASAP7_75t_L g155 ( .A(n_110), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_109), .B(n_2), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_115), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_131), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_113), .Y(n_159) );
INVx5_ASAP7_75t_L g160 ( .A(n_121), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_117), .Y(n_161) );
INVx5_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_111), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
INVx5_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
BUFx12f_ASAP7_75t_L g171 ( .A(n_114), .Y(n_171) );
INVx5_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_109), .B(n_2), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_164), .B(n_118), .Y(n_175) );
AO22x2_ASAP7_75t_L g176 ( .A1(n_173), .A2(n_151), .B1(n_150), .B2(n_147), .Y(n_176) );
AO22x2_ASAP7_75t_L g177 ( .A1(n_173), .A2(n_151), .B1(n_150), .B2(n_147), .Y(n_177) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_173), .B(n_118), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_173), .A2(n_112), .B1(n_148), .B2(n_140), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_164), .B(n_122), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_159), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_164), .A2(n_141), .B1(n_137), .B2(n_144), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
INVxp67_ASAP7_75t_SL g186 ( .A(n_161), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g187 ( .A1(n_158), .A2(n_129), .B1(n_119), .B2(n_149), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_164), .A2(n_125), .B1(n_142), .B2(n_124), .Y(n_188) );
OAI22xp33_ASAP7_75t_L g189 ( .A1(n_158), .A2(n_129), .B1(n_119), .B2(n_126), .Y(n_189) );
OAI22xp33_ASAP7_75t_L g190 ( .A1(n_164), .A2(n_133), .B1(n_108), .B2(n_139), .Y(n_190) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_164), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_164), .A2(n_174), .B1(n_165), .B2(n_156), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_164), .B(n_108), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_164), .B(n_116), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_164), .B(n_120), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_159), .Y(n_201) );
NAND2xp33_ASAP7_75t_SL g202 ( .A(n_165), .B(n_123), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_166), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_164), .B(n_127), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_156), .B(n_3), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_166), .Y(n_207) );
OAI22xp33_ASAP7_75t_L g208 ( .A1(n_156), .A2(n_146), .B1(n_143), .B2(n_138), .Y(n_208) );
OAI22xp33_ASAP7_75t_SL g209 ( .A1(n_165), .A2(n_134), .B1(n_132), .B2(n_130), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_174), .B(n_128), .Y(n_210) );
OAI22xp33_ASAP7_75t_L g211 ( .A1(n_174), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_166), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_170), .A2(n_4), .B1(n_7), .B2(n_8), .Y(n_213) );
INVx1_ASAP7_75t_SL g214 ( .A(n_155), .Y(n_214) );
AO22x2_ASAP7_75t_L g215 ( .A1(n_170), .A2(n_152), .B1(n_157), .B2(n_161), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_161), .B(n_7), .Y(n_216) );
OR2x6_ASAP7_75t_L g217 ( .A(n_154), .B(n_9), .Y(n_217) );
OR2x6_ASAP7_75t_L g218 ( .A(n_154), .B(n_9), .Y(n_218) );
OAI22xp33_ASAP7_75t_SL g219 ( .A1(n_170), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_161), .B(n_10), .Y(n_220) );
AO22x2_ASAP7_75t_L g221 ( .A1(n_170), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_210), .B(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_215), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_193), .B(n_154), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_178), .B(n_161), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_179), .Y(n_226) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_186), .A2(n_152), .B(n_157), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_178), .B(n_161), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_215), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_215), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_206), .B(n_155), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_215), .Y(n_232) );
INVx1_ASAP7_75t_SL g233 ( .A(n_206), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_178), .B(n_163), .Y(n_234) );
XOR2xp5_ASAP7_75t_L g235 ( .A(n_179), .B(n_13), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_214), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_216), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_210), .B(n_155), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_184), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_216), .Y(n_240) );
INVxp67_ASAP7_75t_L g241 ( .A(n_176), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_184), .Y(n_242) );
INVx3_ASAP7_75t_R g243 ( .A(n_199), .Y(n_243) );
INVxp67_ASAP7_75t_SL g244 ( .A(n_220), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_208), .B(n_167), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_193), .B(n_167), .Y(n_246) );
XOR2xp5_ASAP7_75t_L g247 ( .A(n_187), .B(n_15), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_220), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_189), .B(n_163), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_194), .B(n_167), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_185), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_185), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_199), .B(n_167), .Y(n_253) );
AND2x2_ASAP7_75t_SL g254 ( .A(n_199), .B(n_152), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_185), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_194), .B(n_171), .Y(n_256) );
OR2x2_ASAP7_75t_SL g257 ( .A(n_221), .B(n_171), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_175), .Y(n_258) );
XOR2xp5_ASAP7_75t_L g259 ( .A(n_176), .B(n_16), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_175), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_176), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_176), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_177), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_199), .B(n_171), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_177), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_188), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_177), .B(n_163), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_197), .B(n_171), .Y(n_268) );
AO21x1_ASAP7_75t_L g269 ( .A1(n_219), .A2(n_209), .B(n_211), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_183), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_177), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_217), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_217), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_183), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_181), .B(n_169), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_197), .B(n_160), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_217), .B(n_152), .Y(n_277) );
INVxp33_ASAP7_75t_L g278 ( .A(n_188), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_217), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_183), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_192), .Y(n_281) );
NAND2xp33_ASAP7_75t_L g282 ( .A(n_191), .B(n_205), .Y(n_282) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_205), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_277), .A2(n_196), .B(n_200), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_233), .B(n_217), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_229), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_229), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_230), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_230), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_225), .B(n_218), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_257), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_225), .B(n_218), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_238), .B(n_209), .Y(n_293) );
INVx3_ASAP7_75t_L g294 ( .A(n_251), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_251), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_252), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_259), .Y(n_297) );
BUFx3_ASAP7_75t_L g298 ( .A(n_257), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_244), .Y(n_299) );
INVxp33_ASAP7_75t_L g300 ( .A(n_222), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_228), .B(n_218), .Y(n_301) );
INVx4_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_228), .B(n_218), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_252), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_255), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_278), .B(n_218), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_234), .B(n_213), .Y(n_307) );
BUFx10_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
INVx3_ASAP7_75t_SL g309 ( .A(n_271), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_234), .B(n_213), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_223), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_259), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_254), .B(n_213), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_262), .B(n_153), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_277), .A2(n_195), .B(n_182), .Y(n_316) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_262), .B(n_153), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_254), .B(n_213), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_224), .B(n_190), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_224), .B(n_221), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_224), .B(n_221), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_270), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_265), .B(n_153), .Y(n_323) );
BUFx12f_ASAP7_75t_SL g324 ( .A(n_231), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_231), .B(n_221), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_270), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_231), .B(n_157), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_274), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_223), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_241), .B(n_157), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_232), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_232), .Y(n_332) );
BUFx3_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
INVx5_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_302), .B(n_272), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_322), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_292), .B(n_237), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_322), .Y(n_339) );
INVx11_ASAP7_75t_L g340 ( .A(n_324), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_302), .B(n_272), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_299), .B(n_237), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_299), .B(n_240), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_302), .B(n_273), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_333), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_292), .B(n_240), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g347 ( .A(n_333), .B(n_273), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_292), .B(n_248), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_309), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
OR2x6_ASAP7_75t_L g352 ( .A(n_302), .B(n_261), .Y(n_352) );
NAND2x1_ASAP7_75t_SL g353 ( .A(n_325), .B(n_263), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_322), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_299), .B(n_248), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_292), .B(n_267), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_302), .B(n_279), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_285), .B(n_224), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_285), .B(n_224), .Y(n_359) );
NAND2x1p5_ASAP7_75t_L g360 ( .A(n_333), .B(n_279), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_285), .B(n_224), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_300), .B(n_239), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_322), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g364 ( .A(n_325), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_315), .Y(n_366) );
BUFx8_ASAP7_75t_SL g367 ( .A(n_348), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_352), .B(n_291), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_340), .Y(n_371) );
BUFx12f_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_335), .B(n_291), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_337), .Y(n_377) );
AND2x6_ASAP7_75t_L g378 ( .A(n_345), .B(n_291), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_335), .Y(n_379) );
INVx3_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_352), .Y(n_381) );
INVxp67_ASAP7_75t_SL g382 ( .A(n_337), .Y(n_382) );
INVx3_ASAP7_75t_SL g383 ( .A(n_335), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_335), .B(n_291), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_345), .Y(n_385) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_352), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_339), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_339), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_345), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_339), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_339), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
INVx6_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_345), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_375), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_388), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_373), .B(n_362), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_375), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_388), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_375), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g402 ( .A(n_368), .B(n_302), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_372), .A2(n_297), .B1(n_312), .B2(n_298), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_388), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_372), .A2(n_297), .B1(n_312), .B2(n_298), .Y(n_405) );
INVx4_ASAP7_75t_SL g406 ( .A(n_383), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_297), .Y(n_407) );
INVx5_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_372), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_372), .A2(n_297), .B1(n_312), .B2(n_298), .Y(n_410) );
AOI22xp33_ASAP7_75t_SL g411 ( .A1(n_368), .A2(n_312), .B1(n_298), .B2(n_291), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_368), .A2(n_298), .B1(n_325), .B2(n_302), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_378), .A2(n_306), .B1(n_269), .B2(n_325), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_368), .A2(n_325), .B1(n_364), .B2(n_318), .Y(n_414) );
BUFx2_ASAP7_75t_SL g415 ( .A(n_368), .Y(n_415) );
BUFx2_ASAP7_75t_SL g416 ( .A(n_369), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_378), .A2(n_306), .B1(n_269), .B2(n_235), .Y(n_419) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_383), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_378), .A2(n_306), .B1(n_235), .B2(n_362), .Y(n_421) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_382), .A2(n_321), .B1(n_320), .B2(n_318), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_367), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_369), .Y(n_424) );
OAI21xp5_ASAP7_75t_L g425 ( .A1(n_382), .A2(n_300), .B(n_293), .Y(n_425) );
OAI22xp5_ASAP7_75t_SL g426 ( .A1(n_371), .A2(n_247), .B1(n_226), .B2(n_242), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_378), .A2(n_318), .B1(n_314), .B2(n_285), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_383), .A2(n_364), .B1(n_320), .B2(n_321), .Y(n_428) );
INVx5_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
INVx6_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_383), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_382), .A2(n_320), .B1(n_321), .B2(n_318), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_383), .A2(n_236), .B1(n_300), .B2(n_290), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_378), .A2(n_236), .B1(n_247), .B2(n_239), .Y(n_434) );
INVx6_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_387), .A2(n_314), .B1(n_318), .B2(n_309), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_377), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_378), .A2(n_314), .B1(n_285), .B2(n_358), .Y(n_438) );
CKINVDCx6p67_ASAP7_75t_R g439 ( .A(n_383), .Y(n_439) );
BUFx4f_ASAP7_75t_SL g440 ( .A(n_423), .Y(n_440) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_434), .A2(n_384), .B(n_314), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_439), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
BUFx4f_ASAP7_75t_L g444 ( .A(n_439), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g445 ( .A1(n_420), .A2(n_378), .B1(n_369), .B2(n_376), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_417), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_419), .A2(n_324), .B1(n_370), .B2(n_378), .Y(n_448) );
AOI211xp5_ASAP7_75t_L g449 ( .A1(n_426), .A2(n_219), .B(n_293), .C(n_245), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_408), .Y(n_451) );
OAI222xp33_ASAP7_75t_L g452 ( .A1(n_419), .A2(n_370), .B1(n_384), .B2(n_376), .C1(n_380), .C2(n_374), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_421), .A2(n_324), .B1(n_370), .B2(n_378), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_421), .A2(n_408), .B1(n_403), .B2(n_405), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_396), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_413), .A2(n_414), .B1(n_407), .B2(n_324), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_437), .Y(n_457) );
INVx11_ASAP7_75t_L g458 ( .A(n_408), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_433), .A2(n_293), .B1(n_266), .B2(n_292), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_413), .A2(n_324), .B1(n_370), .B2(n_378), .Y(n_460) );
AOI22xp33_ASAP7_75t_SL g461 ( .A1(n_408), .A2(n_378), .B1(n_376), .B2(n_374), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_415), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_399), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_398), .B(n_266), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_411), .A2(n_370), .B1(n_378), .B2(n_224), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_399), .B(n_387), .Y(n_466) );
AOI22xp33_ASAP7_75t_SL g467 ( .A1(n_416), .A2(n_378), .B1(n_376), .B2(n_374), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_405), .A2(n_370), .B1(n_378), .B2(n_314), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_410), .A2(n_370), .B1(n_378), .B2(n_359), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_397), .Y(n_470) );
BUFx12f_ASAP7_75t_L g471 ( .A(n_429), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_401), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_401), .B(n_387), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_410), .A2(n_370), .B1(n_384), .B2(n_309), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_429), .B(n_374), .Y(n_475) );
CKINVDCx14_ASAP7_75t_R g476 ( .A(n_430), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g477 ( .A1(n_425), .A2(n_249), .B(n_353), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_400), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g479 ( .A1(n_412), .A2(n_384), .B(n_379), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_436), .A2(n_370), .B1(n_361), .B2(n_359), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_402), .A2(n_390), .B(n_377), .Y(n_481) );
AOI221xp5_ASAP7_75t_SL g482 ( .A1(n_427), .A2(n_249), .B1(n_327), .B2(n_307), .C(n_310), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_438), .A2(n_370), .B1(n_358), .B2(n_361), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_429), .B(n_168), .C(n_166), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_438), .A2(n_307), .B1(n_310), .B2(n_386), .Y(n_485) );
OAI21xp5_ASAP7_75t_SL g486 ( .A1(n_402), .A2(n_384), .B(n_379), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_427), .A2(n_307), .B1(n_310), .B2(n_386), .Y(n_487) );
BUFx3_ASAP7_75t_L g488 ( .A(n_431), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_404), .Y(n_489) );
BUFx3_ASAP7_75t_L g490 ( .A(n_431), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_429), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_429), .A2(n_384), .B1(n_309), .B2(n_379), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_430), .A2(n_376), .B1(n_374), .B2(n_380), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_406), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_430), .Y(n_495) );
BUFx2_ASAP7_75t_L g496 ( .A(n_431), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_422), .A2(n_307), .B1(n_310), .B2(n_386), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_424), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_424), .B(n_375), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_432), .B(n_390), .Y(n_500) );
OAI21xp5_ASAP7_75t_SL g501 ( .A1(n_431), .A2(n_379), .B(n_374), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_428), .A2(n_379), .B1(n_380), .B2(n_386), .Y(n_502) );
OAI21xp5_ASAP7_75t_SL g503 ( .A1(n_406), .A2(n_380), .B(n_379), .Y(n_503) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_435), .A2(n_379), .B1(n_380), .B2(n_386), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_435), .A2(n_307), .B1(n_310), .B2(n_386), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_406), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g507 ( .A1(n_435), .A2(n_353), .B(n_327), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_396), .Y(n_508) );
BUFx3_ASAP7_75t_L g509 ( .A(n_408), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_419), .A2(n_391), .B(n_390), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_417), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_421), .A2(n_309), .B1(n_380), .B2(n_340), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_448), .A2(n_381), .B1(n_392), .B2(n_386), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_466), .B(n_381), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_470), .B(n_391), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g516 ( .A1(n_464), .A2(n_327), .B1(n_303), .B2(n_301), .C1(n_338), .C2(n_349), .Y(n_516) );
OAI22xp33_ASAP7_75t_L g517 ( .A1(n_444), .A2(n_380), .B1(n_381), .B2(n_386), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_489), .B(n_391), .Y(n_518) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_451), .A2(n_376), .B1(n_386), .B2(n_392), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_444), .A2(n_376), .B1(n_381), .B2(n_392), .Y(n_520) );
AOI222xp33_ASAP7_75t_L g521 ( .A1(n_454), .A2(n_327), .B1(n_303), .B2(n_301), .C1(n_346), .C2(n_338), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_444), .A2(n_381), .B1(n_392), .B2(n_386), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_460), .A2(n_381), .B1(n_392), .B2(n_386), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g524 ( .A(n_449), .B(n_168), .C(n_166), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_453), .A2(n_392), .B1(n_381), .B2(n_376), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_456), .A2(n_381), .B1(n_392), .B2(n_393), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_446), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_511), .B(n_375), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_466), .B(n_381), .Y(n_529) );
OAI22x1_ASAP7_75t_L g530 ( .A1(n_462), .A2(n_394), .B1(n_309), .B2(n_350), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_451), .A2(n_392), .B1(n_381), .B2(n_393), .Y(n_531) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_462), .A2(n_392), .B1(n_381), .B2(n_393), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_482), .A2(n_303), .B1(n_301), .B2(n_356), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_469), .A2(n_392), .B1(n_393), .B2(n_348), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_465), .A2(n_392), .B1(n_393), .B2(n_348), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_445), .A2(n_461), .B1(n_467), .B2(n_442), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_442), .A2(n_393), .B1(n_385), .B2(n_371), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_468), .A2(n_393), .B1(n_348), .B2(n_366), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_477), .A2(n_393), .B1(n_348), .B2(n_366), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_497), .A2(n_393), .B1(n_348), .B2(n_366), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_473), .B(n_455), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_450), .B(n_327), .C(n_202), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_447), .B(n_394), .Y(n_543) );
OAI222xp33_ASAP7_75t_L g544 ( .A1(n_506), .A2(n_476), .B1(n_493), .B2(n_474), .C1(n_475), .C2(n_491), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_441), .A2(n_303), .B1(n_301), .B2(n_356), .Y(n_545) );
AOI222xp33_ASAP7_75t_L g546 ( .A1(n_452), .A2(n_301), .B1(n_303), .B2(n_338), .C1(n_346), .C2(n_349), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_480), .A2(n_348), .B1(n_366), .B2(n_367), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_476), .A2(n_385), .B1(n_350), .B2(n_394), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_512), .A2(n_366), .B1(n_356), .B2(n_352), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_485), .A2(n_366), .B1(n_352), .B2(n_341), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_483), .A2(n_366), .B1(n_352), .B2(n_341), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_471), .A2(n_385), .B1(n_394), .B2(n_395), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_487), .A2(n_366), .B1(n_341), .B2(n_336), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_447), .B(n_351), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_457), .B(n_351), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_505), .A2(n_336), .B1(n_357), .B2(n_344), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_459), .A2(n_346), .B1(n_349), .B2(n_319), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_457), .B(n_354), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_479), .A2(n_389), .B1(n_385), .B2(n_395), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_473), .B(n_354), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_478), .B(n_354), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_507), .A2(n_344), .B1(n_341), .B2(n_336), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_486), .A2(n_267), .B(n_290), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_455), .B(n_363), .Y(n_565) );
OAI222xp33_ASAP7_75t_L g566 ( .A1(n_475), .A2(n_389), .B1(n_395), .B2(n_385), .C1(n_290), .C2(n_342), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_498), .A2(n_344), .B1(n_336), .B2(n_357), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g568 ( .A1(n_501), .A2(n_319), .B1(n_355), .B2(n_343), .C(n_342), .Y(n_568) );
AOI222xp33_ASAP7_75t_L g569 ( .A1(n_440), .A2(n_319), .B1(n_166), .B2(n_168), .C1(n_343), .C2(n_355), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_363), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_498), .A2(n_344), .B1(n_336), .B2(n_341), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_471), .A2(n_344), .B1(n_357), .B2(n_389), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_499), .B(n_363), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_510), .A2(n_357), .B1(n_389), .B2(n_395), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_500), .A2(n_357), .B1(n_395), .B2(n_345), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_463), .B(n_363), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_509), .A2(n_395), .B1(n_333), .B2(n_166), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_494), .A2(n_395), .B1(n_333), .B2(n_166), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_478), .B(n_463), .Y(n_579) );
AOI222xp33_ASAP7_75t_L g580 ( .A1(n_503), .A2(n_166), .B1(n_168), .B2(n_157), .C1(n_330), .C2(n_160), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_502), .A2(n_333), .B1(n_168), .B2(n_166), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_472), .B(n_365), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_492), .A2(n_365), .B1(n_360), .B2(n_347), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_481), .A2(n_168), .B1(n_330), .B2(n_365), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_504), .A2(n_365), .B1(n_308), .B2(n_246), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_472), .A2(n_308), .B1(n_347), .B2(n_360), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_488), .A2(n_168), .B1(n_330), .B2(n_311), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_488), .A2(n_168), .B1(n_330), .B2(n_311), .Y(n_588) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_495), .A2(n_253), .B1(n_264), .B2(n_260), .C(n_258), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_496), .B(n_347), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_475), .A2(n_308), .B1(n_347), .B2(n_360), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_458), .A2(n_340), .B1(n_360), .B2(n_311), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_490), .A2(n_496), .B1(n_484), .B2(n_443), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_490), .A2(n_168), .B1(n_330), .B2(n_331), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_443), .B(n_168), .Y(n_595) );
OAI221xp5_ASAP7_75t_SL g596 ( .A1(n_508), .A2(n_258), .B1(n_260), .B2(n_250), .C(n_256), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g597 ( .A1(n_458), .A2(n_331), .B1(n_311), .B2(n_329), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_508), .A2(n_331), .B1(n_311), .B2(n_329), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_444), .A2(n_311), .B1(n_331), .B2(n_332), .Y(n_599) );
AOI221x1_ASAP7_75t_SL g600 ( .A1(n_449), .A2(n_17), .B1(n_18), .B2(n_19), .C(n_20), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_466), .B(n_160), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_444), .A2(n_331), .B1(n_332), .B2(n_295), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_444), .A2(n_331), .B1(n_332), .B2(n_295), .Y(n_603) );
AOI222xp33_ASAP7_75t_L g604 ( .A1(n_464), .A2(n_160), .B1(n_162), .B2(n_282), .C1(n_315), .C2(n_323), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_444), .A2(n_295), .B1(n_296), .B2(n_305), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_448), .A2(n_329), .B1(n_323), .B2(n_315), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_451), .A2(n_308), .B1(n_334), .B2(n_329), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_448), .A2(n_329), .B1(n_323), .B2(n_315), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g609 ( .A1(n_451), .A2(n_308), .B1(n_334), .B2(n_323), .Y(n_609) );
OA21x2_ASAP7_75t_L g610 ( .A1(n_510), .A2(n_227), .B(n_287), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_448), .A2(n_323), .B1(n_315), .B2(n_287), .Y(n_611) );
AOI221xp5_ASAP7_75t_SL g612 ( .A1(n_449), .A2(n_19), .B1(n_20), .B2(n_21), .C(n_22), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_600), .B(n_268), .C(n_276), .D(n_23), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_514), .B(n_21), .Y(n_614) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_564), .A2(n_334), .B1(n_287), .B2(n_288), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_541), .B(n_22), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_612), .A2(n_160), .B(n_162), .Y(n_617) );
OA211x2_ASAP7_75t_L g618 ( .A1(n_557), .A2(n_23), .B(n_24), .C(n_25), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_527), .B(n_25), .Y(n_619) );
AOI21xp5_ASAP7_75t_SL g620 ( .A1(n_536), .A2(n_323), .B(n_315), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_514), .B(n_26), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_527), .B(n_26), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_519), .A2(n_305), .B1(n_295), .B2(n_296), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_541), .B(n_27), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_524), .B(n_162), .C(n_160), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_565), .B(n_27), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_529), .B(n_28), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_593), .B(n_162), .C(n_160), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_565), .B(n_29), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_521), .A2(n_289), .B1(n_287), .B2(n_288), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_561), .B(n_30), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_561), .B(n_30), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_529), .B(n_31), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_517), .B(n_153), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_570), .B(n_32), .Y(n_635) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_542), .B(n_160), .C(n_162), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_570), .B(n_33), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_573), .B(n_33), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_573), .B(n_34), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_579), .B(n_34), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_576), .B(n_160), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_576), .B(n_160), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_515), .B(n_162), .Y(n_643) );
NAND4xp25_ASAP7_75t_L g644 ( .A(n_569), .B(n_284), .C(n_316), .D(n_323), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_546), .B(n_284), .C(n_316), .D(n_323), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_518), .B(n_162), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_601), .B(n_162), .Y(n_647) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_544), .A2(n_317), .B(n_315), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_580), .B(n_162), .C(n_153), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_601), .B(n_162), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_543), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_548), .B(n_162), .C(n_153), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_532), .B(n_153), .C(n_169), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_523), .B(n_590), .C(n_526), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_554), .B(n_555), .Y(n_655) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_590), .B(n_153), .C(n_169), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_528), .B(n_169), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_568), .B(n_35), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_531), .B(n_36), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_513), .B(n_38), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_583), .A2(n_313), .B(n_305), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_574), .B(n_169), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_575), .B(n_169), .Y(n_663) );
OA21x2_ASAP7_75t_L g664 ( .A1(n_539), .A2(n_525), .B(n_534), .Y(n_664) );
OA21x2_ASAP7_75t_L g665 ( .A1(n_566), .A2(n_288), .B(n_289), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_595), .B(n_153), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_559), .B(n_169), .Y(n_667) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_545), .B(n_284), .C(n_316), .D(n_275), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_552), .A2(n_317), .B(n_212), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_562), .B(n_169), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_595), .B(n_153), .Y(n_671) );
NAND4xp25_ASAP7_75t_SL g672 ( .A(n_545), .B(n_288), .C(n_289), .D(n_313), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_582), .B(n_169), .Y(n_673) );
OA21x2_ASAP7_75t_L g674 ( .A1(n_520), .A2(n_289), .B(n_212), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_586), .B(n_295), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_558), .B(n_169), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_558), .B(n_169), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_572), .A2(n_296), .B1(n_313), .B2(n_305), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_610), .B(n_172), .Y(n_679) );
OAI22xp33_ASAP7_75t_SL g680 ( .A1(n_596), .A2(n_317), .B1(n_153), .B2(n_172), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_610), .B(n_172), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_586), .B(n_39), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_549), .B(n_40), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_551), .B(n_45), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_535), .B(n_172), .C(n_313), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_567), .B(n_46), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_537), .A2(n_313), .B1(n_305), .B2(n_296), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_547), .B(n_172), .C(n_296), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_610), .B(n_172), .Y(n_689) );
OAI21xp5_ASAP7_75t_SL g690 ( .A1(n_560), .A2(n_317), .B(n_286), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_610), .B(n_172), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_563), .B(n_172), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_571), .B(n_47), .Y(n_693) );
NAND4xp25_ASAP7_75t_L g694 ( .A(n_550), .B(n_195), .C(n_196), .D(n_200), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_591), .A2(n_317), .B1(n_286), .B2(n_328), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_589), .B(n_286), .C(n_304), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_585), .B(n_49), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_591), .A2(n_317), .B1(n_286), .B2(n_328), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_522), .A2(n_172), .B1(n_283), .B2(n_182), .C(n_192), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_540), .B(n_172), .Y(n_700) );
AOI21xp5_ASAP7_75t_SL g701 ( .A1(n_530), .A2(n_317), .B(n_308), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_585), .B(n_172), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_538), .B(n_286), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_581), .B(n_51), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_556), .B(n_52), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_553), .A2(n_212), .B1(n_192), .B2(n_204), .C(n_207), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_605), .B(n_286), .C(n_204), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_584), .B(n_286), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_604), .B(n_207), .C(n_204), .D(n_180), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_533), .B(n_286), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_533), .A2(n_304), .B1(n_294), .B2(n_328), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_516), .B(n_328), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_609), .B(n_53), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_592), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_602), .B(n_326), .Y(n_715) );
NAND3xp33_ASAP7_75t_L g716 ( .A(n_654), .B(n_607), .C(n_578), .Y(n_716) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_648), .B(n_603), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_624), .B(n_599), .Y(n_718) );
NOR3xp33_ASAP7_75t_SL g719 ( .A(n_644), .B(n_597), .C(n_611), .Y(n_719) );
BUFx3_ASAP7_75t_L g720 ( .A(n_614), .Y(n_720) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_614), .Y(n_721) );
XOR2x2_ASAP7_75t_L g722 ( .A(n_616), .B(n_608), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_714), .B(n_606), .Y(n_723) );
AND2x2_ASAP7_75t_SL g724 ( .A(n_621), .B(n_577), .Y(n_724) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_620), .A2(n_594), .B(n_588), .C(n_587), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_651), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_655), .B(n_57), .Y(n_727) );
NAND3xp33_ASAP7_75t_SL g728 ( .A(n_696), .B(n_598), .C(n_326), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_621), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_620), .B(n_207), .C(n_326), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_628), .B(n_326), .C(n_203), .Y(n_731) );
AO21x2_ASAP7_75t_L g732 ( .A1(n_619), .A2(n_203), .B(n_198), .Y(n_732) );
AOI211x1_ASAP7_75t_L g733 ( .A1(n_615), .A2(n_59), .B(n_60), .C(n_61), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_627), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_627), .B(n_62), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_622), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_633), .Y(n_737) );
NAND4xp75_ASAP7_75t_L g738 ( .A(n_618), .B(n_243), .C(n_63), .D(n_66), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_658), .B(n_201), .C(n_198), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_635), .B(n_67), .Y(n_740) );
AO21x2_ASAP7_75t_L g741 ( .A1(n_626), .A2(n_201), .B(n_180), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_640), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_645), .A2(n_308), .B1(n_304), .B2(n_294), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_629), .Y(n_744) );
OAI211xp5_ASAP7_75t_SL g745 ( .A1(n_615), .A2(n_304), .B(n_294), .C(n_70), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_637), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_638), .B(n_68), .Y(n_747) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_658), .B(n_304), .C(n_294), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_639), .B(n_69), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_664), .B(n_642), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_675), .B(n_631), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g752 ( .A1(n_696), .A2(n_304), .B1(n_294), .B2(n_308), .C(n_78), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_632), .B(n_72), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_664), .B(n_73), .Y(n_754) );
NAND3xp33_ASAP7_75t_SL g755 ( .A(n_690), .B(n_74), .C(n_79), .Y(n_755) );
AND2x4_ASAP7_75t_L g756 ( .A(n_634), .B(n_80), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_664), .B(n_81), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_674), .Y(n_758) );
OAI21xp33_ASAP7_75t_SL g759 ( .A1(n_701), .A2(n_304), .B(n_294), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_647), .B(n_83), .Y(n_760) );
INVx1_ASAP7_75t_SL g761 ( .A(n_666), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_636), .B(n_85), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_701), .B(n_87), .Y(n_763) );
OAI21xp5_ASAP7_75t_L g764 ( .A1(n_652), .A2(n_294), .B(n_89), .Y(n_764) );
AOI22xp33_ASAP7_75t_SL g765 ( .A1(n_682), .A2(n_294), .B1(n_90), .B2(n_93), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_659), .B(n_88), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_697), .B(n_96), .Y(n_767) );
NAND4xp75_ASAP7_75t_L g768 ( .A(n_697), .B(n_97), .C(n_98), .D(n_99), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_672), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_769) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_649), .B(n_103), .C(n_104), .D(n_105), .Y(n_770) );
OAI21xp5_ASAP7_75t_L g771 ( .A1(n_680), .A2(n_280), .B(n_281), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_641), .Y(n_772) );
AO21x2_ASAP7_75t_L g773 ( .A1(n_679), .A2(n_280), .B(n_281), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g774 ( .A(n_656), .B(n_625), .C(n_653), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g775 ( .A1(n_665), .A2(n_623), .B1(n_713), .B2(n_705), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_665), .B(n_666), .Y(n_776) );
NAND4xp75_ASAP7_75t_L g777 ( .A(n_683), .B(n_684), .C(n_705), .D(n_660), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_681), .B(n_691), .Y(n_778) );
CKINVDCx8_ASAP7_75t_R g779 ( .A(n_669), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g780 ( .A(n_686), .B(n_693), .C(n_704), .D(n_650), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_688), .B(n_613), .C(n_685), .Y(n_781) );
INVx2_ASAP7_75t_SL g782 ( .A(n_671), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_643), .B(n_646), .C(n_617), .Y(n_783) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_694), .B(n_657), .C(n_702), .Y(n_784) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_689), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_711), .A2(n_712), .B1(n_687), .B2(n_630), .Y(n_786) );
NOR3xp33_ASAP7_75t_L g787 ( .A(n_667), .B(n_673), .C(n_670), .Y(n_787) );
OR2x2_ASAP7_75t_L g788 ( .A(n_715), .B(n_671), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_711), .A2(n_704), .B1(n_677), .B2(n_676), .Y(n_789) );
AOI22xp33_ASAP7_75t_SL g790 ( .A1(n_695), .A2(n_698), .B1(n_707), .B2(n_678), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_630), .A2(n_710), .B1(n_692), .B2(n_668), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_703), .B(n_699), .Y(n_792) );
XNOR2xp5_ASAP7_75t_L g793 ( .A(n_722), .B(n_662), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_750), .B(n_661), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_736), .B(n_708), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_726), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_721), .B(n_700), .Y(n_797) );
XOR2x2_ASAP7_75t_L g798 ( .A(n_717), .B(n_663), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_742), .Y(n_799) );
NAND3x1_ASAP7_75t_SL g800 ( .A(n_763), .B(n_709), .C(n_706), .Y(n_800) );
NAND4xp75_ASAP7_75t_SL g801 ( .A(n_776), .B(n_767), .C(n_718), .D(n_792), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_734), .Y(n_802) );
NAND4xp75_ASAP7_75t_L g803 ( .A(n_759), .B(n_733), .C(n_724), .D(n_754), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_720), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_729), .B(n_737), .Y(n_805) );
AND2x4_ASAP7_75t_L g806 ( .A(n_785), .B(n_761), .Y(n_806) );
XNOR2xp5_ASAP7_75t_L g807 ( .A(n_777), .B(n_780), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_744), .B(n_746), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_758), .Y(n_809) );
OR2x2_ASAP7_75t_L g810 ( .A(n_761), .B(n_778), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_772), .B(n_723), .Y(n_811) );
NOR4xp25_ASAP7_75t_L g812 ( .A(n_754), .B(n_757), .C(n_716), .D(n_728), .Y(n_812) );
XNOR2x2_ASAP7_75t_L g813 ( .A(n_755), .B(n_728), .Y(n_813) );
AND2x4_ASAP7_75t_SL g814 ( .A(n_782), .B(n_719), .Y(n_814) );
AOI22x1_ASAP7_75t_SL g815 ( .A1(n_770), .A2(n_775), .B1(n_755), .B2(n_779), .Y(n_815) );
NAND4xp75_ASAP7_75t_SL g816 ( .A(n_735), .B(n_762), .C(n_727), .D(n_740), .Y(n_816) );
INVx1_ASAP7_75t_SL g817 ( .A(n_747), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_778), .B(n_751), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_788), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_781), .A2(n_775), .B1(n_730), .B2(n_783), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_773), .B(n_787), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_732), .B(n_790), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_732), .B(n_790), .Y(n_823) );
NAND4xp75_ASAP7_75t_SL g824 ( .A(n_749), .B(n_760), .C(n_738), .D(n_768), .Y(n_824) );
XNOR2x2_ASAP7_75t_L g825 ( .A(n_752), .B(n_748), .Y(n_825) );
AND2x2_ASAP7_75t_L g826 ( .A(n_741), .B(n_784), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_789), .B(n_791), .Y(n_827) );
INVx4_ASAP7_75t_L g828 ( .A(n_756), .Y(n_828) );
AND2x2_ASAP7_75t_L g829 ( .A(n_786), .B(n_743), .Y(n_829) );
XOR2x2_ASAP7_75t_L g830 ( .A(n_752), .B(n_769), .Y(n_830) );
NAND4xp75_ASAP7_75t_L g831 ( .A(n_764), .B(n_771), .C(n_745), .D(n_765), .Y(n_831) );
NAND2xp5_ASAP7_75t_SL g832 ( .A(n_766), .B(n_739), .Y(n_832) );
XOR2xp5_ASAP7_75t_L g833 ( .A(n_753), .B(n_766), .Y(n_833) );
XOR2x2_ASAP7_75t_L g834 ( .A(n_807), .B(n_731), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_810), .Y(n_835) );
INVx1_ASAP7_75t_SL g836 ( .A(n_804), .Y(n_836) );
AND2x2_ASAP7_75t_L g837 ( .A(n_806), .B(n_774), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_810), .Y(n_838) );
AND2x2_ASAP7_75t_L g839 ( .A(n_806), .B(n_756), .Y(n_839) );
XNOR2xp5_ASAP7_75t_L g840 ( .A(n_807), .B(n_725), .Y(n_840) );
XOR2x2_ASAP7_75t_L g841 ( .A(n_801), .B(n_725), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_806), .B(n_818), .Y(n_842) );
XNOR2x2_ASAP7_75t_L g843 ( .A(n_813), .B(n_825), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_818), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_796), .Y(n_845) );
INVx2_ASAP7_75t_SL g846 ( .A(n_809), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_805), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_805), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_826), .B(n_821), .Y(n_849) );
XOR2x2_ASAP7_75t_L g850 ( .A(n_793), .B(n_798), .Y(n_850) );
XOR2x2_ASAP7_75t_L g851 ( .A(n_793), .B(n_798), .Y(n_851) );
INVx1_ASAP7_75t_SL g852 ( .A(n_817), .Y(n_852) );
INVx1_ASAP7_75t_SL g853 ( .A(n_814), .Y(n_853) );
INVxp67_ASAP7_75t_L g854 ( .A(n_826), .Y(n_854) );
XOR2x2_ASAP7_75t_L g855 ( .A(n_800), .B(n_816), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_819), .Y(n_856) );
INVx2_ASAP7_75t_SL g857 ( .A(n_809), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_820), .A2(n_827), .B1(n_830), .B2(n_814), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_802), .Y(n_859) );
XNOR2xp5_ASAP7_75t_L g860 ( .A(n_833), .B(n_800), .Y(n_860) );
XNOR2x1_ASAP7_75t_L g861 ( .A(n_827), .B(n_830), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_858), .A2(n_828), .B1(n_803), .B2(n_831), .Y(n_862) );
INVx2_ASAP7_75t_L g863 ( .A(n_846), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g864 ( .A(n_853), .Y(n_864) );
INVx3_ASAP7_75t_L g865 ( .A(n_843), .Y(n_865) );
INVx2_ASAP7_75t_SL g866 ( .A(n_836), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g867 ( .A1(n_861), .A2(n_828), .B1(n_803), .B2(n_831), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_846), .Y(n_868) );
XNOR2x1_ASAP7_75t_L g869 ( .A(n_843), .B(n_825), .Y(n_869) );
HB1xp67_ASAP7_75t_L g870 ( .A(n_835), .Y(n_870) );
AO22x2_ASAP7_75t_L g871 ( .A1(n_861), .A2(n_822), .B1(n_823), .B2(n_799), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_841), .A2(n_829), .B1(n_815), .B2(n_821), .Y(n_872) );
BUFx3_ASAP7_75t_L g873 ( .A(n_852), .Y(n_873) );
XOR2x2_ASAP7_75t_L g874 ( .A(n_850), .B(n_824), .Y(n_874) );
OA22x2_ASAP7_75t_L g875 ( .A1(n_840), .A2(n_828), .B1(n_829), .B2(n_808), .Y(n_875) );
OA22x2_ASAP7_75t_L g876 ( .A1(n_860), .A2(n_832), .B1(n_794), .B2(n_811), .Y(n_876) );
BUFx12f_ASAP7_75t_L g877 ( .A(n_864), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_873), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_870), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_870), .Y(n_880) );
INVx5_ASAP7_75t_SL g881 ( .A(n_869), .Y(n_881) );
AOI22x1_ASAP7_75t_L g882 ( .A1(n_865), .A2(n_871), .B1(n_875), .B2(n_874), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_866), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_865), .Y(n_884) );
AOI22x1_ASAP7_75t_L g885 ( .A1(n_884), .A2(n_871), .B1(n_854), .B2(n_875), .Y(n_885) );
OA22x2_ASAP7_75t_L g886 ( .A1(n_878), .A2(n_872), .B1(n_867), .B2(n_862), .Y(n_886) );
OAI222xp33_ASAP7_75t_L g887 ( .A1(n_882), .A2(n_876), .B1(n_867), .B2(n_862), .C1(n_854), .C2(n_849), .Y(n_887) );
NAND4xp75_ASAP7_75t_L g888 ( .A(n_881), .B(n_837), .C(n_855), .D(n_876), .Y(n_888) );
OAI222xp33_ASAP7_75t_L g889 ( .A1(n_883), .A2(n_871), .B1(n_868), .B2(n_863), .C1(n_841), .C2(n_839), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_886), .Y(n_890) );
NOR4xp25_ASAP7_75t_L g891 ( .A(n_887), .B(n_881), .C(n_880), .D(n_879), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_888), .A2(n_881), .B1(n_855), .B2(n_851), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_890), .Y(n_893) );
OAI21xp5_ASAP7_75t_L g894 ( .A1(n_891), .A2(n_886), .B(n_889), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_893), .Y(n_895) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_894), .Y(n_896) );
AND4x1_ASAP7_75t_L g897 ( .A(n_895), .B(n_892), .C(n_877), .D(n_812), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_896), .Y(n_898) );
INVx1_ASAP7_75t_SL g899 ( .A(n_898), .Y(n_899) );
OAI22xp5_ASAP7_75t_L g900 ( .A1(n_898), .A2(n_877), .B1(n_885), .B2(n_838), .Y(n_900) );
NOR4xp25_ASAP7_75t_L g901 ( .A(n_899), .B(n_897), .C(n_850), .D(n_851), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_901), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g903 ( .A1(n_902), .A2(n_900), .B1(n_834), .B2(n_842), .Y(n_903) );
INVxp67_ASAP7_75t_SL g904 ( .A(n_903), .Y(n_904) );
NAND4xp25_ASAP7_75t_L g905 ( .A(n_904), .B(n_844), .C(n_856), .D(n_834), .Y(n_905) );
INVx1_ASAP7_75t_SL g906 ( .A(n_905), .Y(n_906) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_906), .A2(n_848), .B1(n_847), .B2(n_845), .C(n_857), .Y(n_907) );
AOI211xp5_ASAP7_75t_L g908 ( .A1(n_907), .A2(n_859), .B(n_795), .C(n_797), .Y(n_908) );
endmodule