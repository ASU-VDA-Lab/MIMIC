module fake_jpeg_15672_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_64),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_0),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_51),
.B1(n_49),
.B2(n_44),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_0),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_52),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_80),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_51),
.B1(n_41),
.B2(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_41),
.B1(n_54),
.B2(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_50),
.B1(n_40),
.B2(n_57),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_47),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_2),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_67),
.Y(n_83)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_48),
.Y(n_85)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_95),
.CI(n_96),
.CON(n_106),
.SN(n_106)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_50),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_93),
.C(n_97),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_70),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_1),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_101),
.B1(n_102),
.B2(n_5),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_3),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OR2x2_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_4),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_74),
.B1(n_6),
.B2(n_7),
.Y(n_108)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_87),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_90),
.C(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_88),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_113),
.B(n_95),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_120),
.A2(n_122),
.B1(n_117),
.B2(n_113),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_117),
.A2(n_108),
.B1(n_84),
.B2(n_104),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_125),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_109),
.B1(n_107),
.B2(n_111),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_111),
.B1(n_103),
.B2(n_11),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_100),
.C(n_9),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_126),
.C(n_13),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_127),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_134),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_131),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_137),
.B(n_12),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_139)
);

OAI21x1_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_20),
.B(n_21),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_24),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_26),
.B(n_28),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_29),
.C(n_31),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_33),
.B(n_34),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_35),
.Y(n_145)
);


endmodule