module fake_jpeg_27942_n_46 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_4),
.B(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_5),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_5),
.B(n_2),
.Y(n_10)
);

OAI21xp33_ASAP7_75t_L g11 ( 
.A1(n_4),
.A2(n_3),
.B(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx24_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_17),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_3),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_18),
.A2(n_7),
.B1(n_9),
.B2(n_20),
.Y(n_27)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_2),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_23),
.Y(n_29)
);

AND2x6_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_12),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_10),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_14),
.C(n_13),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_32),
.C(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_16),
.B1(n_25),
.B2(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.C(n_36),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_19),
.C(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_16),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_26),
.C(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_24),
.C(n_36),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_35),
.B(n_33),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_33),
.B(n_40),
.C(n_44),
.Y(n_46)
);


endmodule