module fake_netlist_1_7629_n_10 (n_1, n_2, n_0, n_10);
input n_1;
input n_2;
input n_0;
output n_10;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_8;
NAND2xp5_ASAP7_75t_L g3 ( .A(n_2), .B(n_1), .Y(n_3) );
NAND2xp33_ASAP7_75t_SL g4 ( .A(n_0), .B(n_1), .Y(n_4) );
NAND2xp5_ASAP7_75t_L g5 ( .A(n_3), .B(n_0), .Y(n_5) );
INVx4_ASAP7_75t_L g6 ( .A(n_5), .Y(n_6) );
OAI222xp33_ASAP7_75t_L g7 ( .A1(n_6), .A2(n_0), .B1(n_1), .B2(n_2), .C1(n_4), .C2(n_5), .Y(n_7) );
OAI22xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_6), .B1(n_1), .B2(n_2), .Y(n_8) );
XNOR2xp5_ASAP7_75t_L g9 ( .A(n_8), .B(n_7), .Y(n_9) );
AOI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_0), .B1(n_2), .B2(n_6), .Y(n_10) );
endmodule