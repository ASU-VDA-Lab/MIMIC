module real_aes_16677_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_867, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_867;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_0), .Y(n_230) );
AND2x4_ASAP7_75t_L g108 ( .A(n_1), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g845 ( .A(n_2), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_3), .A2(n_5), .B1(n_177), .B2(n_580), .Y(n_579) );
AOI21xp33_ASAP7_75t_SL g849 ( .A1(n_4), .A2(n_850), .B(n_857), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_6), .A2(n_22), .B1(n_140), .B2(n_180), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_7), .A2(n_54), .B1(n_228), .B2(n_529), .Y(n_528) );
BUFx3_ASAP7_75t_L g171 ( .A(n_8), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_9), .A2(n_15), .B1(n_516), .B2(n_543), .Y(n_554) );
INVx1_ASAP7_75t_L g109 ( .A(n_10), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_11), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_12), .B(n_143), .Y(n_142) );
BUFx2_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
OR2x2_ASAP7_75t_L g834 ( .A(n_13), .B(n_32), .Y(n_834) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_14), .Y(n_141) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_16), .A2(n_83), .B1(n_822), .B2(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_16), .Y(n_823) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_17), .B(n_165), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_18), .B(n_190), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_19), .A2(n_84), .B1(n_140), .B2(n_165), .Y(n_239) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_20), .A2(n_49), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g864 ( .A(n_21), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_23), .B(n_180), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_24), .Y(n_652) );
INVx4_ASAP7_75t_R g568 ( .A(n_25), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_26), .B(n_145), .Y(n_601) );
AO32x2_ASAP7_75t_L g236 ( .A1(n_27), .A2(n_157), .A3(n_158), .B1(n_237), .B2(n_240), .Y(n_236) );
AO32x1_ASAP7_75t_L g274 ( .A1(n_27), .A2(n_157), .A3(n_158), .B1(n_237), .B2(n_240), .Y(n_274) );
INVx1_ASAP7_75t_L g582 ( .A(n_28), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_29), .B(n_180), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_SL g515 ( .A1(n_30), .A2(n_144), .B(n_516), .C(n_517), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_31), .A2(n_46), .B1(n_148), .B2(n_516), .Y(n_650) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_32), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_33), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_34), .A2(n_52), .B1(n_168), .B2(n_180), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_35), .A2(n_89), .B1(n_140), .B2(n_148), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_36), .B(n_147), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_37), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_37), .Y(n_848) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_38), .B(n_203), .Y(n_263) );
INVx1_ASAP7_75t_L g604 ( .A(n_39), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_40), .A2(n_67), .B1(n_148), .B2(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_41), .B(n_516), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_42), .Y(n_544) );
INVx2_ASAP7_75t_L g829 ( .A(n_43), .Y(n_829) );
INVx1_ASAP7_75t_L g111 ( .A(n_44), .Y(n_111) );
BUFx3_ASAP7_75t_L g832 ( .A(n_44), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_45), .B(n_265), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_47), .A2(n_85), .B1(n_148), .B2(n_516), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_48), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_50), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_51), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_53), .A2(n_77), .B1(n_202), .B2(n_203), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_55), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_56), .A2(n_81), .B1(n_140), .B2(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g136 ( .A(n_57), .Y(n_136) );
AND2x4_ASAP7_75t_L g154 ( .A(n_58), .B(n_155), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_59), .A2(n_90), .B1(n_148), .B2(n_578), .Y(n_577) );
AO22x1_ASAP7_75t_L g533 ( .A1(n_60), .A2(n_72), .B1(n_534), .B2(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_61), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g155 ( .A(n_62), .Y(n_155) );
AND2x2_ASAP7_75t_L g519 ( .A(n_63), .B(n_157), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_64), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_65), .A2(n_228), .B(n_229), .C(n_231), .Y(n_227) );
NAND3xp33_ASAP7_75t_L g152 ( .A(n_66), .B(n_140), .C(n_150), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_68), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_69), .B(n_228), .Y(n_548) );
AND2x2_ASAP7_75t_L g233 ( .A(n_70), .B(n_234), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_71), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_73), .B(n_180), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_74), .A2(n_94), .B1(n_165), .B2(n_202), .Y(n_206) );
INVx2_ASAP7_75t_L g145 ( .A(n_75), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_76), .B(n_184), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_78), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_79), .B(n_157), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_80), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_82), .B(n_134), .Y(n_531) );
INVx1_ASAP7_75t_L g822 ( .A(n_83), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_86), .B(n_150), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_87), .A2(n_100), .B1(n_148), .B2(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_88), .B(n_203), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_91), .B(n_157), .Y(n_540) );
INVx1_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_92), .B(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_93), .B(n_190), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_95), .A2(n_205), .B(n_228), .C(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g571 ( .A(n_96), .B(n_234), .Y(n_571) );
INVxp67_ASAP7_75t_SL g862 ( .A(n_97), .Y(n_862) );
NAND2xp33_ASAP7_75t_L g547 ( .A(n_98), .B(n_143), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_99), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_118), .B(n_863), .Y(n_101) );
CKINVDCx6p67_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g865 ( .A(n_104), .Y(n_865) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_114), .Y(n_105) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .C(n_112), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AND3x2_ASAP7_75t_L g841 ( .A(n_110), .B(n_112), .C(n_833), .Y(n_841) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g861 ( .A(n_111), .Y(n_861) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g497 ( .A(n_113), .Y(n_497) );
NOR2x1p5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AO21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_825), .B(n_835), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_820), .B1(n_821), .B2(n_824), .Y(n_119) );
INVxp33_ASAP7_75t_SL g824 ( .A(n_120), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_496), .B1(n_498), .B2(n_502), .Y(n_120) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_406), .Y(n_121) );
NAND4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_311), .C(n_338), .D(n_374), .Y(n_122) );
AOI221x1_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_216), .B1(n_250), .B2(n_286), .C(n_290), .Y(n_123) );
NAND3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_192), .C(n_214), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_159), .Y(n_127) );
INVx2_ASAP7_75t_L g251 ( .A(n_128), .Y(n_251) );
AND2x2_ASAP7_75t_L g424 ( .A(n_128), .B(n_368), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_128), .B(n_215), .Y(n_433) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g439 ( .A(n_129), .Y(n_439) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g284 ( .A(n_130), .Y(n_284) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g367 ( .A(n_131), .B(n_213), .Y(n_367) );
OAI21x1_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_137), .B(n_156), .Y(n_131) );
OAI21xp5_ASAP7_75t_L g296 ( .A1(n_132), .A2(n_137), .B(n_156), .Y(n_296) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AO31x2_ASAP7_75t_L g552 ( .A1(n_133), .A2(n_553), .A3(n_557), .B(n_558), .Y(n_552) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
INVx2_ASAP7_75t_L g211 ( .A(n_134), .Y(n_211) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_134), .A2(n_232), .B(n_531), .Y(n_537) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_135), .Y(n_158) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_146), .B(n_153), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_142), .B(n_144), .Y(n_138) );
INVx2_ASAP7_75t_SL g203 ( .A(n_140), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_140), .B(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_141), .Y(n_143) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
INVx1_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx1_ASAP7_75t_L g228 ( .A(n_141), .Y(n_228) );
INVx3_ASAP7_75t_L g516 ( .A(n_141), .Y(n_516) );
INVx1_ASAP7_75t_L g530 ( .A(n_141), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_143), .A2(n_168), .B1(n_568), .B2(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g578 ( .A(n_143), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g163 ( .A1(n_144), .A2(n_164), .B1(n_166), .B2(n_167), .Y(n_163) );
INVx6_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_144), .A2(n_181), .B1(n_238), .B2(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_144), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_144), .A2(n_547), .B(n_548), .Y(n_546) );
A2O1A1Ixp33_ASAP7_75t_L g590 ( .A1(n_144), .A2(n_527), .B(n_533), .C(n_537), .Y(n_590) );
BUFx8_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g151 ( .A(n_145), .Y(n_151) );
INVx2_ASAP7_75t_L g186 ( .A(n_145), .Y(n_186) );
INVx1_ASAP7_75t_L g205 ( .A(n_145), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B(n_152), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g580 ( .A(n_148), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_148), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_151), .B(n_604), .Y(n_603) );
AOI31xp67_ASAP7_75t_L g161 ( .A1(n_153), .A2(n_162), .A3(n_163), .B(n_169), .Y(n_161) );
OAI21x1_ASAP7_75t_L g174 ( .A1(n_153), .A2(n_175), .B(n_182), .Y(n_174) );
INVx1_ASAP7_75t_L g550 ( .A(n_153), .Y(n_550) );
AND2x2_ASAP7_75t_L g608 ( .A(n_153), .B(n_158), .Y(n_608) );
AO31x2_ASAP7_75t_L g647 ( .A1(n_153), .A2(n_162), .A3(n_648), .B(n_651), .Y(n_647) );
BUFx10_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
INVx1_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_154), .A2(n_199), .A3(n_243), .B(n_248), .Y(n_242) );
BUFx10_ASAP7_75t_L g557 ( .A(n_154), .Y(n_557) );
INVx2_ASAP7_75t_L g162 ( .A(n_157), .Y(n_162) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_157), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_158), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
BUFx3_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_158), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_SL g257 ( .A(n_158), .Y(n_257) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_159), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_159), .B(n_395), .Y(n_394) );
INVxp67_ASAP7_75t_L g437 ( .A(n_159), .Y(n_437) );
AND2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_172), .Y(n_159) );
AND2x2_ASAP7_75t_L g215 ( .A(n_160), .B(n_198), .Y(n_215) );
INVx2_ASAP7_75t_L g293 ( .A(n_160), .Y(n_293) );
AND2x2_ASAP7_75t_L g358 ( .A(n_160), .B(n_296), .Y(n_358) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g213 ( .A(n_161), .Y(n_213) );
INVx3_ASAP7_75t_L g265 ( .A(n_165), .Y(n_265) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_165), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_166), .A2(n_201), .B1(n_204), .B2(n_206), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_166), .A2(n_244), .B1(n_246), .B2(n_247), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_166), .A2(n_263), .B(n_264), .Y(n_262) );
OAI22x1_ASAP7_75t_L g553 ( .A1(n_166), .A2(n_554), .B1(n_555), .B2(n_556), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_166), .A2(n_556), .B1(n_577), .B2(n_579), .Y(n_576) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_166), .A2(n_247), .B1(n_649), .B2(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_168), .A2(n_180), .B1(n_224), .B2(n_225), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
INVx1_ASAP7_75t_L g285 ( .A(n_172), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_172), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g357 ( .A(n_172), .B(n_198), .Y(n_357) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_189), .Y(n_172) );
OA21x2_ASAP7_75t_L g195 ( .A1(n_173), .A2(n_174), .B(n_189), .Y(n_195) );
O2A1O1Ixp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B(n_179), .C(n_181), .Y(n_175) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_178), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g245 ( .A(n_180), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_180), .B(n_512), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_181), .A2(n_511), .B(n_513), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_185), .B1(n_187), .B2(n_188), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_184), .A2(n_543), .B(n_544), .C(n_545), .Y(n_542) );
INVx2_ASAP7_75t_SL g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx3_ASAP7_75t_L g231 ( .A(n_186), .Y(n_231) );
INVx2_ASAP7_75t_L g220 ( .A(n_190), .Y(n_220) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g322 ( .A(n_192), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_194), .B(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_194), .B(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_194), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_194), .B(n_392), .Y(n_399) );
INVx2_ASAP7_75t_SL g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g368 ( .A(n_195), .B(n_343), .Y(n_368) );
OR2x2_ASAP7_75t_L g370 ( .A(n_195), .B(n_296), .Y(n_370) );
INVx1_ASAP7_75t_L g429 ( .A(n_195), .Y(n_429) );
BUFx2_ASAP7_75t_L g443 ( .A(n_195), .Y(n_443) );
OR2x2_ASAP7_75t_L g471 ( .A(n_195), .B(n_198), .Y(n_471) );
INVx1_ASAP7_75t_L g490 ( .A(n_196), .Y(n_490) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g337 ( .A(n_197), .Y(n_337) );
OR2x2_ASAP7_75t_L g350 ( .A(n_197), .B(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g369 ( .A(n_197), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_212), .Y(n_197) );
INVx2_ASAP7_75t_L g289 ( .A(n_198), .Y(n_289) );
AND2x2_ASAP7_75t_L g305 ( .A(n_198), .B(n_212), .Y(n_305) );
INVx1_ASAP7_75t_L g343 ( .A(n_198), .Y(n_343) );
INVx1_ASAP7_75t_L g386 ( .A(n_198), .Y(n_386) );
AND2x2_ASAP7_75t_L g428 ( .A(n_198), .B(n_429), .Y(n_428) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .A3(n_207), .B(n_209), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_202), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g535 ( .A(n_202), .Y(n_535) );
INVx1_ASAP7_75t_SL g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g226 ( .A(n_205), .Y(n_226) );
INVx1_ASAP7_75t_L g556 ( .A(n_205), .Y(n_556) );
AO31x2_ASAP7_75t_L g575 ( .A1(n_207), .A2(n_508), .A3(n_576), .B(n_581), .Y(n_575) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_SL g240 ( .A(n_208), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g234 ( .A(n_211), .Y(n_234) );
BUFx2_ASAP7_75t_L g508 ( .A(n_211), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_211), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_211), .B(n_582), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_211), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g484 ( .A(n_214), .Y(n_484) );
AND2x4_ASAP7_75t_L g422 ( .A(n_215), .B(n_282), .Y(n_422) );
INVx2_ASAP7_75t_L g451 ( .A(n_215), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_215), .B(n_443), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_216), .B(n_441), .Y(n_440) );
AND2x4_ASAP7_75t_L g216 ( .A(n_217), .B(n_235), .Y(n_216) );
AND2x2_ASAP7_75t_L g362 ( .A(n_217), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g383 ( .A(n_217), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g254 ( .A(n_218), .B(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g278 ( .A(n_218), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g309 ( .A(n_218), .Y(n_309) );
AND2x2_ASAP7_75t_L g349 ( .A(n_218), .B(n_241), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_218), .B(n_333), .Y(n_390) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g302 ( .A(n_219), .Y(n_302) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_233), .Y(n_219) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_220), .A2(n_562), .B(n_571), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_227), .B(n_232), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_226), .Y(n_222) );
INVx2_ASAP7_75t_L g247 ( .A(n_231), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_232), .A2(n_510), .B(n_515), .Y(n_509) );
INVx3_ASAP7_75t_L g268 ( .A(n_235), .Y(n_268) );
AND2x2_ASAP7_75t_L g313 ( .A(n_235), .B(n_308), .Y(n_313) );
AND2x2_ASAP7_75t_L g468 ( .A(n_235), .B(n_272), .Y(n_468) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_241), .Y(n_235) );
INVx1_ASAP7_75t_L g319 ( .A(n_236), .Y(n_319) );
AND2x2_ASAP7_75t_L g347 ( .A(n_236), .B(n_255), .Y(n_347) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_240), .A2(n_259), .B(n_262), .Y(n_258) );
AND2x4_ASAP7_75t_L g300 ( .A(n_241), .B(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g273 ( .A(n_242), .B(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g310 ( .A(n_242), .B(n_274), .Y(n_310) );
AND2x2_ASAP7_75t_L g320 ( .A(n_242), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_242), .B(n_255), .Y(n_372) );
AND2x2_ASAP7_75t_L g378 ( .A(n_242), .B(n_302), .Y(n_378) );
AOI21x1_ASAP7_75t_L g259 ( .A1(n_247), .A2(n_260), .B(n_261), .Y(n_259) );
OAI21x1_ASAP7_75t_L g527 ( .A1(n_247), .A2(n_528), .B(n_531), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_247), .A2(n_606), .B(n_607), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_269), .Y(n_250) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_251), .A2(n_412), .B(n_416), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_251), .B(n_442), .Y(n_489) );
NAND2x1_ASAP7_75t_SL g252 ( .A(n_253), .B(n_267), .Y(n_252) );
INVx1_ASAP7_75t_L g495 ( .A(n_253), .Y(n_495) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g272 ( .A(n_255), .Y(n_272) );
INVx2_ASAP7_75t_L g277 ( .A(n_255), .Y(n_277) );
INVxp67_ASAP7_75t_L g298 ( .A(n_255), .Y(n_298) );
AND2x2_ASAP7_75t_L g318 ( .A(n_255), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g329 ( .A(n_255), .B(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g333 ( .A(n_255), .Y(n_333) );
INVx1_ASAP7_75t_L g351 ( .A(n_255), .Y(n_351) );
OR2x2_ASAP7_75t_L g384 ( .A(n_255), .B(n_319), .Y(n_384) );
INVx1_ASAP7_75t_L g455 ( .A(n_255), .Y(n_455) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_266), .Y(n_256) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI21xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_275), .B(n_280), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_271), .A2(n_394), .B1(n_396), .B2(n_399), .Y(n_393) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_272), .B(n_320), .Y(n_354) );
BUFx2_ASAP7_75t_L g413 ( .A(n_272), .Y(n_413) );
INVx2_ASAP7_75t_L g363 ( .A(n_273), .Y(n_363) );
OR2x2_ASAP7_75t_L g447 ( .A(n_273), .B(n_277), .Y(n_447) );
INVx1_ASAP7_75t_L g279 ( .A(n_274), .Y(n_279) );
INVx1_ASAP7_75t_L g328 ( .A(n_274), .Y(n_328) );
NOR2x1p5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVxp67_ASAP7_75t_SL g276 ( .A(n_277), .Y(n_276) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_277), .Y(n_398) );
OR2x2_ASAP7_75t_L g482 ( .A(n_277), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g485 ( .A(n_277), .B(n_320), .Y(n_485) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_278), .Y(n_448) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_282), .B(n_342), .Y(n_404) );
AND2x2_ASAP7_75t_L g494 ( .A(n_282), .B(n_292), .Y(n_494) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g403 ( .A(n_283), .B(n_292), .Y(n_403) );
NAND2x1p5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x2_ASAP7_75t_L g360 ( .A(n_284), .B(n_293), .Y(n_360) );
AND2x2_ASAP7_75t_L g395 ( .A(n_284), .B(n_289), .Y(n_395) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g314 ( .A(n_287), .B(n_295), .Y(n_314) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g454 ( .A(n_289), .B(n_455), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_303), .B2(n_306), .Y(n_290) );
O2A1O1Ixp33_ASAP7_75t_L g491 ( .A1(n_291), .A2(n_492), .B(n_493), .C(n_495), .Y(n_491) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g342 ( .A(n_293), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g410 ( .A(n_293), .Y(n_410) );
OR2x2_ASAP7_75t_L g457 ( .A(n_294), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_L g312 ( .A(n_298), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g415 ( .A(n_301), .Y(n_415) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g321 ( .A(n_302), .Y(n_321) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
INVx1_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g458 ( .A(n_305), .Y(n_458) );
AND2x2_ASAP7_75t_L g480 ( .A(n_305), .B(n_443), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_306), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g332 ( .A(n_310), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g388 ( .A(n_310), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_SL g483 ( .A(n_310), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_314), .B1(n_315), .B2(n_322), .C(n_323), .Y(n_311) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx2_ASAP7_75t_L g405 ( .A(n_318), .Y(n_405) );
BUFx2_ASAP7_75t_L g425 ( .A(n_320), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_331), .B(n_334), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
AND2x2_ASAP7_75t_L g467 ( .A(n_326), .B(n_389), .Y(n_467) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
AND2x2_ASAP7_75t_L g463 ( .A(n_328), .B(n_333), .Y(n_463) );
INVx1_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI211xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B(n_352), .C(n_364), .Y(n_338) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B1(n_348), .B2(n_350), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
BUFx2_ASAP7_75t_L g380 ( .A(n_347), .Y(n_380) );
AND2x2_ASAP7_75t_L g473 ( .A(n_347), .B(n_415), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g476 ( .A1(n_348), .A2(n_477), .B(n_479), .Y(n_476) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_355), .B1(n_359), .B2(n_361), .Y(n_352) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_355), .B(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g427 ( .A(n_360), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x4_ASAP7_75t_L g414 ( .A(n_363), .B(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_363), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B(n_371), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
AND2x2_ASAP7_75t_L g441 ( .A(n_366), .B(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g478 ( .A(n_366), .B(n_443), .Y(n_478) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g392 ( .A(n_367), .Y(n_392) );
OR2x2_ASAP7_75t_L g470 ( .A(n_367), .B(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g385 ( .A(n_370), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g417 ( .A(n_370), .Y(n_417) );
OR2x2_ASAP7_75t_L g450 ( .A(n_370), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g421 ( .A(n_371), .Y(n_421) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NOR3xp33_ASAP7_75t_L g374 ( .A(n_375), .B(n_393), .C(n_400), .Y(n_374) );
OAI322xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .A3(n_381), .B1(n_383), .B2(n_385), .C1(n_387), .C2(n_391), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
A2O1A1Ixp33_ASAP7_75t_L g452 ( .A1(n_377), .A2(n_417), .B(n_453), .C(n_456), .Y(n_452) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g397 ( .A(n_378), .B(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g434 ( .A(n_378), .Y(n_434) );
AND2x4_ASAP7_75t_L g462 ( .A(n_378), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g431 ( .A1(n_380), .A2(n_418), .A3(n_432), .B1(n_434), .B2(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g418 ( .A(n_384), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_386), .B(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_404), .C(n_405), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_464), .Y(n_406) );
AOI211xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_411), .B(n_419), .C(n_444), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_412), .A2(n_487), .B(n_488), .C(n_490), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_414), .A2(n_467), .A3(n_468), .B(n_469), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx2_ASAP7_75t_L g426 ( .A(n_418), .Y(n_426) );
NAND4xp25_ASAP7_75t_SL g419 ( .A(n_420), .B(n_423), .C(n_431), .D(n_440), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI32xp33_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .A3(n_426), .B1(n_427), .B2(n_430), .Y(n_423) );
INVx1_ASAP7_75t_L g475 ( .A(n_427), .Y(n_475) );
INVx1_ASAP7_75t_L g487 ( .A(n_430), .Y(n_487) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_445), .B(n_452), .C(n_459), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_448), .B(n_449), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_453), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_476), .C(n_486), .D(n_491), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_472), .Y(n_465) );
OAI21xp33_ASAP7_75t_L g472 ( .A1(n_467), .A2(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B1(n_484), .B2(n_485), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_483), .Y(n_492) );
INVxp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx8_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_497), .Y(n_501) );
AND2x2_ASAP7_75t_L g855 ( .A(n_497), .B(n_856), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx12f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
XNOR2x1_ASAP7_75t_L g842 ( .A(n_502), .B(n_843), .Y(n_842) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_720), .Y(n_502) );
NAND3xp33_ASAP7_75t_SL g503 ( .A(n_504), .B(n_623), .C(n_682), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_520), .B1(n_610), .B2(n_616), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OR2x2_ASAP7_75t_L g679 ( .A(n_506), .B(n_680), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_506), .B(n_597), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_506), .B(n_643), .Y(n_790) );
AND2x2_ASAP7_75t_L g796 ( .A(n_506), .B(n_622), .Y(n_796) );
INVxp67_ASAP7_75t_L g801 ( .A(n_506), .Y(n_801) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g614 ( .A(n_507), .Y(n_614) );
AOI21x1_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B(n_519), .Y(n_507) );
INVx4_ASAP7_75t_L g543 ( .A(n_516), .Y(n_543) );
OAI21xp5_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_572), .B(n_583), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_551), .Y(n_522) );
INVx1_ASAP7_75t_L g717 ( .A(n_523), .Y(n_717) );
AND2x2_ASAP7_75t_L g746 ( .A(n_523), .B(n_708), .Y(n_746) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_538), .Y(n_523) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_561), .Y(n_640) );
INVx1_ASAP7_75t_L g695 ( .A(n_524), .Y(n_695) );
AND2x2_ASAP7_75t_L g745 ( .A(n_524), .B(n_560), .Y(n_745) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g620 ( .A(n_525), .B(n_560), .Y(n_620) );
AND2x4_ASAP7_75t_L g764 ( .A(n_525), .B(n_561), .Y(n_764) );
AOI21x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_532), .B(n_536), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_530), .B(n_565), .Y(n_564) );
OAI21xp33_ASAP7_75t_SL g600 ( .A1(n_535), .A2(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g689 ( .A(n_538), .Y(n_689) );
AND2x2_ASAP7_75t_L g758 ( .A(n_538), .B(n_561), .Y(n_758) );
AND2x2_ASAP7_75t_L g765 ( .A(n_538), .B(n_591), .Y(n_765) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g587 ( .A(n_539), .Y(n_587) );
BUFx3_ASAP7_75t_L g622 ( .A(n_539), .Y(n_622) );
AND2x2_ASAP7_75t_L g633 ( .A(n_539), .B(n_619), .Y(n_633) );
AND2x2_ASAP7_75t_L g696 ( .A(n_539), .B(n_552), .Y(n_696) );
AND2x2_ASAP7_75t_L g701 ( .A(n_539), .B(n_561), .Y(n_701) );
NAND2x1p5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
OAI21x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_546), .B(n_549), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_551), .B(n_707), .Y(n_809) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_560), .Y(n_551) );
INVx2_ASAP7_75t_L g591 ( .A(n_552), .Y(n_591) );
OR2x2_ASAP7_75t_L g594 ( .A(n_552), .B(n_561), .Y(n_594) );
INVx2_ASAP7_75t_L g619 ( .A(n_552), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_552), .B(n_589), .Y(n_635) );
AND2x2_ASAP7_75t_L g708 ( .A(n_552), .B(n_561), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_556), .B(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g570 ( .A(n_557), .Y(n_570) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g636 ( .A(n_561), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B(n_570), .Y(n_562) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_573), .B(n_671), .Y(n_817) );
BUFx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g629 ( .A(n_574), .Y(n_629) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g609 ( .A(n_575), .Y(n_609) );
AND2x2_ASAP7_75t_L g615 ( .A(n_575), .B(n_597), .Y(n_615) );
INVx1_ASAP7_75t_L g663 ( .A(n_575), .Y(n_663) );
OR2x2_ASAP7_75t_L g668 ( .A(n_575), .B(n_647), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_575), .B(n_647), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_575), .B(n_646), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_575), .B(n_614), .Y(n_753) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_592), .B(n_595), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
OR2x2_ASAP7_75t_L g593 ( .A(n_586), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g744 ( .A(n_586), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g774 ( .A(n_586), .B(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_587), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g742 ( .A(n_587), .Y(n_742) );
OR2x2_ASAP7_75t_L g655 ( .A(n_588), .B(n_656), .Y(n_655) );
INVxp33_ASAP7_75t_L g773 ( .A(n_588), .Y(n_773) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVx2_ASAP7_75t_L g677 ( .A(n_589), .Y(n_677) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g631 ( .A(n_591), .Y(n_631) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_SL g739 ( .A1(n_593), .A2(n_664), .B1(n_669), .B2(n_740), .C(n_743), .Y(n_739) );
OR2x2_ASAP7_75t_L g726 ( .A(n_594), .B(n_677), .Y(n_726) );
INVx2_ASAP7_75t_L g775 ( .A(n_594), .Y(n_775) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g675 ( .A(n_596), .Y(n_675) );
OR2x2_ASAP7_75t_L g678 ( .A(n_596), .B(n_679), .Y(n_678) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_596), .Y(n_719) );
OR2x2_ASAP7_75t_L g732 ( .A(n_596), .B(n_733), .Y(n_732) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_609), .Y(n_596) );
NAND2x1p5_ASAP7_75t_SL g628 ( .A(n_597), .B(n_613), .Y(n_628) );
INVx3_ASAP7_75t_L g643 ( .A(n_597), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_597), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g666 ( .A(n_597), .Y(n_666) );
AND2x2_ASAP7_75t_L g747 ( .A(n_597), .B(n_748), .Y(n_747) );
AND2x2_ASAP7_75t_L g754 ( .A(n_597), .B(n_661), .Y(n_754) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_605), .B(n_608), .Y(n_599) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_615), .Y(n_610) );
AND2x2_ASAP7_75t_L g806 ( .A(n_611), .B(n_665), .Y(n_806) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g710 ( .A(n_613), .B(n_680), .Y(n_710) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g645 ( .A(n_614), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g671 ( .A(n_614), .B(n_647), .Y(n_671) );
AND2x4_ASAP7_75t_L g768 ( .A(n_615), .B(n_738), .Y(n_768) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g687 ( .A(n_620), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_621), .B(n_708), .Y(n_792) );
AND2x2_ASAP7_75t_L g799 ( .A(n_621), .B(n_759), .Y(n_799) );
INVx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx2_ASAP7_75t_L g724 ( .A(n_622), .Y(n_724) );
AOI321xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_637), .A3(n_653), .B1(n_654), .B2(n_657), .C(n_672), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_625), .B(n_634), .Y(n_624) );
AOI21xp33_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_630), .B(n_632), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g637 ( .A1(n_627), .A2(n_638), .B(n_641), .Y(n_637) );
OR2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OR2x2_ASAP7_75t_L g736 ( .A(n_628), .B(n_668), .Y(n_736) );
INVx1_ASAP7_75t_L g728 ( .A(n_629), .Y(n_728) );
INVx2_ASAP7_75t_L g713 ( .A(n_630), .Y(n_713) );
OAI32xp33_ASAP7_75t_L g816 ( .A1(n_630), .A2(n_778), .A3(n_789), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g731 ( .A(n_631), .Y(n_731) );
INVx1_ASAP7_75t_L g681 ( .A(n_632), .Y(n_681) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x4_ASAP7_75t_SL g769 ( .A(n_633), .B(n_676), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_634), .B(n_638), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_634), .A2(n_710), .B1(n_771), .B2(n_792), .Y(n_791) );
OR2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g759 ( .A(n_635), .Y(n_759) );
INVx1_ASAP7_75t_L g656 ( .A(n_636), .Y(n_656) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g741 ( .A(n_640), .Y(n_741) );
NAND4xp25_ASAP7_75t_L g657 ( .A(n_641), .B(n_658), .C(n_664), .D(n_669), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVxp67_ASAP7_75t_L g683 ( .A(n_642), .Y(n_683) );
AND2x2_ASAP7_75t_L g762 ( .A(n_642), .B(n_671), .Y(n_762) );
OR2x2_ASAP7_75t_L g771 ( .A(n_642), .B(n_645), .Y(n_771) );
AND2x2_ASAP7_75t_L g795 ( .A(n_642), .B(n_667), .Y(n_795) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g709 ( .A(n_643), .B(n_710), .Y(n_709) );
AND2x4_ASAP7_75t_L g716 ( .A(n_643), .B(n_663), .Y(n_716) );
INVx1_ASAP7_75t_L g780 ( .A(n_644), .Y(n_780) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g688 ( .A(n_645), .B(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g738 ( .A(n_645), .Y(n_738) );
INVx1_ASAP7_75t_L g680 ( .A(n_646), .Y(n_680) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g661 ( .A(n_647), .Y(n_661) );
INVx3_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .Y(n_659) );
AND2x4_ASAP7_75t_L g674 ( .A(n_660), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g715 ( .A(n_660), .Y(n_715) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_662), .Y(n_779) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
AND2x2_ASAP7_75t_L g670 ( .A(n_666), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g756 ( .A(n_668), .Y(n_756) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g733 ( .A(n_671), .Y(n_733) );
AND2x2_ASAP7_75t_L g776 ( .A(n_671), .B(n_716), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_676), .B(n_678), .C(n_681), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g787 ( .A(n_676), .B(n_765), .Y(n_787) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g691 ( .A(n_679), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B(n_697), .C(n_711), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_688), .B(n_690), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g793 ( .A1(n_686), .A2(n_794), .B(n_797), .Y(n_793) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g707 ( .A(n_689), .Y(n_707) );
AND2x2_ASAP7_75t_L g767 ( .A(n_689), .B(n_764), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g786 ( .A(n_694), .Y(n_786) );
AND2x2_ASAP7_75t_L g812 ( .A(n_694), .B(n_775), .Y(n_812) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_695), .Y(n_700) );
INVx2_ASAP7_75t_L g751 ( .A(n_696), .Y(n_751) );
NAND2x1_ASAP7_75t_L g785 ( .A(n_696), .B(n_786), .Y(n_785) );
AOI33xp33_ASAP7_75t_L g803 ( .A1(n_696), .A2(n_716), .A3(n_754), .B1(n_764), .B2(n_796), .B3(n_867), .Y(n_803) );
OAI22xp33_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_702), .B1(n_705), .B2(n_709), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
AND2x2_ASAP7_75t_L g730 ( .A(n_701), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_702), .B(n_789), .Y(n_788) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
OR2x2_ASAP7_75t_L g815 ( .A(n_704), .B(n_749), .Y(n_815) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
OAI22xp33_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_714), .B1(n_717), .B2(n_718), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_715), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_715), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g737 ( .A(n_716), .B(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g802 ( .A(n_716), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_781), .Y(n_720) );
NOR4xp25_ASAP7_75t_L g721 ( .A(n_722), .B(n_739), .C(n_760), .D(n_777), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_727), .B1(n_729), .B2(n_732), .C(n_734), .Y(n_722) );
O2A1O1Ixp33_ASAP7_75t_SL g777 ( .A1(n_723), .A2(n_778), .B(n_779), .C(n_780), .Y(n_777) );
NAND2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g810 ( .A(n_726), .Y(n_810) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g734 ( .A1(n_730), .A2(n_735), .B(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OR2x6_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_746), .B(n_747), .C(n_750), .Y(n_743) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OR2x2_ASAP7_75t_L g789 ( .A(n_749), .B(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_SL g813 ( .A(n_749), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_752), .B1(n_755), .B2(n_757), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_763), .B(n_766), .C(n_772), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_764), .A2(n_812), .B1(n_813), .B2(n_814), .C(n_816), .Y(n_811) );
INVx3_ASAP7_75t_L g819 ( .A(n_764), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_766) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI21xp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B(n_776), .Y(n_772) );
INVx1_ASAP7_75t_L g778 ( .A(n_775), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_804), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_793), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B(n_788), .C(n_791), .Y(n_783) );
INVx2_ASAP7_75t_SL g784 ( .A(n_785), .Y(n_784) );
NOR3xp33_ASAP7_75t_L g807 ( .A(n_787), .B(n_808), .C(n_810), .Y(n_807) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
OAI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_800), .B(n_803), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
OR2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B(n_811), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx3_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx6_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x6_ASAP7_75t_SL g827 ( .A(n_828), .B(n_830), .Y(n_827) );
BUFx3_ASAP7_75t_L g836 ( .A(n_828), .Y(n_836) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_829), .B(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2x1_ASAP7_75t_L g856 ( .A(n_832), .B(n_834), .Y(n_856) );
AND2x6_ASAP7_75t_SL g859 ( .A(n_833), .B(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
OAI21xp33_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_837), .B(n_849), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_842), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx4_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AOI22x1_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_848), .Y(n_847) );
INVx3_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx6_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx10_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_862), .Y(n_857) );
INVx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_R g863 ( .A(n_864), .B(n_865), .Y(n_863) );
endmodule