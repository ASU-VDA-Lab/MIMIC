module real_aes_16944_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_93;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OAI22xp33_ASAP7_75t_SL g571 ( .A1(n_0), .A2(n_37), .B1(n_572), .B2(n_575), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_0), .A2(n_7), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_1), .A2(n_32), .B1(n_115), .B2(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_2), .B(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g542 ( .A(n_2), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_3), .A2(n_13), .B1(n_108), .B2(n_222), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_4), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_5), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_6), .Y(n_489) );
OAI22xp33_ASAP7_75t_SL g564 ( .A1(n_7), .A2(n_67), .B1(n_565), .B2(n_568), .Y(n_564) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_8), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_9), .A2(n_14), .B1(n_89), .B2(n_148), .Y(n_147) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_10), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_11), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g497 ( .A(n_12), .Y(n_497) );
INVx1_ASAP7_75t_L g470 ( .A(n_15), .Y(n_470) );
INVx1_ASAP7_75t_L g476 ( .A(n_15), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_16), .A2(n_76), .B1(n_108), .B2(n_110), .Y(n_107) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_17), .A2(n_29), .B1(n_191), .B2(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g463 ( .A(n_18), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_19), .B(n_109), .Y(n_188) );
OAI21x1_ASAP7_75t_L g123 ( .A1(n_20), .A2(n_40), .B(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_21), .Y(n_126) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_22), .A2(n_35), .B1(n_132), .B2(n_135), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_23), .A2(n_39), .B1(n_108), .B2(n_135), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_24), .Y(n_206) );
INVx1_ASAP7_75t_L g554 ( .A(n_25), .Y(n_554) );
OAI211xp5_ASAP7_75t_SL g589 ( .A1(n_25), .A2(n_590), .B(n_595), .C(n_605), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_26), .B(n_191), .Y(n_190) );
BUFx2_ASAP7_75t_L g635 ( .A(n_26), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_27), .Y(n_180) );
INVx1_ASAP7_75t_L g638 ( .A(n_28), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_30), .A2(n_63), .B1(n_115), .B2(n_200), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_31), .A2(n_34), .B1(n_115), .B2(n_150), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_33), .A2(n_41), .B1(n_108), .B2(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g462 ( .A(n_36), .Y(n_462) );
INVx1_ASAP7_75t_L g506 ( .A(n_36), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_37), .A2(n_67), .B1(n_586), .B2(n_588), .Y(n_585) );
INVx2_ASAP7_75t_L g648 ( .A(n_38), .Y(n_648) );
BUFx3_ASAP7_75t_L g468 ( .A(n_42), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_43), .A2(n_55), .B1(n_114), .B2(n_132), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_44), .A2(n_57), .B1(n_115), .B2(n_150), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_45), .A2(n_74), .B1(n_108), .B2(n_148), .Y(n_177) );
AND2x4_ASAP7_75t_L g82 ( .A(n_46), .B(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_46), .Y(n_622) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_48), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g630 ( .A(n_49), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_50), .Y(n_479) );
INVx1_ASAP7_75t_L g83 ( .A(n_51), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_52), .Y(n_501) );
OAI211xp5_ASAP7_75t_L g544 ( .A1(n_53), .A2(n_545), .B(n_546), .C(n_553), .Y(n_544) );
INVx1_ASAP7_75t_L g604 ( .A(n_53), .Y(n_604) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_54), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_56), .Y(n_471) );
INVx2_ASAP7_75t_L g87 ( .A(n_58), .Y(n_87) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_59), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_59), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_60), .A2(n_75), .B1(n_135), .B2(n_203), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_61), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_62), .Y(n_172) );
BUFx3_ASAP7_75t_L g512 ( .A(n_64), .Y(n_512) );
INVx1_ASAP7_75t_L g574 ( .A(n_64), .Y(n_574) );
XNOR2xp5_ASAP7_75t_L g450 ( .A(n_65), .B(n_451), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_66), .Y(n_558) );
INVx1_ASAP7_75t_L g460 ( .A(n_68), .Y(n_460) );
INVx2_ASAP7_75t_L g504 ( .A(n_68), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_69), .B(n_169), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_70), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_71), .Y(n_493) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_72), .B(n_109), .Y(n_192) );
INVx1_ASAP7_75t_L g636 ( .A(n_73), .Y(n_636) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_74), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_93), .B(n_449), .Y(n_77) );
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_84), .Y(n_80) );
INVx2_ASAP7_75t_L g105 ( .A(n_81), .Y(n_105) );
AO31x2_ASAP7_75t_L g145 ( .A1(n_81), .A2(n_146), .A3(n_153), .B(n_155), .Y(n_145) );
AO31x2_ASAP7_75t_L g163 ( .A1(n_81), .A2(n_164), .A3(n_168), .B(n_171), .Y(n_163) );
AO31x2_ASAP7_75t_L g216 ( .A1(n_81), .A2(n_197), .A3(n_217), .B(n_224), .Y(n_216) );
BUFx10_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_L g137 ( .A(n_82), .Y(n_137) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_83), .Y(n_624) );
INVxp67_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AO21x1_ASAP7_75t_L g668 ( .A1(n_85), .A2(n_623), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_86), .B(n_88), .Y(n_85) );
INVx6_ASAP7_75t_L g112 ( .A(n_86), .Y(n_112) );
O2A1O1Ixp5_ASAP7_75t_L g186 ( .A1(n_86), .A2(n_150), .B(n_187), .C(n_188), .Y(n_186) );
BUFx8_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g118 ( .A(n_87), .Y(n_118) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_92), .Y(n_109) );
INVx1_ASAP7_75t_L g111 ( .A(n_92), .Y(n_111) );
INVx3_ASAP7_75t_L g115 ( .A(n_92), .Y(n_115) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_92), .Y(n_133) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_92), .Y(n_166) );
INVx2_ASAP7_75t_L g201 ( .A(n_92), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_92), .Y(n_203) );
INVx1_ASAP7_75t_L g220 ( .A(n_92), .Y(n_220) );
INVx1_ASAP7_75t_L g223 ( .A(n_92), .Y(n_223) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND3x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_311), .C(n_365), .Y(n_95) );
NOR2x1_ASAP7_75t_L g96 ( .A(n_97), .B(n_271), .Y(n_96) );
NAND3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_207), .C(n_253), .Y(n_97) );
OAI21xp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_140), .B(n_158), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OR2x2_ASAP7_75t_L g303 ( .A(n_101), .B(n_211), .Y(n_303) );
INVx2_ASAP7_75t_L g329 ( .A(n_101), .Y(n_329) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_128), .Y(n_101) );
INVx1_ASAP7_75t_L g228 ( .A(n_102), .Y(n_228) );
INVx2_ASAP7_75t_L g343 ( .A(n_102), .Y(n_343) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
AND2x4_ASAP7_75t_L g286 ( .A(n_103), .B(n_248), .Y(n_286) );
AO31x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_106), .A3(n_119), .B(n_125), .Y(n_103) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_104), .A2(n_153), .A3(n_176), .B(n_179), .Y(n_175) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_112), .B1(n_113), .B2(n_116), .Y(n_106) );
INVx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_112), .A2(n_116), .B1(n_131), .B2(n_134), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_112), .A2(n_147), .B1(n_149), .B2(n_151), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_112), .A2(n_116), .B1(n_165), .B2(n_167), .Y(n_164) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_112), .A2(n_151), .B1(n_177), .B2(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_112), .A2(n_190), .B(n_192), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_112), .A2(n_199), .B1(n_202), .B2(n_204), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_112), .A2(n_116), .B1(n_218), .B2(n_221), .Y(n_217) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g148 ( .A(n_115), .Y(n_148) );
INVx4_ASAP7_75t_L g150 ( .A(n_115), .Y(n_150) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AO31x2_ASAP7_75t_L g129 ( .A1(n_119), .A2(n_130), .A3(n_136), .B(n_138), .Y(n_129) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp33_ASAP7_75t_SL g155 ( .A(n_121), .B(n_156), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_121), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g127 ( .A(n_122), .Y(n_127) );
INVx2_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_123), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_127), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g339 ( .A(n_128), .Y(n_339) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
AND2x4_ASAP7_75t_L g214 ( .A(n_129), .B(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_129), .Y(n_245) );
INVx2_ASAP7_75t_L g248 ( .A(n_129), .Y(n_248) );
OR2x2_ASAP7_75t_L g262 ( .A(n_129), .B(n_216), .Y(n_262) );
AND2x2_ASAP7_75t_L g364 ( .A(n_129), .B(n_145), .Y(n_364) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
AO31x2_ASAP7_75t_L g196 ( .A1(n_136), .A2(n_197), .A3(n_198), .B(n_205), .Y(n_196) );
INVx2_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_SL g193 ( .A(n_137), .Y(n_193) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_141), .B(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
OR2x2_ASAP7_75t_L g246 ( .A(n_142), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_142), .B(n_265), .Y(n_310) );
AND2x2_ASAP7_75t_L g375 ( .A(n_142), .B(n_351), .Y(n_375) );
INVx4_ASAP7_75t_L g409 ( .A(n_142), .Y(n_409) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g244 ( .A(n_143), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g282 ( .A(n_143), .B(n_213), .Y(n_282) );
AND2x2_ASAP7_75t_L g392 ( .A(n_143), .B(n_216), .Y(n_392) );
AND2x2_ASAP7_75t_L g426 ( .A(n_143), .B(n_248), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_145), .B(n_157), .Y(n_144) );
INVx4_ASAP7_75t_SL g213 ( .A(n_145), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_145), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g327 ( .A(n_145), .B(n_216), .Y(n_327) );
BUFx2_ASAP7_75t_L g345 ( .A(n_145), .Y(n_345) );
INVx1_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g204 ( .A(n_152), .Y(n_204) );
BUFx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI222xp33_ASAP7_75t_L g253 ( .A1(n_157), .A2(n_254), .B1(n_259), .B2(n_260), .C1(n_263), .C2(n_267), .Y(n_253) );
INVx1_ASAP7_75t_L g384 ( .A(n_157), .Y(n_384) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_173), .Y(n_158) );
AND2x2_ASAP7_75t_L g421 ( .A(n_159), .B(n_233), .Y(n_421) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g442 ( .A(n_160), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g251 ( .A(n_161), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_161), .B(n_234), .Y(n_390) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_162), .B(n_238), .Y(n_280) );
AND2x2_ASAP7_75t_L g308 ( .A(n_162), .B(n_182), .Y(n_308) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g237 ( .A(n_163), .B(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g270 ( .A(n_163), .B(n_196), .Y(n_270) );
INVx1_ASAP7_75t_L g298 ( .A(n_163), .Y(n_298) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_163), .Y(n_404) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_170), .B(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_170), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_SL g184 ( .A(n_170), .Y(n_184) );
BUFx3_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_170), .B(n_225), .Y(n_224) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_173), .A2(n_296), .B1(n_354), .B2(n_355), .C1(n_357), .C2(n_359), .Y(n_353) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_181), .Y(n_173) );
INVx1_ASAP7_75t_L g288 ( .A(n_174), .Y(n_288) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx3_ASAP7_75t_L g234 ( .A(n_175), .Y(n_234) );
AND2x2_ASAP7_75t_L g239 ( .A(n_175), .B(n_196), .Y(n_239) );
AND2x2_ASAP7_75t_L g299 ( .A(n_175), .B(n_195), .Y(n_299) );
AND2x2_ASAP7_75t_L g287 ( .A(n_181), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g382 ( .A(n_181), .B(n_298), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_181), .B(n_389), .Y(n_388) );
AND3x1_ASAP7_75t_L g447 ( .A(n_181), .B(n_214), .C(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_195), .Y(n_181) );
AND2x2_ASAP7_75t_L g268 ( .A(n_182), .B(n_234), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_182), .B(n_370), .Y(n_417) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g231 ( .A(n_183), .Y(n_231) );
OAI21x1_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_194), .Y(n_183) );
OAI21x1_ASAP7_75t_L g238 ( .A1(n_184), .A2(n_185), .B(n_194), .Y(n_238) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_189), .B(n_193), .Y(n_185) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x4_ASAP7_75t_L g233 ( .A(n_196), .B(n_234), .Y(n_233) );
OR2x2_ASAP7_75t_L g266 ( .A(n_196), .B(n_252), .Y(n_266) );
INVx1_ASAP7_75t_L g276 ( .A(n_196), .Y(n_276) );
BUFx2_ASAP7_75t_L g370 ( .A(n_196), .Y(n_370) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_229), .B(n_235), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2x1_ASAP7_75t_L g209 ( .A(n_210), .B(n_226), .Y(n_209) );
AOI221xp5_ASAP7_75t_SL g293 ( .A1(n_210), .A2(n_294), .B1(n_300), .B2(n_304), .C(n_309), .Y(n_293) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_212), .B(n_228), .Y(n_414) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_213), .B(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g256 ( .A(n_213), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g292 ( .A(n_213), .Y(n_292) );
INVx1_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
AND2x2_ASAP7_75t_L g321 ( .A(n_213), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g333 ( .A(n_213), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_213), .B(n_339), .Y(n_446) );
INVx2_ASAP7_75t_L g281 ( .A(n_214), .Y(n_281) );
AND2x2_ASAP7_75t_L g291 ( .A(n_214), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_214), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_214), .B(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_216), .Y(n_285) );
INVx1_ASAP7_75t_L g322 ( .A(n_216), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_216), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g261 ( .A(n_227), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_227), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_228), .Y(n_320) );
NOR2xp33_ASAP7_75t_R g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR3xp33_ASAP7_75t_L g309 ( .A(n_231), .B(n_301), .C(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g332 ( .A(n_231), .B(n_239), .Y(n_332) );
AND2x2_ASAP7_75t_L g361 ( .A(n_231), .B(n_331), .Y(n_361) );
OR2x2_ASAP7_75t_L g428 ( .A(n_231), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x4_ASAP7_75t_L g354 ( .A(n_233), .B(n_237), .Y(n_354) );
INVx2_ASAP7_75t_SL g438 ( .A(n_233), .Y(n_438) );
INVx2_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_234), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g307 ( .A(n_234), .Y(n_307) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_234), .Y(n_380) );
OAI32xp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_240), .A3(n_243), .B1(n_246), .B2(n_249), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
AND2x2_ASAP7_75t_L g259 ( .A(n_237), .B(n_239), .Y(n_259) );
AND2x2_ASAP7_75t_L g317 ( .A(n_237), .B(n_299), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_237), .B(n_299), .Y(n_325) );
INVx1_ASAP7_75t_L g252 ( .A(n_238), .Y(n_252) );
AND2x4_ASAP7_75t_SL g250 ( .A(n_239), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g394 ( .A(n_239), .Y(n_394) );
INVx2_ASAP7_75t_L g429 ( .A(n_239), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_239), .B(n_308), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g371 ( .A(n_240), .B(n_362), .C(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g257 ( .A(n_242), .Y(n_257) );
AOI321xp33_ASAP7_75t_L g440 ( .A1(n_243), .A2(n_302), .A3(n_441), .B1(n_442), .B2(n_444), .C(n_447), .Y(n_440) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g258 ( .A(n_245), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_247), .A2(n_266), .B1(n_445), .B2(n_446), .Y(n_444) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g347 ( .A(n_251), .B(n_306), .Y(n_347) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_256), .B(n_258), .Y(n_255) );
INVx1_ASAP7_75t_L g381 ( .A(n_256), .Y(n_381) );
NAND2x1_ASAP7_75t_L g408 ( .A(n_256), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_256), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g406 ( .A(n_258), .B(n_392), .Y(n_406) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g346 ( .A(n_262), .Y(n_346) );
OR2x2_ASAP7_75t_L g413 ( .A(n_262), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_265), .B(n_266), .Y(n_290) );
NOR2x1p5_ASAP7_75t_L g331 ( .A(n_265), .B(n_270), .Y(n_331) );
INVx1_ASAP7_75t_L g401 ( .A(n_265), .Y(n_401) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_266), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_268), .Y(n_445) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_283), .C(n_293), .Y(n_271) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_281), .C(n_282), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g423 ( .A(n_277), .Y(n_423) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g315 ( .A(n_280), .Y(n_315) );
INVx1_ASAP7_75t_L g351 ( .A(n_280), .Y(n_351) );
NAND2xp33_ASAP7_75t_L g355 ( .A(n_281), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_281), .Y(n_359) );
INVx1_ASAP7_75t_L g385 ( .A(n_282), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_287), .B(n_289), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx3_ASAP7_75t_L g334 ( .A(n_286), .Y(n_334) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g411 ( .A(n_298), .B(n_401), .Y(n_411) );
AND2x2_ASAP7_75t_L g314 ( .A(n_299), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g379 ( .A(n_299), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
OR2x2_ASAP7_75t_L g337 ( .A(n_302), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g316 ( .A(n_303), .Y(n_316) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g350 ( .A(n_307), .B(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g439 ( .A(n_308), .Y(n_439) );
NOR2xp67_ASAP7_75t_L g311 ( .A(n_312), .B(n_348), .Y(n_311) );
NAND3xp33_ASAP7_75t_SL g312 ( .A(n_313), .B(n_323), .C(n_335), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_317), .B2(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g356 ( .A(n_321), .Y(n_356) );
AND2x2_ASAP7_75t_L g431 ( .A(n_321), .B(n_342), .Y(n_431) );
INVx1_ASAP7_75t_L g378 ( .A(n_322), .Y(n_378) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .A3(n_328), .B1(n_330), .B2(n_333), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
NAND2x1_ASAP7_75t_L g396 ( .A(n_327), .B(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g357 ( .A(n_329), .B(n_358), .Y(n_357) );
NOR2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_334), .A2(n_377), .B(n_384), .C(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g397 ( .A(n_334), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B(n_347), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_341), .Y(n_352) );
NAND2x1_ASAP7_75t_L g341 ( .A(n_342), .B(n_344), .Y(n_341) );
INVx2_ASAP7_75t_L g435 ( .A(n_342), .Y(n_435) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g443 ( .A(n_343), .B(n_378), .Y(n_443) );
AND2x2_ASAP7_75t_L g448 ( .A(n_343), .B(n_404), .Y(n_448) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
OAI211xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B(n_353), .C(n_360), .Y(n_348) );
INVxp67_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g367 ( .A(n_350), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_398), .C(n_427), .Y(n_365) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B(n_374), .C(n_386), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_372), .A2(n_411), .B1(n_412), .B2(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_376), .B1(n_382), .B2(n_383), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B1(n_380), .B2(n_381), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_377), .B(n_409), .Y(n_420) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g391 ( .A(n_384), .B(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_391), .B1(n_393), .B2(n_395), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g416 ( .A(n_390), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_405), .B(n_410), .C(n_418), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B1(n_422), .B2(n_424), .Y(n_418) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI211xp5_ASAP7_75t_SL g427 ( .A1(n_428), .A2(n_430), .B(n_432), .C(n_440), .Y(n_427) );
INVxp67_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_618), .B2(n_625), .C(n_662), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_451), .A2(n_656), .B1(n_663), .B2(n_666), .Y(n_662) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_543), .C(n_584), .Y(n_453) );
NOR2xp33_ASAP7_75t_SL g454 ( .A(n_455), .B(n_508), .Y(n_454) );
OAI33xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_464), .A3(n_478), .B1(n_490), .B2(n_498), .B3(n_502), .Y(n_455) );
BUFx4f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .Y(n_457) );
AND2x2_ASAP7_75t_SL g540 ( .A(n_458), .B(n_541), .Y(n_540) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_458), .Y(n_617) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g583 ( .A(n_459), .Y(n_583) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx2_ASAP7_75t_L g653 ( .A(n_461), .Y(n_653) );
NAND2xp33_ASAP7_75t_SL g461 ( .A(n_462), .B(n_463), .Y(n_461) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_462), .Y(n_615) );
INVx1_ASAP7_75t_L g647 ( .A(n_462), .Y(n_647) );
INVx3_ASAP7_75t_L g507 ( .A(n_463), .Y(n_507) );
BUFx3_ASAP7_75t_L g593 ( .A(n_463), .Y(n_593) );
OAI22xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B1(n_471), .B2(n_472), .Y(n_464) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_465), .A2(n_499), .B1(n_514), .B2(n_520), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_466), .A2(n_499), .B1(n_500), .B2(n_501), .Y(n_498) );
BUFx4f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x4_ASAP7_75t_L g586 ( .A(n_467), .B(n_587), .Y(n_586) );
OR2x4_ASAP7_75t_L g609 ( .A(n_467), .B(n_507), .Y(n_609) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_468), .Y(n_477) );
INVx2_ASAP7_75t_L g484 ( .A(n_468), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_468), .B(n_476), .Y(n_488) );
AND2x4_ASAP7_75t_L g607 ( .A(n_468), .B(n_599), .Y(n_607) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_L g483 ( .A(n_470), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_471), .A2(n_501), .B1(n_526), .B2(n_530), .Y(n_534) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx3_ASAP7_75t_L g500 ( .A(n_474), .Y(n_500) );
NAND2x1p5_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
BUFx2_ASAP7_75t_L g603 ( .A(n_475), .Y(n_603) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g599 ( .A(n_476), .Y(n_599) );
BUFx2_ASAP7_75t_L g594 ( .A(n_477), .Y(n_594) );
INVx2_ASAP7_75t_L g601 ( .A(n_477), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_485), .B2(n_489), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_479), .A2(n_493), .B1(n_526), .B2(n_530), .Y(n_525) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
BUFx8_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_482), .Y(n_492) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_482), .Y(n_612) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x6_ASAP7_75t_L g588 ( .A(n_487), .B(n_507), .Y(n_588) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_488), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g535 ( .A1(n_489), .A2(n_497), .B1(n_520), .B2(n_536), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_493), .B1(n_494), .B2(n_497), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
AND2x4_ASAP7_75t_L g510 ( .A(n_503), .B(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2x1p5_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g587 ( .A(n_507), .Y(n_587) );
AND2x4_ASAP7_75t_L g606 ( .A(n_507), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g646 ( .A(n_507), .B(n_647), .Y(n_646) );
OAI33xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_513), .A3(n_525), .B1(n_534), .B2(n_535), .B3(n_539), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x4_ASAP7_75t_L g541 ( .A(n_512), .B(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g549 ( .A(n_512), .Y(n_549) );
BUFx2_ASAP7_75t_L g556 ( .A(n_512), .Y(n_556) );
AND2x4_ASAP7_75t_L g561 ( .A(n_512), .B(n_562), .Y(n_561) );
INVx4_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx4f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g538 ( .A(n_516), .Y(n_538) );
INVx3_ASAP7_75t_L g567 ( .A(n_516), .Y(n_567) );
INVx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g524 ( .A(n_518), .Y(n_524) );
INVx2_ASAP7_75t_L g529 ( .A(n_518), .Y(n_529) );
NAND2x1_ASAP7_75t_L g533 ( .A(n_518), .B(n_519), .Y(n_533) );
AND2x2_ASAP7_75t_L g552 ( .A(n_518), .B(n_519), .Y(n_552) );
INVx1_ASAP7_75t_L g563 ( .A(n_518), .Y(n_563) );
AND2x2_ASAP7_75t_L g577 ( .A(n_518), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_519), .B(n_524), .Y(n_523) );
OR2x2_ASAP7_75t_L g528 ( .A(n_519), .B(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g557 ( .A(n_519), .Y(n_557) );
INVx2_ASAP7_75t_L g578 ( .A(n_519), .Y(n_578) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx8_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g570 ( .A(n_522), .B(n_556), .Y(n_570) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx4_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx4f_ASAP7_75t_L g545 ( .A(n_532), .Y(n_545) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OR2x6_ASAP7_75t_L g572 ( .A(n_538), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
OAI31xp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_564), .A3(n_571), .B(n_579), .Y(n_543) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVxp67_ASAP7_75t_L g566 ( .A(n_549), .Y(n_566) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_558), .B2(n_559), .Y(n_553) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
AOI32xp33_ASAP7_75t_L g595 ( .A1(n_558), .A2(n_596), .A3(n_600), .B1(n_602), .B2(n_604), .Y(n_595) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x6_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x4_ASAP7_75t_L g576 ( .A(n_573), .B(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx16_ASAP7_75t_R g575 ( .A(n_576), .Y(n_575) );
BUFx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI31xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_589), .A3(n_608), .B(n_613), .Y(n_584) );
AND2x2_ASAP7_75t_L g611 ( .A(n_587), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
AND2x2_ASAP7_75t_L g602 ( .A(n_592), .B(n_603), .Y(n_602) );
INVx3_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g596 ( .A(n_593), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x6_ASAP7_75t_L g645 ( .A(n_600), .B(n_646), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_600), .B(n_650), .C(n_653), .Y(n_649) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
CKINVDCx8_ASAP7_75t_R g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_619), .Y(n_618) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_620), .Y(n_619) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx1_ASAP7_75t_L g655 ( .A(n_622), .Y(n_655) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_624), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g669 ( .A(n_624), .B(n_655), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_640), .B1(n_656), .B2(n_657), .Y(n_625) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_626), .A2(n_656), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_632), .B2(n_633), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_633) );
INVx1_ASAP7_75t_L g639 ( .A(n_634), .Y(n_639) );
XNOR2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_636), .Y(n_634) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx12f_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx12f_ASAP7_75t_L g664 ( .A(n_642), .Y(n_664) );
BUFx8_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B(n_649), .C(n_654), .Y(n_643) );
AND2x2_ASAP7_75t_L g661 ( .A(n_644), .B(n_649), .Y(n_661) );
INVx4_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx3_ASAP7_75t_L g652 ( .A(n_648), .Y(n_652) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g660 ( .A(n_654), .Y(n_660) );
CKINVDCx14_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
BUFx3_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g665 ( .A(n_659), .Y(n_665) );
OR2x6_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
endmodule