module fake_jpeg_428_n_507 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_507);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_507;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_50),
.B(n_14),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_56),
.B(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_57),
.B(n_62),
.Y(n_123)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_58),
.Y(n_141)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_41),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g151 ( 
.A(n_64),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_67),
.Y(n_184)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_69),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_13),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_76),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_73),
.Y(n_152)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_75),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_39),
.B(n_14),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx6_ASAP7_75t_SL g78 ( 
.A(n_30),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g170 ( 
.A(n_78),
.Y(n_170)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_22),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_80),
.A2(n_94),
.B1(n_43),
.B2(n_35),
.Y(n_171)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_82),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_41),
.A2(n_0),
.B(n_1),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_30),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_84),
.Y(n_169)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_44),
.A2(n_0),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_88),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_32),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_92),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_44),
.B(n_0),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_93),
.B(n_99),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_46),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_95),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_97),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_46),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_98),
.A2(n_55),
.B1(n_43),
.B2(n_34),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_33),
.B(n_8),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_112),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_101),
.Y(n_180)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_104),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_110),
.Y(n_196)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_28),
.B(n_6),
.C(n_7),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_24),
.B(n_8),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_6),
.Y(n_178)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_47),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

CKINVDCx11_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_42),
.B1(n_21),
.B2(n_38),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g214 ( 
.A1(n_125),
.A2(n_166),
.B1(n_193),
.B2(n_195),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_67),
.B(n_6),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_148),
.B(n_202),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_60),
.B(n_34),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_153),
.B(n_159),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_122),
.A2(n_32),
.B1(n_47),
.B2(n_45),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_157),
.A2(n_164),
.B1(n_182),
.B2(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_98),
.B(n_48),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_95),
.A2(n_32),
.B1(n_45),
.B2(n_34),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_64),
.B(n_52),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_165),
.B(n_168),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_42),
.B1(n_21),
.B2(n_38),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_171),
.A2(n_173),
.B1(n_147),
.B2(n_167),
.Y(n_224)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_64),
.B(n_54),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_176),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_65),
.B(n_54),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_178),
.B(n_138),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_96),
.B(n_52),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_188),
.Y(n_232)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_101),
.B(n_48),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_85),
.Y(n_189)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_74),
.A2(n_55),
.B1(n_45),
.B2(n_25),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_L g194 ( 
.A1(n_66),
.A2(n_77),
.B1(n_70),
.B2(n_108),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_110),
.A2(n_55),
.B1(n_7),
.B2(n_8),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_65),
.B(n_82),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_151),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_92),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_104),
.A2(n_113),
.B1(n_105),
.B2(n_121),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_206),
.B1(n_125),
.B2(n_183),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_103),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_110),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_111),
.A2(n_59),
.B1(n_69),
.B2(n_81),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_209),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_210),
.Y(n_311)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_194),
.B1(n_166),
.B2(n_195),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_212),
.A2(n_224),
.B1(n_234),
.B2(n_245),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_134),
.A2(n_75),
.B1(n_68),
.B2(n_97),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_213),
.A2(n_269),
.B1(n_231),
.B2(n_230),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_215),
.B(n_219),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_145),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_216),
.Y(n_288)
);

AO22x2_ASAP7_75t_L g217 ( 
.A1(n_148),
.A2(n_75),
.B1(n_182),
.B2(n_158),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_217),
.A2(n_258),
.B1(n_274),
.B2(n_252),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_141),
.Y(n_218)
);

INVx6_ASAP7_75t_SL g282 ( 
.A(n_218),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_220),
.B(n_238),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_142),
.C(n_140),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_221),
.B(n_272),
.C(n_218),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_123),
.B(n_131),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_223),
.B(n_228),
.Y(n_325)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_152),
.Y(n_225)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_226),
.Y(n_321)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_192),
.A2(n_136),
.B1(n_143),
.B2(n_190),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_229),
.A2(n_237),
.B1(n_247),
.B2(n_271),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_139),
.B1(n_160),
.B2(n_150),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

BUFx16f_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_236),
.Y(n_292)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_152),
.Y(n_242)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_133),
.A2(n_153),
.B(n_146),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_246),
.Y(n_287)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_244),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_127),
.A2(n_160),
.B1(n_150),
.B2(n_198),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_137),
.B(n_141),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_143),
.A2(n_155),
.B1(n_205),
.B2(n_162),
.Y(n_247)
);

AO22x1_ASAP7_75t_SL g248 ( 
.A1(n_172),
.A2(n_130),
.B1(n_124),
.B2(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

INVx3_ASAP7_75t_SL g249 ( 
.A(n_156),
.Y(n_249)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_249),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_163),
.A2(n_177),
.B1(n_191),
.B2(n_187),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_250),
.A2(n_251),
.B1(n_265),
.B2(n_267),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_129),
.A2(n_180),
.B1(n_183),
.B2(n_177),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_199),
.A2(n_151),
.B(n_144),
.C(n_181),
.Y(n_252)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_252),
.A2(n_257),
.B(n_263),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_132),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_253),
.B(n_260),
.Y(n_307)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_129),
.B(n_180),
.Y(n_257)
);

AO22x1_ASAP7_75t_SL g258 ( 
.A1(n_163),
.A2(n_126),
.B1(n_135),
.B2(n_197),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_155),
.B(n_187),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_262),
.Y(n_301)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_126),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_185),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_261),
.B(n_264),
.Y(n_322)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_131),
.B(n_178),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_196),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_193),
.A2(n_88),
.B1(n_202),
.B2(n_168),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_266),
.B(n_270),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_134),
.A2(n_159),
.B1(n_133),
.B2(n_182),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_134),
.A2(n_159),
.B1(n_182),
.B2(n_161),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_170),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_206),
.A2(n_78),
.B1(n_84),
.B2(n_38),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_147),
.B(n_158),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_131),
.B(n_178),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_273),
.B(n_275),
.Y(n_319)
);

AO22x1_ASAP7_75t_SL g274 ( 
.A1(n_171),
.A2(n_164),
.B1(n_148),
.B2(n_157),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_145),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_134),
.A2(n_159),
.B1(n_133),
.B2(n_182),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_224),
.B1(n_232),
.B2(n_221),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_236),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_277),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_283),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_268),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_272),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_291),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_286),
.B(n_294),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_272),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g299 ( 
.A1(n_271),
.A2(n_274),
.B1(n_265),
.B2(n_212),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_304),
.B1(n_309),
.B2(n_312),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_210),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_300),
.B(n_313),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_208),
.B(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_314),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_274),
.A2(n_217),
.B1(n_214),
.B2(n_213),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_301),
.C(n_314),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_217),
.A2(n_214),
.B1(n_207),
.B2(n_229),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_217),
.A2(n_214),
.B1(n_247),
.B2(n_227),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_256),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_233),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_323),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_239),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_254),
.A2(n_258),
.B1(n_241),
.B2(n_240),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_279),
.B1(n_281),
.B2(n_309),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_286),
.A2(n_258),
.B1(n_235),
.B2(n_249),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_328),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_303),
.A2(n_261),
.B1(n_211),
.B2(n_248),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_303),
.A2(n_248),
.B1(n_255),
.B2(n_222),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_343),
.Y(n_363)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_302),
.A2(n_284),
.B(n_291),
.C(n_306),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_335),
.B(n_358),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_312),
.A2(n_264),
.B1(n_226),
.B2(n_253),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_336),
.A2(n_348),
.B1(n_340),
.B2(n_329),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_310),
.A2(n_244),
.B(n_260),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_337),
.A2(n_352),
.B(n_320),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_282),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_339),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_282),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_340),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_317),
.Y(n_341)
);

INVx13_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_304),
.A2(n_314),
.B1(n_294),
.B2(n_324),
.Y(n_343)
);

HAxp5_ASAP7_75t_SL g344 ( 
.A(n_287),
.B(n_280),
.CON(n_344),
.SN(n_344)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_344),
.B(n_350),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_295),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_351),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_297),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_279),
.A2(n_281),
.B1(n_326),
.B2(n_325),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_292),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_319),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_283),
.A2(n_313),
.B1(n_323),
.B2(n_322),
.Y(n_352)
);

OR2x4_ASAP7_75t_L g354 ( 
.A(n_318),
.B(n_322),
.Y(n_354)
);

OAI211xp5_ASAP7_75t_SL g370 ( 
.A1(n_354),
.A2(n_296),
.B(n_308),
.C(n_285),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_316),
.A2(n_296),
.B1(n_293),
.B2(n_322),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_297),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_292),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_356),
.B(n_307),
.Y(n_371)
);

INVx5_ASAP7_75t_SL g357 ( 
.A(n_277),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_357),
.Y(n_360)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_346),
.A2(n_278),
.B(n_307),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_368),
.A2(n_370),
.B(n_337),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_376),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_341),
.B(n_307),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_372),
.B(n_382),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_331),
.Y(n_373)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_373),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_374),
.A2(n_343),
.B1(n_327),
.B2(n_349),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_375),
.A2(n_377),
.B(n_352),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_329),
.A2(n_315),
.B1(n_289),
.B2(n_290),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_349),
.A2(n_311),
.B(n_298),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_383),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_381),
.B(n_342),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_351),
.B(n_290),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_321),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_359),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_384),
.Y(n_401)
);

AND2x2_ASAP7_75t_SL g385 ( 
.A(n_349),
.B(n_311),
.Y(n_385)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_385),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_378),
.Y(n_386)
);

BUFx2_ASAP7_75t_SL g423 ( 
.A(n_386),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_388),
.A2(n_404),
.B1(n_362),
.B2(n_394),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_378),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_390),
.B(n_410),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_393),
.A2(n_412),
.B(n_377),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_394),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_367),
.A2(n_348),
.B1(n_334),
.B2(n_347),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_396),
.A2(n_399),
.B1(n_407),
.B2(n_365),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_356),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_397),
.B(n_384),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_383),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_367),
.A2(n_354),
.B1(n_335),
.B2(n_336),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_345),
.Y(n_400)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_400),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_353),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_402),
.B(n_405),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_355),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_385),
.C(n_380),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_373),
.A2(n_339),
.B1(n_338),
.B2(n_332),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_358),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_363),
.A2(n_328),
.B1(n_330),
.B2(n_333),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_408),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_368),
.A2(n_350),
.B(n_357),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_409),
.A2(n_375),
.B(n_377),
.Y(n_414)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_411),
.B(n_365),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_375),
.A2(n_357),
.B(n_298),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_414),
.A2(n_421),
.B(n_389),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_391),
.B(n_372),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_420),
.B(n_431),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_399),
.A2(n_374),
.B1(n_363),
.B2(n_366),
.Y(n_421)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_424),
.B(n_392),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_402),
.B(n_385),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_427),
.B(n_429),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_428),
.B(n_393),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_398),
.B(n_385),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_430),
.B(n_407),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_288),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_371),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_432),
.B(n_390),
.C(n_386),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_401),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_435),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_442),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_396),
.C(n_395),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_441),
.C(n_443),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_395),
.C(n_412),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_405),
.C(n_409),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_452),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_446),
.A2(n_428),
.B(n_387),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_430),
.B(n_388),
.C(n_389),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_424),
.C(n_414),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_427),
.B(n_387),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_448),
.B(n_417),
.Y(n_454)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_416),
.Y(n_450)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_450),
.Y(n_455)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_416),
.Y(n_453)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_453),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_454),
.B(n_457),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_451),
.A2(n_421),
.B1(n_415),
.B2(n_413),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_456),
.B(n_459),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_444),
.B(n_449),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_436),
.A2(n_413),
.B1(n_423),
.B2(n_425),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_463),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_439),
.A2(n_425),
.B1(n_376),
.B2(n_362),
.Y(n_461)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_462),
.B(n_467),
.Y(n_471)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_441),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_459),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_473),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_462),
.B(n_447),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_464),
.B(n_466),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_474),
.B(n_475),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_445),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_438),
.C(n_443),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_476),
.B(n_477),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_458),
.B(n_440),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_477),
.B(n_460),
.C(n_465),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_481),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_468),
.B(n_455),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_469),
.B(n_465),
.C(n_456),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_487),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_484),
.B(n_486),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_463),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_376),
.B1(n_433),
.B2(n_426),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_476),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_488),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_478),
.C(n_442),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_489),
.B(n_491),
.C(n_452),
.Y(n_498)
);

XOR2x2_ASAP7_75t_L g490 ( 
.A(n_482),
.B(n_478),
.Y(n_490)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_490),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_483),
.B(n_440),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_494),
.B(n_485),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_497),
.Y(n_500)
);

AOI31xp67_ASAP7_75t_L g497 ( 
.A1(n_490),
.A2(n_379),
.A3(n_433),
.B(n_426),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_493),
.Y(n_501)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_501),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_495),
.B(n_492),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_492),
.B(n_499),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_503),
.B(n_500),
.C(n_360),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_505),
.A2(n_504),
.B(n_360),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_410),
.Y(n_507)
);


endmodule