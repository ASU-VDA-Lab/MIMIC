module fake_jpeg_27739_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_15),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_44),
.Y(n_47)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_52),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_71),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_17),
.B1(n_32),
.B2(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_36),
.B1(n_29),
.B2(n_38),
.Y(n_86)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_68),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_17),
.B(n_33),
.Y(n_79)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_29),
.A3(n_23),
.B1(n_32),
.B2(n_21),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_23),
.C(n_21),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_32),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_17),
.B1(n_45),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_84),
.B1(n_66),
.B2(n_70),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_17),
.B1(n_45),
.B2(n_19),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_25),
.B(n_33),
.C(n_20),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_29),
.B1(n_23),
.B2(n_25),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_53),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_97),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_36),
.B1(n_16),
.B2(n_32),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_72),
.B1(n_67),
.B2(n_62),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_57),
.B1(n_73),
.B2(n_62),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_29),
.B1(n_24),
.B2(n_31),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_98),
.A2(n_94),
.B1(n_93),
.B2(n_90),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_101),
.Y(n_139)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_49),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_97),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_105),
.Y(n_134)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_121),
.B(n_124),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_113),
.Y(n_141)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_118),
.B1(n_116),
.B2(n_124),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_20),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_112),
.B(n_122),
.Y(n_136)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_88),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_69),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_117),
.Y(n_146)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_15),
.C(n_1),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_16),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g124 ( 
.A(n_82),
.B(n_59),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_76),
.B(n_95),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_103),
.B1(n_119),
.B2(n_107),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_126),
.A2(n_132),
.B1(n_143),
.B2(n_150),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_111),
.B1(n_93),
.B2(n_109),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_19),
.B(n_20),
.Y(n_182)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_144),
.B(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_75),
.C(n_77),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_151),
.C(n_121),
.Y(n_161)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_154),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_94),
.B1(n_80),
.B2(n_76),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_148),
.A2(n_105),
.B1(n_93),
.B2(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_94),
.B1(n_64),
.B2(n_80),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_85),
.C(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_140),
.Y(n_176)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_166),
.B1(n_170),
.B2(n_132),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_157),
.B(n_178),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_137),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_182),
.B1(n_183),
.B2(n_147),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_112),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_165),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_162),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_169),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_121),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g167 ( 
.A(n_129),
.B(n_111),
.C(n_85),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_167),
.A2(n_154),
.B1(n_128),
.B2(n_26),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_111),
.C(n_100),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_165),
.C(n_161),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_79),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_90),
.B1(n_78),
.B2(n_113),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_90),
.B1(n_108),
.B2(n_117),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_173),
.B1(n_177),
.B2(n_148),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_46),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_152),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_59),
.B1(n_54),
.B2(n_50),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_50),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_21),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_143),
.A2(n_54),
.B1(n_33),
.B2(n_24),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_136),
.B(n_149),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_32),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_146),
.B(n_131),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_184),
.A2(n_210),
.B(n_182),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_186),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_23),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_199),
.B1(n_208),
.B2(n_157),
.Y(n_214)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_192),
.B(n_202),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_155),
.A2(n_130),
.B1(n_141),
.B2(n_131),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_201),
.B1(n_203),
.B2(n_205),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_23),
.C(n_21),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_139),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_155),
.A2(n_130),
.B1(n_144),
.B2(n_143),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_153),
.B1(n_150),
.B2(n_134),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_136),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_135),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_172),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_135),
.B1(n_137),
.B2(n_31),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_173),
.A2(n_19),
.B1(n_26),
.B2(n_25),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_156),
.B1(n_170),
.B2(n_163),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_216),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_224),
.B1(n_186),
.B2(n_193),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_232),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_219),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_181),
.Y(n_218)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_167),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_183),
.B1(n_158),
.B2(n_24),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_158),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_226),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_185),
.A2(n_26),
.B1(n_22),
.B2(n_27),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_27),
.Y(n_223)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_188),
.B(n_22),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_27),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_27),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_194),
.C(n_206),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_198),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_21),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_192),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_203),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_201),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_247),
.B1(n_213),
.B2(n_215),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_250),
.C(n_253),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_2),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_194),
.C(n_189),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_231),
.A2(n_191),
.B1(n_184),
.B2(n_204),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_259),
.B1(n_224),
.B2(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_200),
.C(n_210),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_209),
.C(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_256),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_0),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_229),
.C(n_226),
.Y(n_256)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_223),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_213),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_262),
.B1(n_269),
.B2(n_275),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_252),
.B1(n_249),
.B2(n_239),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_258),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_263),
.B(n_272),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_219),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_267),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_211),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_266),
.B(n_257),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_268),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_236),
.B1(n_218),
.B2(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_243),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_254),
.Y(n_285)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_245),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_251),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_276),
.B(n_237),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_241),
.Y(n_277)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_241),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_242),
.C(n_256),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_291),
.C(n_264),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_248),
.B(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_5),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_286),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g288 ( 
.A(n_271),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_285),
.B1(n_291),
.B2(n_292),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_237),
.C(n_253),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_297),
.C(n_302),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_262),
.C(n_265),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_283),
.B(n_273),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_260),
.B(n_266),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_299),
.A2(n_303),
.B(n_306),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_306),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_278),
.B1(n_269),
.B2(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_304),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_14),
.C(n_6),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_293),
.A2(n_289),
.B(n_287),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_5),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_5),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_297),
.C(n_296),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_313),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_299),
.A2(n_290),
.B1(n_9),
.B2(n_10),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_8),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_317),
.B(n_11),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_300),
.B(n_10),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_318),
.B(n_320),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_9),
.B(n_10),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_9),
.B(n_10),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_321),
.A2(n_11),
.B(n_12),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_9),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_314),
.B(n_308),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_327),
.A2(n_329),
.B(n_330),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_310),
.B(n_12),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_326),
.A2(n_325),
.B(n_319),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_328),
.B(n_12),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_331),
.C(n_13),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_11),
.B(n_13),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_14),
.Y(n_337)
);


endmodule