module fake_aes_4835_n_487 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_487);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_487;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g72 ( .A(n_59), .Y(n_72) );
INVxp33_ASAP7_75t_L g73 ( .A(n_63), .Y(n_73) );
INVx2_ASAP7_75t_L g74 ( .A(n_0), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_28), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_47), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_36), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_62), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_40), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_20), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_4), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_16), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_2), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_27), .Y(n_87) );
NOR2xp67_ASAP7_75t_L g88 ( .A(n_0), .B(n_38), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_9), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_57), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_56), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_8), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_10), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_70), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_43), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_9), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_58), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_32), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_41), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_69), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_66), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_26), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_52), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_55), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_50), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_29), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_14), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_101), .Y(n_112) );
NOR2xp67_ASAP7_75t_L g113 ( .A(n_91), .B(n_1), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_87), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_87), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_77), .Y(n_117) );
OAI21x1_ASAP7_75t_L g118 ( .A1(n_78), .A2(n_30), .B(n_68), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_78), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_90), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_90), .Y(n_123) );
CKINVDCx11_ASAP7_75t_R g124 ( .A(n_86), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_107), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_73), .B(n_1), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_97), .B(n_2), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_107), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_98), .B(n_3), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_100), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_111), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_116), .B(n_74), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_119), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_119), .Y(n_138) );
OR2x2_ASAP7_75t_L g139 ( .A(n_128), .B(n_83), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_119), .Y(n_140) );
NAND2x1p5_ASAP7_75t_L g141 ( .A(n_116), .B(n_81), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_132), .B(n_100), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g144 ( .A(n_127), .B(n_92), .C(n_83), .Y(n_144) );
HB1xp67_ASAP7_75t_L g145 ( .A(n_115), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_119), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_119), .Y(n_147) );
INVx4_ASAP7_75t_L g148 ( .A(n_133), .Y(n_148) );
OAI22xp33_ASAP7_75t_L g149 ( .A1(n_112), .A2(n_93), .B1(n_89), .B2(n_82), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_133), .Y(n_151) );
CKINVDCx16_ASAP7_75t_R g152 ( .A(n_127), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_118), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_117), .B(n_74), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_133), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
NAND3xp33_ASAP7_75t_L g158 ( .A(n_120), .B(n_110), .C(n_109), .Y(n_158) );
INVx6_ASAP7_75t_L g159 ( .A(n_127), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_120), .B(n_109), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_141), .B(n_121), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_144), .B(n_128), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_157), .A2(n_126), .B(n_131), .C(n_121), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g165 ( .A1(n_152), .A2(n_134), .B1(n_124), .B2(n_123), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_159), .B(n_122), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_145), .Y(n_167) );
INVx4_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_152), .B(n_128), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_136), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_159), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_141), .B(n_126), .Y(n_173) );
OAI22xp33_ASAP7_75t_L g174 ( .A1(n_159), .A2(n_129), .B1(n_125), .B2(n_134), .Y(n_174) );
OR2x2_ASAP7_75t_SL g175 ( .A(n_139), .B(n_124), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_159), .A2(n_131), .B1(n_130), .B2(n_106), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_139), .B(n_113), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_151), .A2(n_118), .B(n_130), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_156), .Y(n_181) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_141), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_160), .B(n_106), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_137), .Y(n_189) );
NOR2xp33_ASAP7_75t_R g190 ( .A(n_143), .B(n_84), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_135), .Y(n_191) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_135), .Y(n_192) );
NAND2xp33_ASAP7_75t_SL g193 ( .A(n_153), .B(n_84), .Y(n_193) );
OR2x2_ASAP7_75t_L g194 ( .A(n_169), .B(n_149), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_182), .A2(n_158), .B1(n_135), .B2(n_154), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_169), .B(n_135), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_187), .B(n_154), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_161), .A2(n_158), .B1(n_154), .B2(n_113), .Y(n_198) );
AOI221xp5_ASAP7_75t_L g199 ( .A1(n_174), .A2(n_154), .B1(n_155), .B2(n_153), .C(n_85), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_161), .A2(n_153), .B1(n_155), .B2(n_85), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_167), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_187), .B(n_153), .Y(n_202) );
BUFx3_ASAP7_75t_L g203 ( .A(n_187), .Y(n_203) );
AOI222xp33_ASAP7_75t_L g204 ( .A1(n_165), .A2(n_88), .B1(n_110), .B2(n_72), .C1(n_103), .C2(n_75), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_184), .Y(n_205) );
BUFx3_ASAP7_75t_L g206 ( .A(n_188), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_185), .B(n_155), .Y(n_208) );
AOI221xp5_ASAP7_75t_L g209 ( .A1(n_162), .A2(n_155), .B1(n_108), .B2(n_105), .C(n_94), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_184), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_162), .B(n_155), .Y(n_211) );
NAND2xp33_ASAP7_75t_L g212 ( .A(n_173), .B(n_136), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_176), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_184), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_188), .B(n_76), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_184), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_162), .B(n_95), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_173), .B(n_96), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_185), .B(n_99), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_177), .B(n_102), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_188), .Y(n_221) );
BUFx4_ASAP7_75t_SL g222 ( .A(n_189), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_165), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_184), .Y(n_224) );
OAI21xp33_ASAP7_75t_L g225 ( .A1(n_186), .A2(n_150), .B(n_147), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_168), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_207), .Y(n_228) );
INVx6_ASAP7_75t_SL g229 ( .A(n_221), .Y(n_229) );
OAI21xp33_ASAP7_75t_L g230 ( .A1(n_217), .A2(n_190), .B(n_177), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_208), .A2(n_184), .B(n_180), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_196), .B(n_162), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_226), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_207), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_196), .B(n_186), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_213), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_216), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_203), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_194), .B(n_175), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_218), .A2(n_163), .B1(n_191), .B2(n_192), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_197), .B(n_179), .Y(n_242) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_201), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_203), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_216), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_221), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_197), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_203), .B(n_191), .Y(n_248) );
AND2x2_ASAP7_75t_SL g249 ( .A(n_216), .B(n_168), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_220), .B(n_179), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_194), .B(n_179), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g252 ( .A1(n_219), .A2(n_179), .B1(n_191), .B2(n_166), .C(n_172), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_211), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_206), .B(n_191), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_230), .A2(n_204), .B1(n_199), .B2(n_223), .Y(n_256) );
AOI222xp33_ASAP7_75t_L g257 ( .A1(n_251), .A2(n_209), .B1(n_215), .B2(n_175), .C1(n_195), .C2(n_218), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_228), .B(n_215), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_230), .A2(n_204), .B1(n_195), .B2(n_198), .Y(n_259) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_231), .A2(n_200), .B(n_198), .Y(n_260) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_240), .A2(n_172), .B1(n_206), .B2(n_227), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_228), .B(n_206), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_240), .A2(n_227), .B1(n_226), .B2(n_183), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_246), .Y(n_264) );
OAI22xp33_ASAP7_75t_L g265 ( .A1(n_241), .A2(n_200), .B1(n_226), .B2(n_227), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_234), .B(n_226), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_234), .Y(n_267) );
NAND2x1_ASAP7_75t_L g268 ( .A(n_238), .B(n_216), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_241), .A2(n_216), .B1(n_227), .B2(n_224), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_243), .Y(n_270) );
AOI22xp33_ASAP7_75t_SL g271 ( .A1(n_249), .A2(n_222), .B1(n_104), .B2(n_212), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_236), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_236), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_249), .Y(n_274) );
OAI211xp5_ASAP7_75t_L g275 ( .A1(n_252), .A2(n_250), .B(n_254), .C(n_237), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_237), .B(n_183), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_232), .B(n_168), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_232), .B(n_171), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_249), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_257), .A2(n_256), .B1(n_259), .B2(n_261), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_272), .B(n_254), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_259), .A2(n_247), .B1(n_242), .B2(n_235), .C(n_248), .Y(n_283) );
AOI33xp33_ASAP7_75t_L g284 ( .A1(n_256), .A2(n_263), .A3(n_261), .B1(n_271), .B2(n_247), .B3(n_265), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_272), .Y(n_285) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_257), .A2(n_202), .B(n_193), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_271), .A2(n_242), .B1(n_255), .B2(n_248), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g288 ( .A1(n_265), .A2(n_235), .B1(n_248), .B2(n_255), .C(n_233), .Y(n_288) );
OAI33xp33_ASAP7_75t_L g289 ( .A1(n_267), .A2(n_142), .A3(n_147), .B1(n_150), .B2(n_146), .B3(n_140), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_267), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_273), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_264), .B(n_246), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_273), .Y(n_293) );
AO21x1_ASAP7_75t_SL g294 ( .A1(n_279), .A2(n_229), .B(n_225), .Y(n_294) );
NOR2xp33_ASAP7_75t_R g295 ( .A(n_270), .B(n_239), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_274), .B(n_233), .Y(n_296) );
AND2x6_ASAP7_75t_L g297 ( .A(n_274), .B(n_238), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_263), .A2(n_229), .B1(n_244), .B2(n_239), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_274), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_258), .B(n_248), .Y(n_300) );
CKINVDCx16_ASAP7_75t_R g301 ( .A(n_279), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_297), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_282), .B(n_260), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_297), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_290), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_285), .B(n_260), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_280), .B(n_275), .C(n_269), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_301), .B(n_285), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_285), .B(n_260), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_287), .A2(n_258), .B1(n_277), .B2(n_278), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_258), .B1(n_275), .B2(n_276), .C1(n_266), .C2(n_278), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_286), .A2(n_269), .B(n_260), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_291), .Y(n_317) );
OAI21xp33_ASAP7_75t_SL g318 ( .A1(n_284), .A2(n_291), .B(n_293), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_281), .B(n_276), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_288), .A2(n_278), .B1(n_277), .B2(n_255), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_281), .B(n_276), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_299), .B(n_266), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_300), .A2(n_277), .B1(n_266), .B2(n_262), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_297), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
OAI31xp33_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_262), .A3(n_255), .B(n_233), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_297), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_301), .B(n_268), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_329), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_319), .B(n_292), .Y(n_331) );
NAND4xp25_ASAP7_75t_L g332 ( .A(n_315), .B(n_296), .C(n_233), .D(n_142), .Y(n_332) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_329), .B(n_297), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_319), .B(n_299), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_317), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_321), .B(n_296), .Y(n_336) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_307), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_307), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_328), .B(n_297), .Y(n_339) );
NAND2xp33_ASAP7_75t_SL g340 ( .A(n_306), .B(n_295), .Y(n_340) );
NAND2xp33_ASAP7_75t_R g341 ( .A(n_328), .B(n_294), .Y(n_341) );
NAND4xp25_ASAP7_75t_L g342 ( .A(n_315), .B(n_296), .C(n_4), .D(n_5), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_317), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_326), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_302), .Y(n_345) );
NAND2x2_ASAP7_75t_L g346 ( .A(n_303), .B(n_294), .Y(n_346) );
OAI33xp33_ASAP7_75t_L g347 ( .A1(n_310), .A2(n_3), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_347) );
OR2x2_ASAP7_75t_L g348 ( .A(n_321), .B(n_296), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_324), .B(n_6), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_304), .B(n_7), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_302), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_327), .B(n_253), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_318), .B(n_289), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_328), .B(n_268), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_311), .B(n_10), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_311), .B(n_329), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_304), .B(n_11), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_327), .B(n_253), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_328), .B(n_253), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_308), .B(n_12), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_303), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_310), .B(n_12), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_324), .B(n_13), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_313), .Y(n_364) );
INVxp33_ASAP7_75t_L g365 ( .A(n_303), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_313), .B(n_13), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_314), .B1(n_320), .B2(n_306), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_356), .B(n_312), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_342), .B(n_323), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_350), .B(n_312), .Y(n_370) );
OAI32xp33_ASAP7_75t_L g371 ( .A1(n_340), .A2(n_325), .A3(n_322), .B1(n_306), .B2(n_323), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_337), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_334), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
OAI22xp33_ASAP7_75t_SL g378 ( .A1(n_346), .A2(n_322), .B1(n_325), .B2(n_317), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_L g379 ( .A1(n_362), .A2(n_305), .B(n_312), .C(n_309), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_332), .A2(n_309), .B1(n_304), .B2(n_316), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_362), .A2(n_316), .B1(n_305), .B2(n_136), .C(n_146), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_344), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_335), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_345), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_330), .Y(n_386) );
NAND2xp33_ASAP7_75t_SL g387 ( .A(n_341), .B(n_316), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_364), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_347), .A2(n_245), .B1(n_238), .B2(n_205), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_353), .B(n_136), .C(n_138), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_333), .A2(n_229), .B1(n_245), .B2(n_15), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_SL g392 ( .A1(n_355), .A2(n_17), .B(n_229), .C(n_245), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_349), .A2(n_224), .B1(n_214), .B2(n_210), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_357), .B(n_140), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_331), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_352), .A2(n_214), .B(n_210), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_348), .B(n_18), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_363), .A2(n_366), .B1(n_360), .B2(n_357), .C(n_336), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_343), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_352), .A2(n_205), .B(n_225), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_365), .B(n_19), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_365), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_181), .B1(n_178), .B2(n_171), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_358), .A2(n_138), .B(n_171), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_359), .B(n_21), .Y(n_406) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_375), .B(n_339), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_369), .B(n_354), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_368), .B(n_339), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_382), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
AOI221x1_ASAP7_75t_SL g412 ( .A1(n_369), .A2(n_354), .B1(n_359), .B2(n_341), .C(n_33), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_403), .B(n_395), .Y(n_414) );
NOR4xp25_ASAP7_75t_SL g415 ( .A(n_376), .B(n_354), .C(n_25), .D(n_31), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_386), .B(n_23), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_372), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_388), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_372), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_402), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_370), .B(n_35), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_373), .B(n_37), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_397), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_398), .B(n_42), .Y(n_425) );
XNOR2xp5_ASAP7_75t_L g426 ( .A(n_367), .B(n_44), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_374), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_383), .Y(n_428) );
XNOR2x1_ASAP7_75t_L g429 ( .A(n_380), .B(n_45), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g431 ( .A1(n_378), .A2(n_46), .B(n_48), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_379), .B(n_49), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
NAND2xp33_ASAP7_75t_SL g435 ( .A(n_404), .B(n_51), .Y(n_435) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_390), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g437 ( .A1(n_391), .A2(n_53), .B(n_54), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_381), .B(n_61), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g439 ( .A1(n_408), .A2(n_391), .B1(n_387), .B2(n_401), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g440 ( .A(n_413), .B(n_405), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_413), .B(n_400), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_414), .B(n_393), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_417), .B(n_400), .Y(n_443) );
OAI322xp33_ASAP7_75t_L g444 ( .A1(n_408), .A2(n_406), .A3(n_389), .B1(n_396), .B2(n_392), .C1(n_371), .C2(n_404), .Y(n_444) );
XNOR2xp5_ASAP7_75t_L g445 ( .A(n_407), .B(n_64), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_429), .B(n_178), .C(n_181), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g447 ( .A(n_412), .B(n_164), .C(n_170), .D(n_71), .Y(n_447) );
NAND3xp33_ASAP7_75t_L g448 ( .A(n_429), .B(n_170), .C(n_425), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_411), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_418), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_410), .B(n_434), .Y(n_452) );
BUFx3_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_428), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_430), .A2(n_424), .B1(n_426), .B2(n_437), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_436), .Y(n_456) );
O2A1O1Ixp5_ASAP7_75t_L g457 ( .A1(n_435), .A2(n_431), .B(n_432), .C(n_423), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_427), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_458), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_452), .Y(n_460) );
NOR2xp67_ASAP7_75t_L g461 ( .A(n_447), .B(n_409), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_453), .Y(n_462) );
OAI21xp33_ASAP7_75t_L g463 ( .A1(n_439), .A2(n_422), .B(n_433), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_440), .A2(n_415), .B(n_438), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_457), .A2(n_455), .B(n_440), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_445), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_446), .A2(n_441), .B(n_448), .C(n_442), .Y(n_467) );
AOI211x1_ASAP7_75t_L g468 ( .A1(n_441), .A2(n_449), .B(n_451), .C(n_450), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_454), .B(n_457), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_443), .B(n_420), .Y(n_470) );
NOR4xp25_ASAP7_75t_L g471 ( .A(n_456), .B(n_447), .C(n_444), .D(n_421), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_456), .A2(n_444), .B1(n_412), .B2(n_408), .C(n_452), .Y(n_472) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_455), .A2(n_447), .B(n_439), .C(n_456), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g474 ( .A1(n_473), .A2(n_465), .B1(n_467), .B2(n_469), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_460), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_470), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_466), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_459), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_474), .B(n_472), .C(n_464), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_478), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_476), .A2(n_468), .B1(n_462), .B2(n_461), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_480), .Y(n_482) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_479), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_482), .Y(n_484) );
INVxp67_ASAP7_75t_L g485 ( .A(n_483), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_485), .A2(n_481), .B1(n_477), .B2(n_475), .Y(n_486) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_486), .A2(n_484), .B1(n_471), .B2(n_477), .C(n_463), .Y(n_487) );
endmodule