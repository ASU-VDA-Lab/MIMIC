module fake_jpeg_9255_n_312 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_312);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_312;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_33),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_46),
.A2(n_55),
.B1(n_21),
.B2(n_23),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_47),
.B(n_57),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_22),
.B(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_24),
.B1(n_22),
.B2(n_16),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_21),
.B1(n_16),
.B2(n_28),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_30),
.C(n_28),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_29),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_67),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_68),
.Y(n_82)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_27),
.B1(n_16),
.B2(n_21),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_67),
.B1(n_62),
.B2(n_44),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_53),
.B1(n_69),
.B2(n_65),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_80),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_21),
.B1(n_42),
.B2(n_39),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_61),
.B1(n_44),
.B2(n_41),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_79),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_83),
.A2(n_23),
.B1(n_42),
.B2(n_44),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_57),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_25),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_54),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_30),
.B1(n_25),
.B2(n_39),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_30),
.B1(n_17),
.B2(n_29),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_80),
.B(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_104),
.Y(n_131)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_103),
.Y(n_144)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_56),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_105),
.B(n_115),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_107),
.A2(n_109),
.B(n_74),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_108),
.B(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_110),
.A2(n_111),
.B1(n_122),
.B2(n_82),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_62),
.B1(n_53),
.B2(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_45),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_113),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_45),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_110),
.B(n_111),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_120),
.Y(n_150)
);

O2A1O1Ixp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_26),
.B(n_31),
.C(n_20),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_84),
.B(n_77),
.C(n_72),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_63),
.Y(n_121)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_84),
.A2(n_41),
.B1(n_18),
.B2(n_31),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_130),
.Y(n_165)
);

XNOR2x2_ASAP7_75t_SL g173 ( 
.A(n_128),
.B(n_26),
.Y(n_173)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_92),
.C(n_76),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_133),
.C(n_143),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_95),
.C(n_93),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_102),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g135 ( 
.A1(n_123),
.A2(n_73),
.B(n_94),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_33),
.B(n_32),
.Y(n_175)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_136),
.B(n_138),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_78),
.B1(n_73),
.B2(n_87),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_117),
.B1(n_99),
.B2(n_82),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_95),
.C(n_90),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_148),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_116),
.B(n_106),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_74),
.C(n_96),
.Y(n_143)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_26),
.C(n_32),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_108),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_17),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_124),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_100),
.B(n_113),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_119),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_114),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_130),
.C(n_132),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_120),
.Y(n_156)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_156),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_149),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_173),
.B(n_175),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_162),
.B(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_163),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_107),
.B1(n_99),
.B2(n_124),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_175),
.B1(n_167),
.B2(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_115),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_125),
.B1(n_97),
.B2(n_96),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_103),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_174),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_180),
.C(n_184),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_135),
.B(n_147),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_177),
.A2(n_182),
.B(n_189),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_137),
.C(n_133),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_142),
.B1(n_126),
.B2(n_136),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_162),
.B1(n_170),
.B2(n_173),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_137),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_142),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_188),
.C(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_187),
.B(n_192),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_145),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_126),
.B(n_148),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_145),
.B(n_146),
.Y(n_193)
);

NOR4xp25_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_11),
.C(n_15),
.D(n_14),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_141),
.C(n_138),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_171),
.B1(n_82),
.B2(n_68),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_97),
.Y(n_205)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_160),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_156),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_188),
.C(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_210),
.Y(n_238)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_207),
.B(n_178),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_153),
.Y(n_209)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_221),
.B(n_222),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_213),
.C(n_180),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_166),
.C(n_173),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_154),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_33),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_171),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_219),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_217),
.A2(n_183),
.B1(n_191),
.B2(n_192),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_12),
.C(n_9),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_10),
.B(n_15),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_177),
.B(n_10),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_10),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_223),
.A2(n_195),
.B(n_197),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_235),
.B1(n_236),
.B2(n_215),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_222),
.B1(n_211),
.B2(n_221),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_194),
.B1(n_178),
.B2(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_R g244 ( 
.A(n_232),
.B(n_220),
.C(n_7),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_184),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_234),
.C(n_237),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_177),
.B1(n_68),
.B2(n_60),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_202),
.B(n_60),
.C(n_33),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_206),
.C(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_60),
.C(n_33),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_32),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_247),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_236),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_204),
.B(n_203),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_6),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_31),
.B1(n_20),
.B2(n_18),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_252),
.A2(n_239),
.B1(n_227),
.B2(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_214),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_256),
.C(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_203),
.C(n_217),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_224),
.A2(n_8),
.B(n_13),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_33),
.C(n_32),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_32),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_20),
.C(n_1),
.Y(n_273)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_253),
.A2(n_238),
.B1(n_243),
.B2(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_264),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_240),
.B1(n_232),
.B2(n_31),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_273),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_269),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_267),
.B(n_20),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_5),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_258),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_255),
.C(n_245),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_0),
.C(n_1),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_268),
.B1(n_264),
.B2(n_265),
.Y(n_286)
);

NOR2xp67_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_255),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_254),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_268),
.B(n_245),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_285),
.B(n_275),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_4),
.CI(n_8),
.CON(n_285),
.SN(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_286),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_261),
.B(n_273),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_4),
.B(n_6),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_4),
.C(n_6),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_299),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_281),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_296),
.A2(n_2),
.B(n_3),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_279),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_300),
.A2(n_302),
.B(n_9),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_5),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_307),
.Y(n_309)
);

O2A1O1Ixp33_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_1),
.C(n_2),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_309),
.B(n_296),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_304),
.B(n_308),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_301),
.Y(n_312)
);


endmodule