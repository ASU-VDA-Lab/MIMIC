module fake_jpeg_11837_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_6),
.B(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_1),
.B(n_7),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_16),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_14),
.B(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_15),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_10),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_21),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_32),
.B(n_33),
.Y(n_41)
);

AOI21x1_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_22),
.B(n_19),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_11),
.B1(n_8),
.B2(n_20),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.C(n_32),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_9),
.C(n_30),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.C(n_8),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_50),
.A2(n_51),
.B1(n_11),
.B2(n_20),
.Y(n_52)
);

AOI321xp33_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_49),
.A3(n_20),
.B1(n_15),
.B2(n_46),
.C(n_5),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_15),
.C(n_1),
.Y(n_54)
);


endmodule