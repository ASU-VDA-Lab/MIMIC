module fake_jpeg_1215_n_268 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_9),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_0),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_45),
.Y(n_82)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_43),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_21),
.B(n_0),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_32),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_69),
.Y(n_88)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_62),
.Y(n_83)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_64),
.Y(n_87)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_75),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_32),
.B(n_1),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_67),
.Y(n_96)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_16),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_70),
.B(n_29),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_74),
.C(n_76),
.Y(n_91)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_16),
.B(n_2),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_79),
.Y(n_105)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_25),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_41),
.B1(n_40),
.B2(n_22),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_86),
.A2(n_103),
.B1(n_123),
.B2(n_64),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_89),
.B(n_100),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_43),
.A2(n_27),
.B1(n_23),
.B2(n_36),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_99),
.B1(n_104),
.B2(n_116),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_34),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_111),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_48),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_122),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_22),
.B1(n_25),
.B2(n_19),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_54),
.A2(n_25),
.B1(n_19),
.B2(n_6),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_3),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_71),
.B(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_3),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_4),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_57),
.A2(n_19),
.B1(n_8),
.B2(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_128),
.B(n_135),
.Y(n_169)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_144),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_101),
.A2(n_63),
.B1(n_67),
.B2(n_58),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_111),
.B1(n_114),
.B2(n_106),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_8),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_155),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_149),
.B1(n_152),
.B2(n_158),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_78),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_92),
.Y(n_145)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_82),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_114),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_98),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_156),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_84),
.B(n_8),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_89),
.B(n_88),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_159),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_83),
.A2(n_12),
.B1(n_19),
.B2(n_87),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_90),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_160),
.A2(n_115),
.B1(n_90),
.B2(n_118),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_110),
.B(n_100),
.C(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_165),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_83),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_168),
.A2(n_183),
.B1(n_114),
.B2(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_83),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_187),
.B1(n_188),
.B2(n_160),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_95),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_132),
.B(n_95),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_150),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_139),
.A2(n_95),
.B1(n_106),
.B2(n_112),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_125),
.B1(n_127),
.B2(n_140),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_131),
.A2(n_106),
.B1(n_112),
.B2(n_118),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_143),
.B1(n_134),
.B2(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_187),
.A2(n_131),
.B1(n_129),
.B2(n_144),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_192),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_137),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_138),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_195),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_149),
.C(n_91),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_197),
.B1(n_208),
.B2(n_209),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_159),
.B1(n_153),
.B2(n_130),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_175),
.B(n_165),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_198),
.A2(n_172),
.B(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_167),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_178),
.A2(n_112),
.B1(n_118),
.B2(n_152),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_174),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_207),
.A2(n_185),
.B1(n_145),
.B2(n_152),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_185),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_162),
.C(n_179),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_219),
.C(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_196),
.A2(n_183),
.B1(n_172),
.B2(n_174),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_205),
.B1(n_203),
.B2(n_200),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_209),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_170),
.B(n_186),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_216),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_186),
.B(n_176),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_224),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_182),
.C(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_181),
.C(n_184),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_223),
.A2(n_201),
.B1(n_189),
.B2(n_195),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_229),
.A2(n_237),
.B1(n_210),
.B2(n_217),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_215),
.A2(n_201),
.B1(n_204),
.B2(n_207),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_230),
.A2(n_215),
.B1(n_222),
.B2(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_219),
.B1(n_188),
.B2(n_214),
.Y(n_241)
);

AO221x1_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_149),
.B1(n_206),
.B2(n_115),
.C(n_136),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_233),
.B(n_234),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_199),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_182),
.C(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_224),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_238),
.B(n_189),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_231),
.A3(n_237),
.B(n_236),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_242),
.B1(n_228),
.B2(n_235),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_227),
.A2(n_220),
.B1(n_218),
.B2(n_216),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_236),
.C(n_220),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_248),
.B1(n_243),
.B2(n_244),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_228),
.B(n_230),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_250),
.A2(n_245),
.B(n_238),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_246),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_252),
.A2(n_243),
.B1(n_164),
.B2(n_115),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_253),
.B(n_255),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_245),
.C(n_241),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_257),
.B(n_252),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_249),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_258),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_259),
.B(n_255),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_261),
.B(n_254),
.Y(n_264)
);

BUFx24_ASAP7_75t_SL g265 ( 
.A(n_264),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_266),
.A2(n_262),
.B(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_265),
.Y(n_268)
);


endmodule