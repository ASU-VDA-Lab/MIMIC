module real_aes_8404_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_729;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g514 ( .A(n_1), .Y(n_514) );
INVx1_ASAP7_75t_L g195 ( .A(n_2), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_3), .A2(n_38), .B1(n_157), .B2(n_456), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_4), .Y(n_753) );
AOI21xp33_ASAP7_75t_L g136 ( .A1(n_5), .A2(n_137), .B(n_144), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_6), .B(n_130), .Y(n_505) );
AND2x6_ASAP7_75t_L g142 ( .A(n_7), .B(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_8), .A2(n_236), .B(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_9), .B(n_39), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_9), .B(n_39), .Y(n_120) );
INVx1_ASAP7_75t_L g154 ( .A(n_10), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_11), .B(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g135 ( .A(n_12), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_13), .B(n_167), .Y(n_451) );
INVx1_ASAP7_75t_L g242 ( .A(n_14), .Y(n_242) );
INVx1_ASAP7_75t_L g509 ( .A(n_15), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_16), .B(n_131), .Y(n_490) );
AO32x2_ASAP7_75t_L g471 ( .A1(n_17), .A2(n_130), .A3(n_164), .B1(n_472), .B2(n_476), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_18), .B(n_157), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_19), .B(n_183), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_20), .B(n_131), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_21), .A2(n_50), .B1(n_157), .B2(n_456), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_22), .B(n_137), .Y(n_207) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_23), .A2(n_77), .B1(n_157), .B2(n_167), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_24), .B(n_157), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_25), .B(n_128), .Y(n_186) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_26), .A2(n_240), .B(n_241), .C(n_243), .Y(n_239) );
OAI22xp5_ASAP7_75t_SL g724 ( .A1(n_27), .A2(n_75), .B1(n_725), .B2(n_726), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_27), .Y(n_726) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_28), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_29), .B(n_160), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_30), .B(n_152), .Y(n_197) );
INVx1_ASAP7_75t_L g173 ( .A(n_31), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_32), .B(n_160), .Y(n_469) );
INVx2_ASAP7_75t_L g140 ( .A(n_33), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_34), .B(n_157), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_35), .B(n_160), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_36), .A2(n_63), .B1(n_745), .B2(n_746), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_36), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_37), .A2(n_142), .B(n_147), .C(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g171 ( .A(n_40), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_41), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_42), .B(n_152), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_43), .B(n_157), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_44), .A2(n_87), .B1(n_214), .B2(n_456), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_45), .B(n_157), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_46), .B(n_157), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g174 ( .A(n_47), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_48), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_49), .B(n_137), .Y(n_230) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_51), .A2(n_61), .B1(n_157), .B2(n_167), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_52), .A2(n_102), .B1(n_111), .B2(n_756), .Y(n_101) );
AOI22xp5_ASAP7_75t_L g166 ( .A1(n_53), .A2(n_147), .B1(n_167), .B2(n_169), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g217 ( .A(n_54), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_55), .B(n_157), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_56), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_57), .B(n_157), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g150 ( .A1(n_58), .A2(n_151), .B(n_153), .C(n_156), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_59), .Y(n_260) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
INVx1_ASAP7_75t_L g143 ( .A(n_62), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_63), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_64), .B(n_157), .Y(n_515) );
INVx1_ASAP7_75t_L g134 ( .A(n_65), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_66), .Y(n_739) );
AO32x2_ASAP7_75t_L g481 ( .A1(n_67), .A2(n_130), .A3(n_222), .B1(n_476), .B2(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g526 ( .A(n_68), .Y(n_526) );
INVx1_ASAP7_75t_L g464 ( .A(n_69), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_SL g182 ( .A1(n_70), .A2(n_156), .B(n_183), .C(n_184), .Y(n_182) );
INVxp67_ASAP7_75t_L g185 ( .A(n_71), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_72), .B(n_167), .Y(n_465) );
INVx1_ASAP7_75t_L g110 ( .A(n_73), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_74), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_75), .Y(n_725) );
INVx1_ASAP7_75t_L g253 ( .A(n_76), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_78), .A2(n_142), .B(n_147), .C(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_79), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_80), .B(n_167), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_81), .B(n_196), .Y(n_210) );
INVx2_ASAP7_75t_L g132 ( .A(n_82), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_83), .B(n_183), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_84), .B(n_167), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_85), .A2(n_142), .B(n_147), .C(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g107 ( .A(n_86), .Y(n_107) );
OR2x2_ASAP7_75t_L g117 ( .A(n_86), .B(n_118), .Y(n_117) );
OR2x2_ASAP7_75t_L g749 ( .A(n_86), .B(n_735), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_88), .A2(n_100), .B1(n_167), .B2(n_168), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_89), .B(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_90), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_91), .A2(n_142), .B(n_147), .C(n_225), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_92), .Y(n_232) );
INVx1_ASAP7_75t_L g181 ( .A(n_93), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g238 ( .A(n_94), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_95), .B(n_196), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_96), .B(n_167), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_97), .B(n_130), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_98), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_99), .A2(n_137), .B(n_180), .Y(n_179) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g756 ( .A(n_104), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g439 ( .A(n_107), .B(n_118), .Y(n_439) );
NOR2x2_ASAP7_75t_L g734 ( .A(n_107), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
AO221x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_737), .B1(n_740), .B2(n_750), .C(n_752), .Y(n_111) );
OAI222xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_723), .B1(n_724), .B2(n_727), .C1(n_731), .C2(n_736), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_121), .B1(n_438), .B2(n_440), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g728 ( .A(n_117), .Y(n_728) );
INVx2_ASAP7_75t_L g735 ( .A(n_118), .Y(n_735) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_121), .A2(n_729), .B1(n_743), .B2(n_744), .Y(n_742) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g729 ( .A(n_122), .Y(n_729) );
AND3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_360), .C(n_405), .Y(n_122) );
NOR4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_283), .C(n_324), .D(n_341), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_187), .B(n_203), .C(n_245), .Y(n_124) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_126), .B(n_188), .Y(n_187) );
NOR4xp25_ASAP7_75t_L g307 ( .A(n_126), .B(n_301), .C(n_308), .D(n_314), .Y(n_307) );
AND2x2_ASAP7_75t_L g380 ( .A(n_126), .B(n_269), .Y(n_380) );
AND2x2_ASAP7_75t_L g399 ( .A(n_126), .B(n_345), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_126), .B(n_394), .Y(n_408) );
AND2x2_ASAP7_75t_L g421 ( .A(n_126), .B(n_202), .Y(n_421) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_SL g266 ( .A(n_127), .Y(n_266) );
AND2x2_ASAP7_75t_L g273 ( .A(n_127), .B(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g323 ( .A(n_127), .B(n_162), .Y(n_323) );
AND2x2_ASAP7_75t_SL g334 ( .A(n_127), .B(n_269), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_127), .B(n_162), .Y(n_338) );
AND2x2_ASAP7_75t_L g347 ( .A(n_127), .B(n_272), .Y(n_347) );
BUFx2_ASAP7_75t_L g370 ( .A(n_127), .Y(n_370) );
AND2x2_ASAP7_75t_L g374 ( .A(n_127), .B(n_178), .Y(n_374) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_136), .B(n_159), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_129), .B(n_217), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g491 ( .A(n_129), .B(n_476), .C(n_492), .Y(n_491) );
AO21x1_ASAP7_75t_L g529 ( .A1(n_129), .A2(n_492), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_130), .A2(n_179), .B(n_186), .Y(n_178) );
OA21x2_ASAP7_75t_L g496 ( .A1(n_130), .A2(n_497), .B(n_505), .Y(n_496) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
AND2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_132), .B(n_133), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
BUFx2_ASAP7_75t_L g236 ( .A(n_137), .Y(n_236) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_142), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_138), .B(n_142), .Y(n_175) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_141), .Y(n_138) );
INVx1_ASAP7_75t_L g504 ( .A(n_139), .Y(n_504) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx1_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
INVx1_ASAP7_75t_L g149 ( .A(n_141), .Y(n_149) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_141), .Y(n_155) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_141), .Y(n_170) );
INVx1_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
INVx4_ASAP7_75t_SL g158 ( .A(n_142), .Y(n_158) );
OAI21xp5_ASAP7_75t_L g448 ( .A1(n_142), .A2(n_449), .B(n_453), .Y(n_448) );
OAI21xp5_ASAP7_75t_L g462 ( .A1(n_142), .A2(n_463), .B(n_466), .Y(n_462) );
BUFx3_ASAP7_75t_L g476 ( .A(n_142), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_142), .A2(n_498), .B(n_501), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_142), .A2(n_508), .B(n_512), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_150), .C(n_158), .Y(n_144) );
O2A1O1Ixp33_ASAP7_75t_L g180 ( .A1(n_146), .A2(n_158), .B(n_181), .C(n_182), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_146), .A2(n_158), .B(n_238), .C(n_239), .Y(n_237) );
INVx5_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_148), .Y(n_157) );
BUFx3_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
INVx1_ASAP7_75t_L g456 ( .A(n_148), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_151), .A2(n_454), .B(n_455), .Y(n_453) );
O2A1O1Ixp5_ASAP7_75t_L g525 ( .A1(n_151), .A2(n_513), .B(n_526), .C(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx4_ASAP7_75t_L g228 ( .A(n_152), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_152), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
OAI22xp5_ASAP7_75t_SL g482 ( .A1(n_152), .A2(n_155), .B1(n_483), .B2(n_484), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_152), .A2(n_474), .B1(n_493), .B2(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_155), .B(n_185), .Y(n_184) );
INVx5_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
O2A1O1Ixp5_ASAP7_75t_SL g463 ( .A1(n_156), .A2(n_196), .B(n_464), .C(n_465), .Y(n_463) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
HB1xp67_ASAP7_75t_L g229 ( .A(n_157), .Y(n_229) );
OAI22xp33_ASAP7_75t_L g165 ( .A1(n_158), .A2(n_166), .B1(n_174), .B2(n_175), .Y(n_165) );
INVx1_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
INVx2_ASAP7_75t_L g222 ( .A(n_160), .Y(n_222) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_160), .A2(n_235), .B(n_244), .Y(n_234) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_160), .A2(n_448), .B(n_457), .Y(n_447) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_160), .A2(n_462), .B(n_469), .Y(n_461) );
OR2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_178), .Y(n_161) );
AND2x2_ASAP7_75t_L g202 ( .A(n_162), .B(n_178), .Y(n_202) );
BUFx2_ASAP7_75t_L g276 ( .A(n_162), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_162), .A2(n_309), .B1(n_311), .B2(n_312), .Y(n_308) );
OR2x2_ASAP7_75t_L g330 ( .A(n_162), .B(n_190), .Y(n_330) );
AND2x2_ASAP7_75t_L g394 ( .A(n_162), .B(n_272), .Y(n_394) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g262 ( .A(n_163), .B(n_190), .Y(n_262) );
AND2x2_ASAP7_75t_L g269 ( .A(n_163), .B(n_178), .Y(n_269) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_163), .Y(n_311) );
OR2x2_ASAP7_75t_L g346 ( .A(n_163), .B(n_189), .Y(n_346) );
AO21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_176), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_164), .B(n_177), .Y(n_176) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_164), .A2(n_191), .B(n_199), .Y(n_190) );
INVx2_ASAP7_75t_L g215 ( .A(n_164), .Y(n_215) );
INVx2_ASAP7_75t_L g198 ( .A(n_167), .Y(n_198) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_170), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_169) );
INVx2_ASAP7_75t_L g172 ( .A(n_170), .Y(n_172) );
INVx4_ASAP7_75t_L g240 ( .A(n_170), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_175), .A2(n_192), .B(n_193), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_175), .A2(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g265 ( .A(n_178), .Y(n_265) );
INVx3_ASAP7_75t_L g274 ( .A(n_178), .Y(n_274) );
BUFx2_ASAP7_75t_L g298 ( .A(n_178), .Y(n_298) );
AND2x2_ASAP7_75t_L g331 ( .A(n_178), .B(n_266), .Y(n_331) );
INVx1_ASAP7_75t_L g452 ( .A(n_183), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_187), .A2(n_417), .B1(n_418), .B2(n_419), .Y(n_416) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_202), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_189), .B(n_274), .Y(n_278) );
INVx1_ASAP7_75t_L g306 ( .A(n_189), .Y(n_306) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g272 ( .A(n_190), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .C(n_198), .Y(n_194) );
INVx2_ASAP7_75t_L g474 ( .A(n_196), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_196), .A2(n_499), .B(n_500), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_196), .A2(n_523), .B(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_198), .A2(n_509), .B(n_510), .C(n_511), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_200), .B(n_201), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_201), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_201), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g284 ( .A(n_202), .Y(n_284) );
NAND2x1_ASAP7_75t_SL g203 ( .A(n_204), .B(n_218), .Y(n_203) );
AND2x2_ASAP7_75t_L g282 ( .A(n_204), .B(n_233), .Y(n_282) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_204), .Y(n_356) );
AND2x2_ASAP7_75t_L g383 ( .A(n_204), .B(n_303), .Y(n_383) );
AND2x2_ASAP7_75t_L g391 ( .A(n_204), .B(n_353), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_204), .B(n_248), .Y(n_418) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g249 ( .A(n_205), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g267 ( .A(n_205), .B(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g288 ( .A(n_205), .Y(n_288) );
INVx1_ASAP7_75t_L g294 ( .A(n_205), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_205), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_205), .B(n_251), .Y(n_327) );
OR2x2_ASAP7_75t_L g365 ( .A(n_205), .B(n_320), .Y(n_365) );
AOI32xp33_ASAP7_75t_L g377 ( .A1(n_205), .A2(n_378), .A3(n_381), .B1(n_382), .B2(n_383), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_205), .B(n_353), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_205), .B(n_313), .Y(n_428) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_216), .Y(n_205) );
AOI21xp5_ASAP7_75t_SL g206 ( .A1(n_207), .A2(n_208), .B(n_215), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_212), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_212), .A2(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g243 ( .A(n_214), .Y(n_243) );
INVx1_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
OA21x2_ASAP7_75t_L g506 ( .A1(n_215), .A2(n_507), .B(n_516), .Y(n_506) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_215), .A2(n_521), .B(n_528), .Y(n_520) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
OR2x2_ASAP7_75t_L g339 ( .A(n_219), .B(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_233), .Y(n_219) );
INVx1_ASAP7_75t_L g301 ( .A(n_220), .Y(n_301) );
AND2x2_ASAP7_75t_L g303 ( .A(n_220), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_220), .B(n_250), .Y(n_320) );
AND2x2_ASAP7_75t_L g353 ( .A(n_220), .B(n_329), .Y(n_353) );
AND2x2_ASAP7_75t_L g390 ( .A(n_220), .B(n_251), .Y(n_390) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g248 ( .A(n_221), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_221), .B(n_250), .Y(n_280) );
AND2x2_ASAP7_75t_L g287 ( .A(n_221), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g328 ( .A(n_221), .B(n_329), .Y(n_328) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_231), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_229), .Y(n_225) );
INVx2_ASAP7_75t_L g304 ( .A(n_233), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_233), .B(n_250), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_233), .B(n_295), .Y(n_376) );
INVx1_ASAP7_75t_L g398 ( .A(n_233), .Y(n_398) );
INVx1_ASAP7_75t_L g415 ( .A(n_233), .Y(n_415) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g268 ( .A(n_234), .B(n_250), .Y(n_268) );
AND2x2_ASAP7_75t_L g290 ( .A(n_234), .B(n_251), .Y(n_290) );
INVx1_ASAP7_75t_L g329 ( .A(n_234), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_240), .B(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_240), .A2(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g511 ( .A(n_240), .Y(n_511) );
AOI221x1_ASAP7_75t_SL g245 ( .A1(n_246), .A2(n_261), .B1(n_267), .B2(n_269), .C(n_270), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_246), .A2(n_334), .B1(n_401), .B2(n_402), .Y(n_400) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
AND2x2_ASAP7_75t_L g292 ( .A(n_247), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g387 ( .A(n_247), .B(n_267), .Y(n_387) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g343 ( .A(n_248), .B(n_268), .Y(n_343) );
INVx1_ASAP7_75t_L g355 ( .A(n_249), .Y(n_355) );
AND2x2_ASAP7_75t_L g366 ( .A(n_249), .B(n_353), .Y(n_366) );
AND2x2_ASAP7_75t_L g433 ( .A(n_249), .B(n_328), .Y(n_433) );
INVx2_ASAP7_75t_L g295 ( .A(n_250), .Y(n_295) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_258), .B(n_259), .Y(n_251) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_262), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g385 ( .A(n_262), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_263), .B(n_346), .Y(n_349) );
INVx3_ASAP7_75t_SL g263 ( .A(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_264), .A2(n_385), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_SL g407 ( .A(n_267), .B(n_293), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_268), .B(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g359 ( .A(n_268), .B(n_287), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_268), .B(n_294), .Y(n_436) );
AND2x2_ASAP7_75t_L g305 ( .A(n_269), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g372 ( .A(n_269), .Y(n_372) );
AOI21xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_275), .B(n_279), .Y(n_270) );
NAND2x1_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_272), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g321 ( .A(n_272), .B(n_322), .Y(n_321) );
INVx1_ASAP7_75t_SL g333 ( .A(n_272), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_272), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g357 ( .A(n_273), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_273), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_273), .B(n_276), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AOI211xp5_ASAP7_75t_L g344 ( .A1(n_276), .A2(n_315), .B(n_345), .C(n_347), .Y(n_344) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_276), .A2(n_363), .B1(n_366), .B2(n_367), .C(n_371), .Y(n_362) );
AND2x2_ASAP7_75t_L g358 ( .A(n_277), .B(n_311), .Y(n_358) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g318 ( .A(n_282), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g389 ( .A(n_282), .B(n_390), .Y(n_389) );
OAI211xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B(n_291), .C(n_316), .Y(n_283) );
NAND3xp33_ASAP7_75t_SL g402 ( .A(n_284), .B(n_403), .C(n_404), .Y(n_402) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
OR2x2_ASAP7_75t_L g375 ( .A(n_286), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_296), .B1(n_299), .B2(n_305), .C(n_307), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_293), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_293), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_298), .A2(n_355), .B1(n_356), .B2(n_357), .Y(n_354) );
OR2x2_ASAP7_75t_L g435 ( .A(n_298), .B(n_346), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVxp67_ASAP7_75t_L g409 ( .A(n_301), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_303), .B(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g310 ( .A(n_304), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_306), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_306), .B(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_306), .B(n_373), .Y(n_412) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_310), .Y(n_336) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g426 ( .A(n_315), .B(n_346), .Y(n_426) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_321), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g404 ( .A(n_321), .Y(n_404) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI322xp33_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_330), .A3(n_331), .B1(n_332), .B2(n_335), .C1(n_337), .C2(n_339), .Y(n_324) );
OAI322xp33_ASAP7_75t_L g406 ( .A1(n_325), .A2(n_407), .A3(n_408), .B1(n_409), .B2(n_410), .C1(n_411), .C2(n_413), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx4_ASAP7_75t_L g340 ( .A(n_327), .Y(n_340) );
AND2x2_ASAP7_75t_L g401 ( .A(n_327), .B(n_353), .Y(n_401) );
AND2x2_ASAP7_75t_L g414 ( .A(n_327), .B(n_415), .Y(n_414) );
CKINVDCx16_ASAP7_75t_R g425 ( .A(n_330), .Y(n_425) );
INVx1_ASAP7_75t_L g403 ( .A(n_331), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OR2x2_ASAP7_75t_L g337 ( .A(n_333), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g420 ( .A(n_333), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_333), .B(n_374), .Y(n_431) );
OR2x2_ASAP7_75t_L g364 ( .A(n_336), .B(n_365), .Y(n_364) );
INVxp33_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
OAI221xp5_ASAP7_75t_SL g341 ( .A1(n_340), .A2(n_342), .B1(n_344), .B2(n_348), .C(n_350), .Y(n_341) );
NOR2xp67_ASAP7_75t_L g397 ( .A(n_340), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g424 ( .A(n_340), .Y(n_424) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AOI322xp5_ASAP7_75t_L g388 ( .A1(n_347), .A2(n_372), .A3(n_389), .B1(n_391), .B2(n_392), .C1(n_395), .C2(n_399), .Y(n_388) );
INVxp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_354), .B1(n_358), .B2(n_359), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_384), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_377), .Y(n_361) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_365), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp33_ASAP7_75t_SL g382 ( .A(n_368), .B(n_379), .Y(n_382) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
OAI322xp33_ASAP7_75t_L g422 ( .A1(n_370), .A2(n_423), .A3(n_425), .B1(n_426), .B2(n_427), .C1(n_429), .C2(n_432), .Y(n_422) );
AOI21xp33_ASAP7_75t_SL g371 ( .A1(n_372), .A2(n_373), .B(n_375), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_380), .B(n_428), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g384 ( .A1(n_385), .A2(n_386), .B(n_388), .C(n_400), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR4xp25_ASAP7_75t_L g405 ( .A(n_406), .B(n_416), .C(n_422), .D(n_434), .Y(n_405) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
CKINVDCx14_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_436), .B(n_437), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx6_ASAP7_75t_L g730 ( .A(n_439), .Y(n_730) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_441), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_645), .Y(n_441) );
NAND5xp2_ASAP7_75t_L g442 ( .A(n_443), .B(n_564), .C(n_579), .D(n_605), .E(n_627), .Y(n_442) );
NOR2xp33_ASAP7_75t_SL g443 ( .A(n_444), .B(n_544), .Y(n_443) );
OAI221xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_485), .B1(n_517), .B2(n_533), .C(n_534), .Y(n_444) );
NOR2xp33_ASAP7_75t_SL g445 ( .A(n_446), .B(n_477), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_446), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g721 ( .A(n_446), .Y(n_721) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_458), .Y(n_446) );
INVx1_ASAP7_75t_L g561 ( .A(n_447), .Y(n_561) );
AND2x2_ASAP7_75t_L g563 ( .A(n_447), .B(n_471), .Y(n_563) );
AND2x2_ASAP7_75t_L g573 ( .A(n_447), .B(n_470), .Y(n_573) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_447), .Y(n_591) );
INVx1_ASAP7_75t_L g601 ( .A(n_447), .Y(n_601) );
OR2x2_ASAP7_75t_L g639 ( .A(n_447), .B(n_538), .Y(n_639) );
INVx2_ASAP7_75t_L g689 ( .A(n_447), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_447), .B(n_537), .Y(n_706) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B(n_452), .Y(n_449) );
NOR2xp67_ASAP7_75t_L g458 ( .A(n_459), .B(n_470), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_460), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_460), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_460), .B(n_561), .Y(n_621) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_461), .Y(n_479) );
INVx2_ASAP7_75t_L g538 ( .A(n_461), .Y(n_538) );
OR2x2_ASAP7_75t_L g600 ( .A(n_461), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g539 ( .A(n_470), .B(n_481), .Y(n_539) );
AND2x2_ASAP7_75t_L g556 ( .A(n_470), .B(n_536), .Y(n_556) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g480 ( .A(n_471), .B(n_481), .Y(n_480) );
BUFx2_ASAP7_75t_L g559 ( .A(n_471), .Y(n_559) );
AND2x2_ASAP7_75t_L g688 ( .A(n_471), .B(n_689), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_474), .A2(n_502), .B(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_474), .A2(n_513), .B(n_514), .C(n_515), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_476), .A2(n_522), .B(n_525), .Y(n_521) );
INVx1_ASAP7_75t_L g533 ( .A(n_477), .Y(n_533) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
AND2x2_ASAP7_75t_L g651 ( .A(n_478), .B(n_539), .Y(n_651) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g652 ( .A(n_479), .B(n_563), .Y(n_652) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_480), .A2(n_620), .B(n_622), .C(n_624), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_480), .B(n_620), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_480), .A2(n_550), .B1(n_693), .B2(n_694), .C(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g536 ( .A(n_481), .Y(n_536) );
INVx1_ASAP7_75t_L g572 ( .A(n_481), .Y(n_572) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_481), .Y(n_581) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_495), .Y(n_486) );
AND2x2_ASAP7_75t_L g598 ( .A(n_487), .B(n_543), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_487), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_488), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g690 ( .A(n_488), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g722 ( .A(n_488), .Y(n_722) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g552 ( .A(n_489), .Y(n_552) );
AND2x2_ASAP7_75t_L g578 ( .A(n_489), .B(n_532), .Y(n_578) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_489), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g594 ( .A(n_489), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx1_ASAP7_75t_L g530 ( .A(n_490), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_495), .B(n_634), .Y(n_669) );
INVx1_ASAP7_75t_SL g673 ( .A(n_495), .Y(n_673) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_506), .Y(n_495) );
INVx3_ASAP7_75t_L g532 ( .A(n_496), .Y(n_532) );
AND2x2_ASAP7_75t_L g543 ( .A(n_496), .B(n_520), .Y(n_543) );
AND2x2_ASAP7_75t_L g565 ( .A(n_496), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g610 ( .A(n_496), .B(n_604), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_496), .B(n_542), .Y(n_691) );
INVx2_ASAP7_75t_L g513 ( .A(n_504), .Y(n_513) );
AND2x2_ASAP7_75t_L g531 ( .A(n_506), .B(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g542 ( .A(n_506), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g603 ( .A(n_506), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_531), .Y(n_518) );
INVx1_ASAP7_75t_L g583 ( .A(n_519), .Y(n_583) );
AND2x2_ASAP7_75t_L g625 ( .A(n_519), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_519), .B(n_546), .Y(n_631) );
AOI21xp5_ASAP7_75t_SL g705 ( .A1(n_519), .A2(n_537), .B(n_560), .Y(n_705) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
OR2x2_ASAP7_75t_L g548 ( .A(n_520), .B(n_529), .Y(n_548) );
AND2x2_ASAP7_75t_L g595 ( .A(n_520), .B(n_532), .Y(n_595) );
INVx2_ASAP7_75t_L g604 ( .A(n_520), .Y(n_604) );
INVx1_ASAP7_75t_L g710 ( .A(n_520), .Y(n_710) );
AND2x2_ASAP7_75t_L g634 ( .A(n_529), .B(n_604), .Y(n_634) );
INVx1_ASAP7_75t_L g659 ( .A(n_529), .Y(n_659) );
AND2x2_ASAP7_75t_L g568 ( .A(n_531), .B(n_552), .Y(n_568) );
AND2x2_ASAP7_75t_L g580 ( .A(n_531), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g698 ( .A(n_531), .Y(n_698) );
INVx2_ASAP7_75t_L g588 ( .A(n_532), .Y(n_588) );
AND2x2_ASAP7_75t_L g626 ( .A(n_532), .B(n_542), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_532), .B(n_710), .Y(n_709) );
OAI21xp33_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_539), .B(n_540), .Y(n_534) );
AND2x2_ASAP7_75t_L g641 ( .A(n_535), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g695 ( .A(n_535), .Y(n_695) );
AND2x2_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g615 ( .A(n_536), .Y(n_615) );
BUFx2_ASAP7_75t_L g714 ( .A(n_536), .Y(n_714) );
BUFx2_ASAP7_75t_L g585 ( .A(n_537), .Y(n_585) );
AND2x2_ASAP7_75t_L g687 ( .A(n_537), .B(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g670 ( .A(n_538), .Y(n_670) );
AND2x4_ASAP7_75t_L g597 ( .A(n_539), .B(n_560), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_539), .B(n_621), .Y(n_633) );
AOI32xp33_ASAP7_75t_L g557 ( .A1(n_540), .A2(n_558), .A3(n_560), .B1(n_562), .B2(n_563), .Y(n_557) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx3_ASAP7_75t_L g546 ( .A(n_541), .Y(n_546) );
OR2x2_ASAP7_75t_L g682 ( .A(n_541), .B(n_638), .Y(n_682) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g551 ( .A(n_542), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g658 ( .A(n_542), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g550 ( .A(n_543), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g562 ( .A(n_543), .B(n_552), .Y(n_562) );
INVx1_ASAP7_75t_L g683 ( .A(n_543), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_543), .B(n_658), .Y(n_716) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_549), .B(n_553), .C(n_557), .Y(n_544) );
OAI322xp33_ASAP7_75t_L g653 ( .A1(n_545), .A2(n_590), .A3(n_654), .B1(n_656), .B2(n_660), .C1(n_661), .C2(n_665), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVxp67_ASAP7_75t_L g618 ( .A(n_546), .Y(n_618) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g672 ( .A(n_548), .B(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_548), .B(n_588), .Y(n_719) );
INVxp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g611 ( .A(n_551), .Y(n_611) );
OR2x2_ASAP7_75t_L g697 ( .A(n_552), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_555), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g606 ( .A(n_556), .B(n_585), .Y(n_606) );
AND2x2_ASAP7_75t_L g677 ( .A(n_556), .B(n_590), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_556), .B(n_664), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g564 ( .A1(n_558), .A2(n_565), .B1(n_568), .B2(n_569), .C(n_574), .Y(n_564) );
OR2x2_ASAP7_75t_L g575 ( .A(n_558), .B(n_571), .Y(n_575) );
AND2x2_ASAP7_75t_L g663 ( .A(n_558), .B(n_664), .Y(n_663) );
AOI32xp33_ASAP7_75t_L g702 ( .A1(n_558), .A2(n_588), .A3(n_703), .B1(n_704), .B2(n_707), .Y(n_702) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g636 ( .A(n_559), .B(n_595), .C(n_618), .Y(n_636) );
AND2x2_ASAP7_75t_L g662 ( .A(n_559), .B(n_655), .Y(n_662) );
INVxp67_ASAP7_75t_L g642 ( .A(n_560), .Y(n_642) );
BUFx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_563), .B(n_615), .Y(n_671) );
INVx2_ASAP7_75t_L g681 ( .A(n_563), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_563), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g650 ( .A(n_566), .Y(n_650) );
OR2x2_ASAP7_75t_L g576 ( .A(n_567), .B(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_569), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_572), .Y(n_655) );
AND2x2_ASAP7_75t_L g614 ( .A(n_573), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g660 ( .A(n_573), .Y(n_660) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_573), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
AOI21xp33_ASAP7_75t_SL g599 ( .A1(n_575), .A2(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g693 ( .A(n_578), .B(n_603), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B(n_592), .C(n_599), .Y(n_579) );
AND2x2_ASAP7_75t_L g623 ( .A(n_581), .B(n_591), .Y(n_623) );
INVx2_ASAP7_75t_L g638 ( .A(n_581), .Y(n_638) );
OR2x2_ASAP7_75t_L g676 ( .A(n_581), .B(n_639), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_581), .B(n_719), .Y(n_718) );
AOI211xp5_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_584), .B(n_586), .C(n_589), .Y(n_582) );
INVxp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_585), .B(n_623), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g704 ( .A1(n_586), .A2(n_681), .B(n_705), .C(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_587), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g644 ( .A(n_588), .B(n_634), .Y(n_644) );
INVx1_ASAP7_75t_L g649 ( .A(n_588), .Y(n_649) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_593), .B(n_596), .Y(n_592) );
INVxp33_ASAP7_75t_L g700 ( .A(n_594), .Y(n_700) );
AND2x2_ASAP7_75t_L g679 ( .A(n_595), .B(n_658), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_600), .A2(n_662), .B(n_663), .Y(n_661) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_602), .A2(n_681), .A3(n_682), .B1(n_683), .B2(n_684), .C1(n_686), .C2(n_690), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_612), .B2(n_616), .C(n_619), .Y(n_605) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g657 ( .A(n_610), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g701 ( .A(n_614), .Y(n_701) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_617), .B(n_637), .Y(n_703) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g666 ( .A(n_626), .B(n_634), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_630), .B1(n_632), .B2(n_634), .C(n_635), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_630), .A2(n_647), .B1(n_651), .B2(n_652), .C(n_653), .Y(n_646) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_634), .B(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_640), .B2(n_643), .Y(n_635) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx2_ASAP7_75t_SL g664 ( .A(n_639), .Y(n_664) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND5xp2_ASAP7_75t_L g645 ( .A(n_646), .B(n_667), .C(n_692), .D(n_702), .E(n_712), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_648), .B(n_650), .Y(n_647) );
NOR4xp25_ASAP7_75t_L g720 ( .A(n_649), .B(n_655), .C(n_721), .D(n_722), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_652), .A2(n_713), .B1(n_715), .B2(n_717), .C(n_720), .Y(n_712) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g711 ( .A(n_658), .Y(n_711) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_662), .A2(n_669), .A3(n_670), .B1(n_671), .B2(n_672), .C1(n_674), .C2(n_678), .Y(n_668) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_668), .B(n_680), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g713 ( .A(n_688), .B(n_714), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_696) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_SL g751 ( .A(n_738), .Y(n_751) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_SL g741 ( .A(n_742), .B(n_747), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g755 ( .A(n_749), .Y(n_755) );
BUFx3_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
endmodule