module real_jpeg_32359_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_0),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_44),
.B1(n_186),
.B2(n_189),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_2),
.A2(n_17),
.B1(n_21),
.B2(n_23),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_3),
.B(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_3),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_3),
.A2(n_294),
.B(n_302),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_3),
.B(n_144),
.Y(n_439)
);

OAI22xp33_ASAP7_75t_SL g466 ( 
.A1(n_3),
.A2(n_31),
.B1(n_450),
.B2(n_467),
.Y(n_466)
);

OAI32xp33_ASAP7_75t_L g487 ( 
.A1(n_3),
.A2(n_175),
.A3(n_383),
.B1(n_488),
.B2(n_489),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g492 ( 
.A1(n_3),
.A2(n_169),
.B1(n_316),
.B2(n_335),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_4),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_6),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_6),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_6),
.A2(n_76),
.B1(n_155),
.B2(n_160),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_6),
.A2(n_76),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_7),
.A2(n_105),
.B1(n_108),
.B2(n_112),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_7),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_7),
.A2(n_112),
.B1(n_165),
.B2(n_230),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_7),
.A2(n_112),
.B1(n_357),
.B2(n_359),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_7),
.A2(n_112),
.B1(n_376),
.B2(n_378),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_8),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_8),
.A2(n_168),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_8),
.A2(n_168),
.B1(n_224),
.B2(n_260),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_8),
.A2(n_168),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_9),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_9),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_10),
.Y(n_149)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_11),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_12),
.A2(n_221),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_12),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_12),
.A2(n_225),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_12),
.A2(n_225),
.B1(n_243),
.B2(n_443),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g459 ( 
.A1(n_12),
.A2(n_50),
.B1(n_225),
.B2(n_460),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_13),
.A2(n_291),
.B1(n_320),
.B2(n_324),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_13),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_13),
.A2(n_324),
.B1(n_340),
.B2(n_343),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_13),
.A2(n_324),
.B1(n_408),
.B2(n_412),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_13),
.A2(n_324),
.B1(n_451),
.B2(n_456),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_14),
.A2(n_91),
.B1(n_92),
.B2(n_97),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_14),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_14),
.A2(n_91),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_14),
.A2(n_91),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_15),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_50),
.B1(n_53),
.B2(n_57),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_16),
.A2(n_57),
.B1(n_205),
.B2(n_242),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_18),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_19),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_19),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_19),
.A2(n_128),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_19),
.A2(n_128),
.B1(n_357),
.B2(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_19),
.A2(n_128),
.B1(n_430),
.B2(n_433),
.Y(n_429)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_267),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_265),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_233),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_26),
.B(n_233),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_182),
.C(n_197),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_28),
.B(n_183),
.Y(n_550)
);

XNOR2x1_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_101),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_29),
.B(n_235),
.C(n_236),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_58),
.Y(n_29)
);

XOR2x2_ASAP7_75t_L g530 ( 
.A(n_30),
.B(n_58),
.Y(n_530)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_37),
.B1(n_45),
.B2(n_49),
.Y(n_30)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_31),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_31),
.A2(n_37),
.B1(n_209),
.B2(n_215),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_31),
.A2(n_429),
.B1(n_435),
.B2(n_437),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_31),
.A2(n_450),
.B1(n_459),
.B2(n_463),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_34),
.Y(n_379)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_36),
.Y(n_332)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_36),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_36),
.Y(n_434)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_36),
.Y(n_458)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_41),
.Y(n_283)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_47),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_47),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_48),
.Y(n_478)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_49),
.Y(n_196)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_51),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_53),
.Y(n_470)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_62),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_56),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_75),
.B1(n_87),
.B2(n_90),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_59),
.A2(n_87),
.B1(n_90),
.B2(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_59),
.A2(n_75),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_59),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_59),
.A2(n_201),
.B1(n_202),
.B2(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_59),
.A2(n_201),
.B1(n_356),
.B2(n_366),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_59),
.A2(n_201),
.B1(n_441),
.B2(n_442),
.Y(n_440)
);

AO21x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_68),
.B(n_72),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_66),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_68),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B(n_81),
.Y(n_75)
);

BUFx2_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_79),
.Y(n_406)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_82),
.Y(n_359)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_86),
.Y(n_370)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_86),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_88),
.A2(n_240),
.B1(n_245),
.B2(n_246),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_88),
.A2(n_245),
.B1(n_367),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_89),
.Y(n_201)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_99),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_100),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_143),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_102),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_113),
.B1(n_124),
.B2(n_133),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_104),
.A2(n_134),
.B1(n_259),
.B2(n_264),
.Y(n_258)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_107),
.Y(n_223)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_107),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_110),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_111),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_113),
.A2(n_124),
.B1(n_133),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_113),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_113),
.B(n_335),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_113),
.A2(n_133),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g533 ( 
.A1(n_113),
.A2(n_124),
.B1(n_133),
.B2(n_220),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_135),
.Y(n_134)
);

AOI22x1_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_117),
.Y(n_290)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_119),
.Y(n_293)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_119),
.Y(n_353)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_119),
.Y(n_390)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_120),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_133),
.Y(n_523)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

AO22x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_154),
.B1(n_162),
.B2(n_173),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_144),
.A2(n_154),
.B1(n_248),
.B2(n_253),
.Y(n_247)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_144),
.Y(n_318)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AO21x2_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_175),
.B(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_152),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_159),
.Y(n_250)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_163),
.A2(n_174),
.B1(n_229),
.B2(n_232),
.Y(n_228)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_164),
.Y(n_307)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_170),
.Y(n_231)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_171),
.Y(n_252)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_171),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_172),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g253 ( 
.A(n_174),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_174),
.A2(n_311),
.B1(n_318),
.B2(n_319),
.Y(n_310)
);

OA22x2_ASAP7_75t_L g347 ( 
.A1(n_174),
.A2(n_311),
.B1(n_318),
.B2(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_174),
.A2(n_232),
.B1(n_319),
.B2(n_492),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_174),
.A2(n_229),
.B1(n_232),
.B2(n_348),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_L g382 ( 
.A1(n_175),
.A2(n_383),
.B(n_389),
.Y(n_382)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_192),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_184),
.B(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_190),
.Y(n_412)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_192),
.A2(n_193),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B(n_196),
.Y(n_193)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_194),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_195),
.A2(n_277),
.B1(n_278),
.B2(n_281),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_195),
.A2(n_281),
.B1(n_327),
.B2(n_333),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_195),
.A2(n_327),
.B1(n_375),
.B2(n_380),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_195),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_197),
.B(n_550),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_218),
.C(n_226),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_199),
.B(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_200),
.B(n_208),
.Y(n_510)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_201),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_201),
.B(n_335),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_210),
.Y(n_417)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_211),
.Y(n_284)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_211),
.Y(n_455)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_216),
.Y(n_333)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_SL g381 ( 
.A(n_217),
.Y(n_381)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_217),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_218),
.A2(n_227),
.B1(n_228),
.B2(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_220),
.Y(n_524)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_254),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_247),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_245),
.A2(n_401),
.B1(n_407),
.B2(n_413),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

AOI22x1_ASAP7_75t_L g521 ( 
.A1(n_264),
.A2(n_522),
.B1(n_523),
.B2(n_524),
.Y(n_521)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_544),
.B(n_551),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_505),
.B(n_541),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_394),
.B(n_504),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_360),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_272),
.B(n_360),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_336),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_309),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_274),
.B(n_309),
.C(n_336),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_285),
.B2(n_308),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_275),
.B(n_285),
.Y(n_526)
);

INVxp67_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_279),
.B(n_335),
.Y(n_469)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_285),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_294),
.B(n_299),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_288),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_300),
.C(n_307),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_325),
.C(n_334),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_310),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_325),
.A2(n_326),
.B1(n_334),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_334),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_384),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_390),
.C(n_391),
.Y(n_389)
);

OAI21xp33_ASAP7_75t_SL g401 ( 
.A1(n_335),
.A2(n_402),
.B(n_404),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_335),
.B(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_337),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_339),
.Y(n_522)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_354),
.B2(n_355),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g512 ( 
.A(n_347),
.B(n_354),
.C(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_365),
.C(n_371),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_361),
.A2(n_362),
.B1(n_498),
.B2(n_499),
.Y(n_497)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_365),
.A2(n_371),
.B1(n_372),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_365),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_370),
.Y(n_443)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_382),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_373),
.A2(n_374),
.B1(n_382),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_391),
.Y(n_489)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_496),
.B(n_503),
.Y(n_394)
);

AOI21x1_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_482),
.B(n_495),
.Y(n_395)
);

OAI21x1_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_446),
.B(n_481),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_427),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_427),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_414),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_399),
.A2(n_400),
.B1(n_414),
.B2(n_415),
.Y(n_479)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_407),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_422),
.B1(n_423),
.B2(n_426),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_438),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_428),
.B(n_440),
.C(n_444),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_440),
.B1(n_444),
.B2(n_445),
.Y(n_438)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_439),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_440),
.Y(n_445)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_472),
.B(n_480),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_465),
.B(n_471),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_464),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_449),
.B(n_464),
.Y(n_471)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx4_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_459),
.Y(n_474)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_468),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_479),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_479),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_484),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_490),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_493),
.C(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_491),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_501),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_501),
.Y(n_503)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_506),
.B(n_536),
.Y(n_505)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_527),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_508),
.B(n_527),
.C(n_543),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_511),
.C(n_514),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_510),
.Y(n_509)
);

XNOR2x1_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_512),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

XNOR2x1_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_539),
.Y(n_538)
);

XNOR2x1_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_526),
.Y(n_514)
);

OAI21x1_ASAP7_75t_L g515 ( 
.A1(n_516),
.A2(n_519),
.B(n_525),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_526),
.C(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_518),
.B(n_521),
.Y(n_525)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_521),
.Y(n_535)
);

XNOR2x1_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_534),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_534),
.C(n_548),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_537),
.Y(n_536)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_540),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_540),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_549),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_547),
.B(n_549),
.Y(n_553)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);


endmodule