module fake_aes_12205_n_658 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_658);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_658;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g77 ( .A(n_74), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_30), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_18), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_16), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_54), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_75), .Y(n_84) );
INVxp33_ASAP7_75t_SL g85 ( .A(n_60), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_31), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_19), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_0), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_21), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_0), .Y(n_91) );
BUFx2_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
CKINVDCx20_ASAP7_75t_R g93 ( .A(n_7), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_7), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_4), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_52), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_62), .Y(n_98) );
INVxp33_ASAP7_75t_SL g99 ( .A(n_33), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_15), .Y(n_100) );
INVxp33_ASAP7_75t_L g101 ( .A(n_8), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_2), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_10), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_26), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_57), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_3), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_51), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_59), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_68), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_50), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_49), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_23), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_56), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_67), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_11), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_48), .Y(n_118) );
BUFx5_ASAP7_75t_L g119 ( .A(n_6), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_119), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_92), .B(n_1), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_119), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_119), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_92), .B(n_1), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_119), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_108), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_119), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_119), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_101), .B(n_2), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_118), .B(n_3), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_91), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_119), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_114), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_114), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_82), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_93), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
BUFx12f_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_95), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_112), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_112), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_82), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_95), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_116), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_88), .B(n_5), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
OAI22xp5_ASAP7_75t_SL g152 ( .A1(n_116), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_95), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_95), .Y(n_154) );
NAND2x1_ASAP7_75t_L g155 ( .A(n_88), .B(n_12), .Y(n_155) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_124), .B(n_87), .Y(n_156) );
INVx1_ASAP7_75t_SL g157 ( .A(n_141), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_149), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_141), .B(n_104), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_133), .B(n_111), .Y(n_161) );
BUFx3_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_149), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_120), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_139), .B(n_105), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_124), .B(n_102), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_135), .B(n_111), .Y(n_171) );
BUFx10_ASAP7_75t_L g172 ( .A(n_124), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_132), .A2(n_85), .B1(n_99), .B2(n_79), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_139), .B(n_98), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_142), .B(n_99), .Y(n_177) );
OR2x2_ASAP7_75t_SL g178 ( .A(n_121), .B(n_102), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_146), .B(n_86), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_146), .B(n_110), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_150), .B(n_110), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_132), .Y(n_184) );
OR2x2_ASAP7_75t_L g185 ( .A(n_130), .B(n_106), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_131), .Y(n_188) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_151), .A2(n_98), .B(n_90), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_130), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_151), .B(n_85), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_122), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_137), .B(n_106), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_122), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_123), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_123), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_131), .Y(n_197) );
NAND3xp33_ASAP7_75t_L g198 ( .A(n_155), .B(n_117), .C(n_100), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_137), .B(n_94), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_155), .B(n_81), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_175), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_172), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_157), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_175), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
NOR2xp33_ASAP7_75t_R g206 ( .A(n_182), .B(n_127), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_156), .B(n_148), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_164), .A2(n_125), .B(n_126), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_176), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_186), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_191), .B(n_125), .Y(n_212) );
AND2x6_ASAP7_75t_SL g213 ( .A(n_200), .B(n_140), .Y(n_213) );
INVx4_ASAP7_75t_L g214 ( .A(n_172), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_189), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_193), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g217 ( .A(n_173), .B(n_136), .C(n_126), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_169), .B(n_136), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_193), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_156), .A2(n_152), .B1(n_115), .B2(n_80), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_182), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_179), .B(n_129), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_163), .A2(n_129), .B(n_138), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_180), .B(n_138), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_193), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_181), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_183), .B(n_77), .Y(n_228) );
NOR2xp67_ASAP7_75t_L g229 ( .A(n_198), .B(n_12), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_184), .B(n_113), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_163), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_190), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_184), .B(n_103), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_170), .B(n_96), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_163), .A2(n_177), .B1(n_170), .B2(n_160), .Y(n_235) );
NOR3xp33_ASAP7_75t_SL g236 ( .A(n_161), .B(n_90), .C(n_78), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_181), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g238 ( .A1(n_200), .A2(n_95), .B1(n_97), .B2(n_109), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_171), .B(n_107), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_199), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_197), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_170), .B(n_145), .Y(n_242) );
BUFx3_ASAP7_75t_L g243 ( .A(n_172), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_199), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_200), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_185), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_189), .Y(n_247) );
BUFx4f_ASAP7_75t_L g248 ( .A(n_200), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_185), .B(n_145), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_199), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_162), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_174), .B(n_134), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_165), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_211), .A2(n_167), .B(n_196), .C(n_168), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_251), .Y(n_257) );
BUFx4f_ASAP7_75t_L g258 ( .A(n_208), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_218), .A2(n_167), .B(n_196), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_222), .A2(n_168), .B(n_195), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_250), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_248), .A2(n_178), .B1(n_194), .B2(n_192), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_243), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_209), .A2(n_166), .B(n_197), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_203), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_211), .Y(n_266) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_215), .B(n_166), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
CKINVDCx8_ASAP7_75t_R g269 ( .A(n_213), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_219), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_215), .A2(n_153), .B(n_143), .Y(n_271) );
INVxp33_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_235), .B(n_178), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_246), .A2(n_143), .B(n_153), .C(n_162), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_251), .Y(n_276) );
INVx2_ASAP7_75t_SL g277 ( .A(n_221), .Y(n_277) );
BUFx6f_ASAP7_75t_L g278 ( .A(n_243), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_234), .B(n_187), .Y(n_279) );
BUFx2_ASAP7_75t_L g280 ( .A(n_248), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_240), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_248), .A2(n_187), .B1(n_134), .B2(n_144), .Y(n_282) );
O2A1O1Ixp5_ASAP7_75t_SL g283 ( .A1(n_249), .A2(n_153), .B(n_143), .C(n_154), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_224), .A2(n_153), .B(n_188), .C(n_145), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_232), .B(n_13), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_245), .A2(n_187), .B1(n_145), .B2(n_144), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_212), .A2(n_188), .B(n_145), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_245), .A2(n_145), .B1(n_144), .B2(n_134), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_223), .A2(n_144), .B(n_134), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_233), .B(n_13), .Y(n_291) );
NOR2xp67_ASAP7_75t_SL g292 ( .A(n_214), .B(n_144), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_220), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_254), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_234), .B(n_144), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_214), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_254), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_214), .B(n_14), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_201), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_234), .A2(n_134), .B1(n_154), .B2(n_147), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_205), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_201), .Y(n_302) );
INVx1_ASAP7_75t_SL g303 ( .A(n_233), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_208), .A2(n_134), .B1(n_154), .B2(n_147), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_252), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_257), .Y(n_306) );
AO31x2_ASAP7_75t_L g307 ( .A1(n_284), .A2(n_247), .A3(n_224), .B(n_207), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_257), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_298), .B(n_202), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_298), .B(n_202), .Y(n_310) );
BUFx12f_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_298), .B(n_231), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_266), .B(n_205), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_276), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_276), .A2(n_207), .B1(n_210), .B2(n_247), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_299), .Y(n_316) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_284), .A2(n_236), .B(n_242), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_256), .A2(n_225), .B(n_228), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_299), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_278), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_301), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_294), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_273), .A2(n_217), .B1(n_210), .B2(n_230), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_273), .A2(n_255), .B1(n_238), .B2(n_229), .Y(n_327) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_239), .B1(n_255), .B2(n_231), .C(n_241), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_278), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_265), .B(n_231), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_268), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_256), .A2(n_253), .B1(n_147), .B2(n_154), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_271), .A2(n_241), .B(n_237), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_262), .B(n_253), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_278), .Y(n_336) );
OAI21x1_ASAP7_75t_L g337 ( .A1(n_283), .A2(n_237), .B(n_227), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_259), .A2(n_253), .B(n_227), .C(n_204), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_316), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_321), .B(n_265), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_335), .A2(n_258), .B1(n_293), .B2(n_291), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_311), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_335), .A2(n_304), .B1(n_258), .B2(n_293), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_314), .B(n_280), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_317), .A2(n_274), .B(n_286), .Y(n_346) );
AO21x2_ASAP7_75t_L g347 ( .A1(n_332), .A2(n_267), .B(n_287), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_321), .B(n_325), .Y(n_348) );
BUFx12f_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_325), .A2(n_272), .B1(n_261), .B2(n_285), .C(n_281), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_323), .B(n_275), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_309), .Y(n_353) );
BUFx12f_ASAP7_75t_L g354 ( .A(n_311), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_331), .A2(n_272), .B1(n_290), .B2(n_279), .C(n_295), .Y(n_355) );
OAI211xp5_ASAP7_75t_L g356 ( .A1(n_327), .A2(n_269), .B(n_289), .C(n_300), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_328), .A2(n_263), .B1(n_296), .B2(n_260), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_315), .A2(n_263), .B1(n_267), .B2(n_296), .Y(n_358) );
OR3x1_ASAP7_75t_L g359 ( .A(n_323), .B(n_15), .C(n_16), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_316), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_331), .A2(n_288), .B1(n_282), .B2(n_264), .C(n_292), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_319), .Y(n_363) );
OAI22xp33_ASAP7_75t_L g364 ( .A1(n_328), .A2(n_302), .B1(n_305), .B2(n_252), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_312), .A2(n_305), .B1(n_252), .B2(n_204), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_351), .B(n_306), .Y(n_366) );
BUFx2_ASAP7_75t_L g367 ( .A(n_339), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_342), .B(n_330), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_351), .B(n_306), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_344), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_348), .B(n_306), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_344), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_360), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_360), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_360), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_352), .B(n_326), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_362), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_341), .A2(n_317), .B1(n_326), .B2(n_318), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g382 ( .A(n_356), .B(n_332), .C(n_318), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_362), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_362), .B(n_308), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_340), .B(n_308), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_363), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_363), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
INVx4_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_353), .B(n_308), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_345), .B(n_319), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_345), .B(n_307), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_343), .B(n_324), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_343), .B(n_307), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_369), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_367), .B(n_307), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_389), .B(n_334), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_367), .B(n_307), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_385), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_389), .B(n_342), .Y(n_403) );
OAI21xp33_ASAP7_75t_L g404 ( .A1(n_381), .A2(n_350), .B(n_327), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_377), .B(n_307), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_381), .A2(n_359), .B1(n_355), .B2(n_334), .C(n_330), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_373), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_368), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_396), .A2(n_317), .B1(n_312), .B2(n_310), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_377), .B(n_307), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_392), .B(n_307), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_372), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_373), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_385), .A2(n_359), .B1(n_310), .B2(n_309), .Y(n_416) );
OAI22xp5_ASAP7_75t_SL g417 ( .A1(n_379), .A2(n_349), .B1(n_354), .B2(n_317), .Y(n_417) );
AOI33xp33_ASAP7_75t_L g418 ( .A1(n_395), .A2(n_330), .A3(n_357), .B1(n_312), .B2(n_365), .B3(n_364), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_392), .B(n_317), .Y(n_420) );
OAI33xp33_ASAP7_75t_L g421 ( .A1(n_396), .A2(n_358), .A3(n_315), .B1(n_313), .B2(n_18), .B3(n_17), .Y(n_421) );
OR2x6_ASAP7_75t_L g422 ( .A(n_390), .B(n_358), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_378), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_379), .B(n_354), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_394), .B(n_324), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_376), .B(n_347), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_376), .B(n_347), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_309), .B1(n_310), .B2(n_349), .Y(n_428) );
INVx4_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx4_ASAP7_75t_L g430 ( .A(n_391), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_395), .A2(n_312), .B1(n_310), .B2(n_309), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_371), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_394), .B(n_324), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_376), .B(n_310), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_378), .B(n_347), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_383), .B(n_336), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_370), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_383), .B(n_336), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_366), .Y(n_439) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_370), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_413), .B(n_393), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_402), .B(n_393), .Y(n_443) );
AND2x4_ASAP7_75t_L g444 ( .A(n_426), .B(n_393), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_432), .B(n_366), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_409), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_426), .B(n_388), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_425), .B(n_388), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_413), .B(n_370), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_405), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_425), .B(n_386), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_398), .B(n_370), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_375), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_404), .A2(n_382), .B1(n_391), .B2(n_309), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_401), .B(n_375), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_439), .B(n_386), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_401), .B(n_375), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_415), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_433), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_426), .B(n_372), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_424), .B(n_382), .C(n_147), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_423), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_399), .B(n_384), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_406), .B(n_387), .Y(n_470) );
AND2x4_ASAP7_75t_SL g471 ( .A(n_419), .B(n_391), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_421), .A2(n_346), .B1(n_391), .B2(n_312), .C(n_147), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_416), .A2(n_384), .B(n_346), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_408), .Y(n_474) );
AND2x4_ASAP7_75t_SL g475 ( .A(n_429), .B(n_387), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_403), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_400), .B(n_380), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_433), .B(n_380), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_427), .B(n_380), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_407), .A2(n_147), .B1(n_154), .B2(n_361), .C(n_374), .Y(n_480) );
NOR2xp67_ASAP7_75t_L g481 ( .A(n_429), .B(n_354), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_397), .B(n_372), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_406), .B(n_387), .Y(n_483) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_397), .B(n_374), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_412), .B(n_420), .Y(n_487) );
NOR2x1p5_ASAP7_75t_L g488 ( .A(n_430), .B(n_349), .Y(n_488) );
NAND4xp25_ASAP7_75t_L g489 ( .A(n_411), .B(n_313), .C(n_338), .D(n_329), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_410), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_412), .B(n_154), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_435), .B(n_17), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_435), .B(n_322), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_430), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_431), .B(n_336), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_410), .B(n_336), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_486), .B(n_428), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_487), .B(n_437), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_461), .B(n_414), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_482), .B(n_417), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_492), .B(n_430), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_446), .B(n_414), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_485), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_487), .B(n_427), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_464), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_441), .B(n_427), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_441), .B(n_422), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_450), .B(n_422), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_459), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_491), .B(n_418), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_450), .B(n_422), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_491), .B(n_436), .Y(n_512) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_464), .B(n_436), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_484), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_443), .B(n_422), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_445), .B(n_436), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_459), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_447), .B(n_438), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_460), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_468), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_454), .B(n_440), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_481), .B(n_434), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_463), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_454), .B(n_438), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_457), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_442), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_456), .B(n_434), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_456), .B(n_434), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_458), .B(n_322), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_449), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_449), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_452), .Y(n_534) );
NAND2xp33_ASAP7_75t_SL g535 ( .A(n_488), .B(n_322), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_458), .B(n_470), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_475), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_462), .B(n_20), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_452), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_469), .B(n_470), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_483), .B(n_336), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_483), .B(n_320), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_442), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_475), .Y(n_544) );
NOR2x1_ASAP7_75t_L g545 ( .A(n_466), .B(n_320), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_476), .B(n_320), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_443), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_477), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_478), .B(n_320), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_453), .B(n_320), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_453), .B(n_322), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_448), .B(n_322), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_527), .B(n_485), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_497), .A2(n_462), .B1(n_485), .B2(n_471), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_505), .Y(n_555) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_537), .A2(n_513), .B1(n_505), .B2(n_544), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_500), .A2(n_494), .B1(n_455), .B2(n_471), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_498), .Y(n_558) );
OAI211xp5_ASAP7_75t_SL g559 ( .A1(n_510), .A2(n_472), .B(n_480), .C(n_495), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_498), .Y(n_560) );
AO22x2_ASAP7_75t_L g561 ( .A1(n_503), .A2(n_494), .B1(n_448), .B2(n_465), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_537), .A2(n_448), .B(n_473), .C(n_465), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_503), .B(n_489), .Y(n_563) );
OAI321xp33_ASAP7_75t_L g564 ( .A1(n_513), .A2(n_493), .A3(n_496), .B1(n_490), .B2(n_474), .C(n_467), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_536), .B(n_493), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_513), .A2(n_479), .B1(n_465), .B2(n_444), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_548), .B(n_479), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_525), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_525), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_547), .B(n_479), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_522), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_501), .A2(n_444), .B(n_474), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_509), .Y(n_573) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_546), .A2(n_444), .B(n_467), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_507), .A2(n_490), .B1(n_451), .B2(n_329), .Y(n_575) );
INVxp67_ASAP7_75t_L g576 ( .A(n_514), .Y(n_576) );
AO22x1_ASAP7_75t_L g577 ( .A1(n_503), .A2(n_451), .B1(n_329), .B2(n_322), .Y(n_577) );
OAI21xp33_ASAP7_75t_L g578 ( .A1(n_507), .A2(n_322), .B(n_337), .Y(n_578) );
INVx4_ASAP7_75t_L g579 ( .A(n_552), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_508), .A2(n_337), .B1(n_333), .B2(n_252), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_532), .B(n_337), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_536), .B(n_22), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_529), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_517), .Y(n_584) );
NAND2xp33_ASAP7_75t_SL g585 ( .A(n_529), .B(n_24), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_519), .Y(n_586) );
OAI21xp33_ASAP7_75t_SL g587 ( .A1(n_524), .A2(n_333), .B(n_27), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_508), .B(n_25), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_506), .B(n_28), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_538), .B(n_333), .C(n_32), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_520), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_535), .A2(n_252), .B1(n_34), .B2(n_35), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_521), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_556), .B(n_535), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_561), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_568), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_569), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_573), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_584), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_586), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_591), .Y(n_601) );
AOI222xp33_ASAP7_75t_L g602 ( .A1(n_587), .A2(n_533), .B1(n_534), .B2(n_539), .C1(n_518), .C2(n_523), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_593), .B(n_540), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_567), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_587), .A2(n_516), .B(n_515), .C(n_499), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_557), .A2(n_511), .B1(n_530), .B2(n_512), .Y(n_606) );
NAND2x1_ASAP7_75t_L g607 ( .A(n_561), .B(n_545), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_565), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_558), .B(n_526), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_583), .B(n_506), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_579), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_553), .Y(n_612) );
XOR2x2_ASAP7_75t_L g613 ( .A(n_554), .B(n_530), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_560), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_554), .A2(n_511), .B1(n_526), .B2(n_504), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_563), .A2(n_504), .B1(n_522), .B2(n_515), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_571), .Y(n_617) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_585), .A2(n_502), .B(n_542), .C(n_541), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_596), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_602), .A2(n_579), .B1(n_559), .B2(n_576), .Y(n_620) );
OAI321xp33_ASAP7_75t_L g621 ( .A1(n_594), .A2(n_562), .A3(n_566), .B1(n_575), .B2(n_582), .C(n_570), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_611), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_598), .Y(n_623) );
AOI21xp33_ASAP7_75t_L g624 ( .A1(n_602), .A2(n_588), .B(n_564), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_595), .A2(n_572), .B(n_592), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g626 ( .A(n_613), .B(n_588), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_605), .A2(n_574), .B1(n_555), .B2(n_578), .C(n_581), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_597), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_616), .A2(n_589), .B1(n_590), .B2(n_592), .Y(n_629) );
OAI211xp5_ASAP7_75t_SL g630 ( .A1(n_606), .A2(n_580), .B(n_549), .C(n_550), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_615), .A2(n_550), .B1(n_549), .B2(n_528), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_612), .A2(n_551), .B1(n_552), .B2(n_531), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_604), .B(n_543), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_624), .A2(n_607), .B1(n_608), .B2(n_603), .Y(n_634) );
AOI221x1_ASAP7_75t_L g635 ( .A1(n_619), .A2(n_600), .B1(n_601), .B2(n_599), .C(n_603), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_625), .A2(n_614), .B1(n_617), .B2(n_618), .C1(n_609), .C2(n_610), .Y(n_636) );
OAI211xp5_ASAP7_75t_SL g637 ( .A1(n_620), .A2(n_618), .B(n_609), .C(n_543), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_630), .A2(n_551), .B1(n_531), .B2(n_528), .Y(n_638) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_621), .A2(n_577), .B(n_36), .C(n_37), .Y(n_639) );
AO221x1_ASAP7_75t_L g640 ( .A1(n_622), .A2(n_76), .B1(n_38), .B2(n_39), .C(n_40), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_626), .B(n_29), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g642 ( .A1(n_627), .A2(n_41), .B(n_42), .C(n_43), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_634), .B(n_623), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_635), .B(n_628), .Y(n_644) );
XNOR2xp5_ASAP7_75t_L g645 ( .A(n_642), .B(n_629), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_638), .B(n_632), .Y(n_646) );
NAND4xp75_ASAP7_75t_L g647 ( .A(n_641), .B(n_633), .C(n_631), .D(n_47), .Y(n_647) );
OA22x2_ASAP7_75t_L g648 ( .A1(n_645), .A2(n_640), .B1(n_636), .B2(n_637), .Y(n_648) );
OR4x2_ASAP7_75t_L g649 ( .A(n_643), .B(n_639), .C(n_46), .D(n_53), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_646), .B(n_643), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_650), .Y(n_651) );
INVx3_ASAP7_75t_L g652 ( .A(n_648), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_651), .Y(n_653) );
AO22x2_ASAP7_75t_L g654 ( .A1(n_652), .A2(n_644), .B1(n_648), .B2(n_647), .Y(n_654) );
AOI22x1_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_652), .B1(n_644), .B2(n_649), .Y(n_655) );
AOI222xp33_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_653), .B1(n_644), .B2(n_58), .C1(n_63), .C2(n_64), .Y(n_656) );
OA22x2_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_45), .B1(n_55), .B2(n_65), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_69), .B1(n_70), .B2(n_72), .C(n_73), .Y(n_658) );
endmodule