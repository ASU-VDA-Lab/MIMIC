module fake_jpeg_31033_n_316 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_316);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_53),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_56),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_18),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_62),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_29),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_45),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_73),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_0),
.C(n_1),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_43),
.C(n_46),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_34),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_76),
.Y(n_113)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_1),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_2),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_34),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_75),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_52),
.A2(n_39),
.B1(n_26),
.B2(n_30),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_24),
.B1(n_28),
.B2(n_32),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_92),
.A2(n_95),
.B1(n_44),
.B2(n_50),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_30),
.B1(n_26),
.B2(n_24),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_30),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_57),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_62),
.A2(n_28),
.B1(n_44),
.B2(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_35),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_35),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_43),
.B1(n_38),
.B2(n_37),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_47),
.A2(n_27),
.B1(n_23),
.B2(n_37),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_114),
.A2(n_117),
.B1(n_142),
.B2(n_112),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_85),
.B(n_81),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_118),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_112),
.A2(n_48),
.B1(n_61),
.B2(n_60),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_38),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_128),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_120),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_130),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_27),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_125),
.B(n_127),
.Y(n_149)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_23),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_87),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_64),
.B1(n_51),
.B2(n_34),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_14),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_134),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_35),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_138),
.C(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_144),
.Y(n_161)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_141),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_17),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_98),
.B(n_35),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_66),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_105),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_57),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_116),
.A2(n_84),
.B1(n_94),
.B2(n_97),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_121),
.B1(n_138),
.B2(n_130),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_127),
.Y(n_168)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_143),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_172),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_150),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_125),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_135),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_177),
.B1(n_160),
.B2(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_138),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_144),
.B1(n_116),
.B2(n_110),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_179),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_139),
.C(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_175),
.C(n_173),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_145),
.B(n_134),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_181),
.A2(n_148),
.B(n_158),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_153),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_182),
.B1(n_168),
.B2(n_160),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_151),
.B1(n_149),
.B2(n_146),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_198),
.C(n_180),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_190),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_192),
.A2(n_181),
.B(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_110),
.B1(n_63),
.B2(n_55),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_164),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_211),
.B(n_214),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_197),
.B(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_155),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_181),
.B(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_199),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_179),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_189),
.C(n_194),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_183),
.B(n_184),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_214),
.B(n_200),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_174),
.B1(n_198),
.B2(n_196),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_229),
.B1(n_202),
.B2(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_230),
.C(n_227),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_206),
.A2(n_169),
.B1(n_178),
.B2(n_194),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_208),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_185),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_208),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_162),
.B1(n_157),
.B2(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_185),
.C(n_154),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_247),
.C(n_166),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_242),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_152),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_225),
.Y(n_251)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_221),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_238),
.B(n_240),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_244),
.B1(n_216),
.B2(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_228),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_207),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_245),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_219),
.A2(n_205),
.B1(n_204),
.B2(n_200),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_153),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_212),
.C(n_154),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_256),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_222),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_254),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_247),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_255),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_239),
.A2(n_220),
.B1(n_216),
.B2(n_157),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_152),
.C(n_148),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_233),
.B1(n_245),
.B2(n_164),
.Y(n_258)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_163),
.C(n_123),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_107),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_264),
.B(n_2),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_166),
.C(n_158),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_267),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_165),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_266),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_165),
.B(n_129),
.Y(n_267)
);

NOR2x1_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_249),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_R g287 ( 
.A(n_268),
.B(n_4),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_272),
.C(n_250),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_163),
.C(n_162),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_163),
.C(n_132),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_162),
.C(n_86),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_134),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_283),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_271),
.A2(n_250),
.B1(n_262),
.B2(n_133),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_286),
.B1(n_111),
.B2(n_83),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_86),
.B1(n_111),
.B2(n_105),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_269),
.A2(n_122),
.B1(n_101),
.B2(n_83),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_285),
.B(n_287),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_2),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_272),
.B(n_270),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_291),
.B(n_294),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_281),
.A2(n_263),
.B(n_268),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_279),
.B(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_295),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_101),
.C(n_124),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_5),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_6),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_5),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_299),
.B(n_301),
.Y(n_305)
);

NOR4xp25_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_8),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_7),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_293),
.B1(n_10),
.B2(n_11),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

AOI321xp33_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_305),
.A3(n_307),
.B1(n_11),
.B2(n_8),
.C(n_10),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_300),
.B(n_109),
.Y(n_309)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_91),
.B(n_109),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_11),
.B1(n_74),
.B2(n_82),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_312),
.A2(n_313),
.B(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_91),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_91),
.Y(n_316)
);


endmodule