module real_jpeg_25773_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_228;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_244;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_31),
.B1(n_41),
.B2(n_42),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_31),
.B1(n_57),
.B2(n_61),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_31),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_9),
.B1(n_55),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_6),
.A2(n_57),
.B1(n_61),
.B2(n_64),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_64),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_44),
.B1(n_57),
.B2(n_61),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_8),
.Y(n_74)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_11),
.A2(n_28),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_11),
.A2(n_28),
.B1(n_57),
.B2(n_61),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_28),
.B1(n_41),
.B2(n_42),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_11),
.A2(n_60),
.B(n_107),
.C(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_11),
.B(n_56),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_11),
.A2(n_61),
.B(n_74),
.C(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_11),
.B(n_26),
.C(n_38),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_11),
.B(n_127),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_11),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_11),
.B(n_36),
.Y(n_232)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_273),
.B1(n_286),
.B2(n_287),
.Y(n_13)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_14),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_131),
.B(n_272),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_108),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_16),
.B(n_108),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.C(n_90),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_17),
.B(n_82),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_49),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_18),
.B(n_50),
.C(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_19),
.B(n_34),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_20),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_24),
.A2(n_32),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_24),
.B(n_32),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_26),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_28),
.A2(n_59),
.B(n_61),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_41),
.B(n_75),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_29),
.A2(n_94),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_29),
.B(n_219),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_84),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_32),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_32),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B(n_45),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_35),
.B(n_123),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_35),
.A2(n_87),
.B(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_36),
.B(n_48),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_36),
.B(n_189),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_47)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_40),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_42),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_42),
.B(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_45),
.B(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_46),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_46),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_69),
.B2(n_70),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_62),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_53),
.B(n_65),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_59),
.B1(n_60),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_63),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_56),
.B(n_105),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_61),
.B1(n_74),
.B2(n_75),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_71),
.B(n_153),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_71),
.A2(n_78),
.B(n_126),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_72),
.B(n_79),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_73),
.A2(n_79),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_73),
.B(n_101),
.Y(n_155)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_77),
.B(n_146),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_79),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_89),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_86),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_83),
.A2(n_89),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_83),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_83),
.A2(n_89),
.B1(n_184),
.B2(n_244),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g283 ( 
.A1(n_83),
.A2(n_112),
.B(n_114),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_88),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_88),
.B(n_188),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_90),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.C(n_102),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_91),
.A2(n_92),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_97),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_96),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_96),
.B(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_98),
.B(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_100),
.A2(n_102),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_100),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_102),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_130),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_119),
.B2(n_120),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_110),
.B(n_120),
.C(n_130),
.Y(n_284)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_125),
.B(n_129),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_125),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_128),
.B(n_145),
.Y(n_144)
);

FAx1_ASAP7_75t_L g275 ( 
.A(n_129),
.B(n_276),
.CI(n_283),
.CON(n_275),
.SN(n_275)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_267),
.B(n_271),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_178),
.B(n_253),
.C(n_266),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_166),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_134),
.B(n_166),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_150),
.B2(n_165),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_148),
.B2(n_149),
.Y(n_136)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_137),
.B(n_149),
.C(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_144),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_140),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_141),
.B(n_157),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_142),
.A2(n_143),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g154 ( 
.A(n_147),
.Y(n_154)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_160),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_152),
.B(n_159),
.C(n_160),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.C(n_173),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_168),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_173),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

FAx1_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.CI(n_177),
.CON(n_173),
.SN(n_173)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_252),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_193),
.B(n_251),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_190),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_181),
.B(n_190),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.C(n_186),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_182),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_186),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_246),
.B(n_250),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_237),
.B(n_245),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_216),
.B(n_236),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_197),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_210),
.B2(n_215),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_209),
.C(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_224),
.B(n_235),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_222),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_221),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_231),
.B(n_234),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_232),
.B(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_255),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_263),
.B2(n_264),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_264),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_285),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_284),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_275),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_282),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_277),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_278),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);


endmodule