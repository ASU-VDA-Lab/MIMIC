module real_jpeg_9127_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_24),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_1),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_1),
.A2(n_3),
.B(n_25),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_1),
.A2(n_78),
.B1(n_80),
.B2(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_1),
.A2(n_28),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_1),
.B(n_28),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_1),
.A2(n_69),
.B1(n_71),
.B2(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_1),
.A2(n_24),
.B(n_65),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_32),
.B1(n_80),
.B2(n_105),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_2),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_24),
.B(n_26),
.C(n_27),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_7),
.B(n_24),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_9),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_60),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_47),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_11),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_14),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_58),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_58),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_109),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_107),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_73),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_19),
.B(n_73),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_51),
.C(n_61),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_20),
.A2(n_21),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_35),
.B1(n_36),
.B2(n_50),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_23),
.A2(n_27),
.B1(n_33),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_155),
.Y(n_154)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_27),
.B(n_78),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_53),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_28),
.B(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_29),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_41),
.C(n_50),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_38),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_39),
.A2(n_40),
.B(n_80),
.C(n_103),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_80),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_42),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_42),
.A2(n_43),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_45),
.B1(n_53),
.B2(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_44),
.B(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_44),
.B(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_45),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_51),
.A2(n_61),
.B1(n_62),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_51),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_51)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_52),
.A2(n_55),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_52),
.A2(n_55),
.B1(n_124),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_52),
.A2(n_55),
.B1(n_57),
.B2(n_147),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_54),
.Y(n_128)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_55),
.B(n_78),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_68),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_63),
.B(n_68),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_69),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_69),
.A2(n_71),
.B1(n_116),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_78),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_89),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_98),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_158),
.B(n_164),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_150),
.B(n_157),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_141),
.B(n_149),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_130),
.B(n_140),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_125),
.B2(n_129),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_129),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_125),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_135),
.B(n_139),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_134),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_143),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_146),
.C(n_148),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_152),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_152),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.CI(n_156),
.CON(n_152),
.SN(n_152)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_160),
.Y(n_164)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);


endmodule