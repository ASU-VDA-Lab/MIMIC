module real_jpeg_6817_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_323;
wire n_166;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_1),
.A2(n_26),
.B1(n_140),
.B2(n_143),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_1),
.B(n_31),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_26),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_1),
.A2(n_26),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g311 ( 
.A1(n_1),
.A2(n_34),
.B(n_312),
.C(n_314),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_1),
.B(n_126),
.C(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_1),
.B(n_114),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_1),
.B(n_179),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_1),
.B(n_128),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_2),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_2),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_15),
.B1(n_18),
.B2(n_20),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_4),
.A2(n_73),
.B1(n_110),
.B2(n_113),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_4),
.A2(n_73),
.B1(n_324),
.B2(n_326),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_4),
.A2(n_73),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_5),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_6),
.Y(n_185)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_6),
.Y(n_204)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_7),
.Y(n_155)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g429 ( 
.A(n_10),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_11),
.A2(n_169),
.B1(n_170),
.B2(n_174),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_11),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_11),
.A2(n_143),
.B1(n_169),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_11),
.A2(n_169),
.B1(n_287),
.B2(n_291),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_11),
.A2(n_169),
.B1(n_428),
.B2(n_430),
.Y(n_427)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_12),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_13),
.A2(n_35),
.B1(n_46),
.B2(n_107),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_13),
.A2(n_46),
.B1(n_134),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_46),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_454),
.Y(n_20)
);

OAI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_57),
.B1(n_61),
.B2(n_449),
.C(n_452),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_22),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_22),
.B(n_57),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_23),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_24),
.B(n_224),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_48),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_29),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g314 ( 
.A1(n_26),
.A2(n_315),
.B(n_317),
.Y(n_314)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_28),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_29),
.Y(n_158)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_30),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_31),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_31),
.B(n_44),
.Y(n_223)
);

AO22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_38),
.B2(n_41),
.Y(n_31)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_32),
.Y(n_166)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_36),
.Y(n_152)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_37),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_37),
.Y(n_290)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_43),
.B(n_70),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_43),
.A2(n_58),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_48),
.B(n_71),
.Y(n_224)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_51),
.Y(n_53)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_57),
.A2(n_268),
.B1(n_272),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_57),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_57),
.A2(n_272),
.B(n_278),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_59),
.B(n_60),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_59),
.A2(n_223),
.B(n_427),
.Y(n_445)
);

A2O1A1O1Ixp25_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_405),
.B(n_438),
.C(n_441),
.D(n_448),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_397),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_256),
.C(n_301),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_232),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_205),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_66),
.B(n_205),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_146),
.C(n_189),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_67),
.B(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_77),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_68),
.B(n_78),
.C(n_116),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_69),
.B(n_223),
.Y(n_412)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_115),
.B1(n_116),
.B2(n_145),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_108),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_80),
.A2(n_114),
.B(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_80),
.B(n_227),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_105),
.Y(n_80)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_94),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_88),
.B1(n_90),
.B2(n_93),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_87),
.Y(n_316)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_94),
.B(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_97),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_99),
.Y(n_218)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_99),
.Y(n_325)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g336 ( 
.A(n_101),
.Y(n_336)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_102),
.Y(n_216)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_102),
.Y(n_328)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_106),
.B(n_114),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_108),
.B(n_266),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_109),
.B(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_112),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_114),
.A2(n_193),
.B(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_115),
.A2(n_116),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_115),
.A2(n_116),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_115),
.B(n_412),
.C(n_416),
.Y(n_436)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_116),
.B(n_434),
.C(n_435),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_137),
.B(n_138),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_117),
.A2(n_213),
.B(n_243),
.Y(n_271)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_118),
.B(n_214),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_118),
.B(n_323),
.Y(n_322)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_128),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_128),
.B(n_323),
.Y(n_341)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_134),
.B2(n_136),
.Y(n_128)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_133),
.Y(n_183)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_133),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_137),
.A2(n_243),
.B(n_247),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_137),
.B(n_138),
.Y(n_294)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_142),
.Y(n_318)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_146),
.A2(n_147),
.B1(n_189),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_167),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_148),
.B(n_167),
.Y(n_220)
);

AOI32xp33_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_153),
.A3(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_177),
.B(n_180),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_201),
.B(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_173),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_174),
.Y(n_349)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_177),
.Y(n_269)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_186),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_181),
.A2(n_198),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_181),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_185),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_188),
.Y(n_371)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_189),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.C(n_196),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_190),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_191),
.B(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_191),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_193),
.B(n_229),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_193),
.A2(n_286),
.B(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_196),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_197),
.B(n_361),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_201),
.B(n_345),
.Y(n_375)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_204),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_219),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_208),
.C(n_219),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_211),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_212),
.B(n_341),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_213),
.B(n_322),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.C(n_225),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_229),
.Y(n_228)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_230),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_232),
.A2(n_400),
.B(n_401),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_255),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_233),
.B(n_255),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_236),
.C(n_248),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_248),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_238),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_241),
.B(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_247),
.B(n_341),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.C(n_253),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_251),
.A2(n_253),
.B1(n_444),
.B2(n_445),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_251),
.B(n_445),
.C(n_446),
.Y(n_451)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_298),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_257),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_274),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_258),
.B(n_274),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_267),
.C(n_273),
.Y(n_258)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_259),
.B(n_267),
.CI(n_273),
.CON(n_299),
.SN(n_299)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_264),
.C(n_265),
.Y(n_297)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_267)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_271),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_268),
.A2(n_272),
.B1(n_311),
.B2(n_388),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_297),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_283),
.B2(n_284),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_277),
.B(n_283),
.C(n_297),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_293),
.B(n_296),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_293),
.Y(n_296)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_296),
.A2(n_409),
.B1(n_410),
.B2(n_418),
.Y(n_408)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_296),
.Y(n_418)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_299),
.B(n_300),
.Y(n_402)
);

BUFx24_ASAP7_75t_SL g456 ( 
.A(n_299),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_329),
.B(n_396),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_306),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_303),
.B(n_306),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.C(n_319),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_307),
.B(n_392),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_310),
.A2(n_319),
.B1(n_320),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_390),
.B(n_395),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_380),
.B(n_389),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_355),
.B(n_379),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_342),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_342),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_340),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_334),
.A2(n_335),
.B1(n_340),
.B2(n_358),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_350),
.Y(n_342)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_351),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_352),
.B(n_353),
.C(n_382),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_364),
.B(n_378),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_357),
.B(n_359),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_359),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_374),
.B(n_377),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_373),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_372),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_375),
.B(n_376),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_383),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_383),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_385),
.B(n_386),
.C(n_387),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_394),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_394),
.Y(n_395)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_399),
.B(n_402),
.C(n_403),
.D(n_404),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_421),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_407),
.B(n_420),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_420),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_419),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_418),
.C(n_419),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_411),
.A2(n_412),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_424),
.C(n_436),
.Y(n_447)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_421),
.A2(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_437),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_437),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_436),
.Y(n_422)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_431),
.B1(n_432),
.B2(n_435),
.Y(n_425)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_426),
.Y(n_435)
);

INVx8_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_447),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_442),
.B(n_447),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g453 ( 
.A(n_451),
.Y(n_453)
);


endmodule