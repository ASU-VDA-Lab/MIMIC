module fake_ibex_1487_n_1749 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_340, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_323, n_143, n_106, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_331, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_335, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_329, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_320, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_324, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_319, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1749);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_323;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_335;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_320;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1749;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_550;
wire n_641;
wire n_557;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_1704;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_650;
wire n_409;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1694;
wire n_1458;
wire n_1460;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_348;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_648;
wire n_571;
wire n_1169;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1740;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1734;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_1744;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

OR2x2_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_33),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_150),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_248),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_253),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_221),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_61),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_236),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_64),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_15),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_302),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_216),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_17),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_70),
.B(n_90),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_39),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_34),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_187),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_20),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_196),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_257),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_214),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_291),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_83),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_311),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_103),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_16),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_107),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_118),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_227),
.Y(n_373)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_270),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_91),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_141),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_237),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_194),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_205),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_288),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_321),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_13),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_259),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_229),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_312),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g386 ( 
.A(n_314),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_91),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_107),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_325),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_322),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_232),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_166),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_271),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_297),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_211),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_207),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_68),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_180),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_319),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_180),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_21),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_316),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_113),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_186),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_71),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_162),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_33),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_25),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_122),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_332),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_228),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_245),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_294),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_63),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_260),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_304),
.B(n_277),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_22),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_284),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_301),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_231),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_39),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_111),
.Y(n_424)
);

BUFx8_ASAP7_75t_SL g425 ( 
.A(n_339),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_268),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_269),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_296),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_252),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_58),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_172),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_100),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_4),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_142),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_110),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_266),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_273),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_144),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_244),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_16),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_36),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_8),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_310),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_73),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_299),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_309),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_330),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_164),
.Y(n_448)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_8),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_49),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_97),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_278),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_142),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g454 ( 
.A(n_233),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_74),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_110),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_84),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_210),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_21),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_109),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_97),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_298),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_307),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_331),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_98),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_335),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_102),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_106),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_52),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_220),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_306),
.B(n_165),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_159),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_275),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_163),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_287),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_184),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_47),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_146),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_206),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_112),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_182),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_106),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_76),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_251),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_315),
.Y(n_485)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_163),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_209),
.Y(n_487)
);

BUFx10_ASAP7_75t_L g488 ( 
.A(n_267),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_274),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_151),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_65),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_81),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_117),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_176),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_3),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_38),
.Y(n_496)
);

BUFx5_ASAP7_75t_L g497 ( 
.A(n_280),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_66),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_255),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_114),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_272),
.Y(n_501)
);

BUFx5_ASAP7_75t_L g502 ( 
.A(n_153),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_254),
.B(n_276),
.Y(n_503)
);

BUFx8_ASAP7_75t_SL g504 ( 
.A(n_204),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_181),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_25),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_139),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_55),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_45),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_324),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_218),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_329),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_0),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_265),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_41),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_203),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_200),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_103),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_308),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_72),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_326),
.Y(n_521)
);

INVxp67_ASAP7_75t_SL g522 ( 
.A(n_202),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_4),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_43),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_1),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_286),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_215),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_305),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_95),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_246),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_264),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_109),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_320),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_121),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_56),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_53),
.Y(n_536)
);

BUFx10_ASAP7_75t_L g537 ( 
.A(n_226),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_80),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_77),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_69),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_80),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_197),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_176),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_38),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_285),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_258),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_141),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_150),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_240),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_105),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_247),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_290),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_303),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_256),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_23),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_43),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_166),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_281),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_10),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_242),
.Y(n_560)
);

CKINVDCx14_ASAP7_75t_R g561 ( 
.A(n_222),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_92),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_313),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_190),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_35),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_292),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_48),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_328),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_116),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_293),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_125),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_50),
.Y(n_572)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_44),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_137),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_113),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_238),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_23),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_94),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_289),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_28),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_27),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_279),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_282),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_6),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_72),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_88),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_384),
.A2(n_188),
.B(n_185),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_368),
.A2(n_191),
.B(n_189),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_425),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_396),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_382),
.B(n_0),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_486),
.B(n_1),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_502),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_520),
.B(n_2),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_375),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_351),
.B(n_2),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_377),
.Y(n_597)
);

AOI22x1_ASAP7_75t_SL g598 ( 
.A1(n_460),
.A2(n_6),
.B1(n_3),
.B2(n_5),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_377),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_375),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_502),
.Y(n_601)
);

AND2x6_ASAP7_75t_L g602 ( 
.A(n_397),
.B(n_192),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_502),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_348),
.B(n_7),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_377),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_425),
.Y(n_606)
);

NOR2x1_ASAP7_75t_L g607 ( 
.A(n_347),
.B(n_9),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_386),
.B(n_9),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_397),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_347),
.B(n_10),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_487),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_487),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_583),
.B(n_193),
.Y(n_616)
);

INVx6_ASAP7_75t_L g617 ( 
.A(n_396),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_359),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_359),
.Y(n_620)
);

OA21x2_ASAP7_75t_L g621 ( 
.A1(n_368),
.A2(n_445),
.B(n_383),
.Y(n_621)
);

AND2x2_ASAP7_75t_SL g622 ( 
.A(n_418),
.B(n_503),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_359),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_359),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_583),
.Y(n_625)
);

BUFx8_ASAP7_75t_SL g626 ( 
.A(n_460),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_441),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_627)
);

OA21x2_ASAP7_75t_L g628 ( 
.A1(n_383),
.A2(n_198),
.B(n_195),
.Y(n_628)
);

AOI22x1_ASAP7_75t_SL g629 ( 
.A1(n_524),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_359),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_396),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_357),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_445),
.Y(n_633)
);

BUFx12f_ASAP7_75t_L g634 ( 
.A(n_488),
.Y(n_634)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_488),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

BUFx3_ASAP7_75t_L g637 ( 
.A(n_458),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_458),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_541),
.B(n_14),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_409),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_470),
.A2(n_579),
.B(n_519),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_443),
.B(n_15),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_357),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_537),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_573),
.B(n_17),
.Y(n_646)
);

OA21x2_ASAP7_75t_L g647 ( 
.A1(n_470),
.A2(n_201),
.B(n_199),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_519),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_374),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_374),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_485),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_474),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_360),
.Y(n_654)
);

BUFx12f_ASAP7_75t_L g655 ( 
.A(n_361),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_409),
.B(n_18),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_374),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_435),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_374),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_374),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_374),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_435),
.Y(n_662)
);

INVx6_ASAP7_75t_L g663 ( 
.A(n_378),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_480),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_361),
.Y(n_665)
);

INVx6_ASAP7_75t_L g666 ( 
.A(n_378),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_491),
.Y(n_667)
);

CKINVDCx8_ASAP7_75t_R g668 ( 
.A(n_390),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_435),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_378),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_505),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_480),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_454),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_505),
.Y(n_674)
);

BUFx12f_ASAP7_75t_L g675 ( 
.A(n_362),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_590),
.B(n_405),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_600),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_612),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_633),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_633),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_637),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_514),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_655),
.Y(n_683)
);

NOR2x1p5_ASAP7_75t_L g684 ( 
.A(n_590),
.B(n_360),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_655),
.Y(n_685)
);

INVx11_ASAP7_75t_L g686 ( 
.A(n_634),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_612),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_591),
.B(n_584),
.C(n_571),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_631),
.B(n_636),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_631),
.B(n_551),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_636),
.B(n_645),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_633),
.Y(n_692)
);

INVx3_ASAP7_75t_L g693 ( 
.A(n_656),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_656),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_622),
.A2(n_449),
.B1(n_405),
.B2(n_560),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_656),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_638),
.B(n_378),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_595),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_595),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_637),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_638),
.B(n_378),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_597),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_650),
.B(n_561),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_617),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_602),
.B(n_378),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_617),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_640),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_632),
.B(n_369),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_638),
.B(n_497),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_650),
.B(n_561),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_617),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_648),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_648),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_638),
.B(n_497),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_617),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_648),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_638),
.B(n_497),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_664),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_643),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_664),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_622),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_622),
.Y(n_724)
);

INVxp33_ASAP7_75t_SL g725 ( 
.A(n_654),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_663),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_638),
.B(n_497),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_672),
.Y(n_728)
);

CKINVDCx11_ASAP7_75t_R g729 ( 
.A(n_668),
.Y(n_729)
);

BUFx6f_ASAP7_75t_SL g730 ( 
.A(n_650),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_611),
.B(n_618),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_675),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_611),
.B(n_497),
.Y(n_733)
);

INVxp67_ASAP7_75t_SL g734 ( 
.A(n_592),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_644),
.B(n_350),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_665),
.B(n_369),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_665),
.B(n_370),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_593),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_593),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_601),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_644),
.B(n_564),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_601),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_603),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_652),
.A2(n_449),
.B1(n_544),
.B2(n_372),
.Y(n_744)
);

AND2x2_ASAP7_75t_SL g745 ( 
.A(n_665),
.B(n_342),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_603),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_608),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_606),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_608),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_613),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_597),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_613),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_610),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_610),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_610),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_644),
.B(n_355),
.Y(n_756)
);

NOR2x1p5_ASAP7_75t_L g757 ( 
.A(n_634),
.B(n_372),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_610),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_663),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_610),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_663),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_619),
.B(n_620),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_610),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_614),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_675),
.Y(n_765)
);

INVx5_ASAP7_75t_L g766 ( 
.A(n_602),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_644),
.B(n_564),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_673),
.B(n_550),
.Y(n_768)
);

AO21x2_ASAP7_75t_L g769 ( 
.A1(n_587),
.A2(n_365),
.B(n_363),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_624),
.Y(n_770)
);

CKINVDCx6p67_ASAP7_75t_R g771 ( 
.A(n_673),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_624),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_592),
.B(n_535),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_SL g774 ( 
.A(n_646),
.B(n_353),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_635),
.B(n_366),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_594),
.B(n_556),
.C(n_555),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_614),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_373),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_614),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_615),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_589),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_670),
.B(n_556),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_615),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_615),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_626),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_624),
.Y(n_786)
);

OAI22xp33_ASAP7_75t_L g787 ( 
.A1(n_627),
.A2(n_569),
.B1(n_565),
.B2(n_524),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_670),
.B(n_569),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_663),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_630),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_670),
.B(n_362),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_668),
.B(n_380),
.Y(n_792)
);

AND2x2_ASAP7_75t_SL g793 ( 
.A(n_642),
.B(n_356),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_623),
.B(n_381),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_653),
.Y(n_795)
);

INVxp67_ASAP7_75t_SL g796 ( 
.A(n_621),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_597),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_L g798 ( 
.A(n_602),
.B(n_364),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_666),
.B(n_364),
.Y(n_799)
);

OAI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_639),
.A2(n_354),
.B1(n_387),
.B2(n_343),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_625),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_646),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_604),
.A2(n_353),
.B1(n_512),
.B2(n_412),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_667),
.B(n_535),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_625),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_621),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_689),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_728),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_804),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_689),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_676),
.B(n_596),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_704),
.B(n_711),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_734),
.B(n_721),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_736),
.B(n_609),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_691),
.B(n_545),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_804),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_711),
.B(n_546),
.Y(n_817)
);

OAI221xp5_ASAP7_75t_L g818 ( 
.A1(n_696),
.A2(n_627),
.B1(n_547),
.B2(n_580),
.C(n_496),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_737),
.B(n_554),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_699),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_700),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_766),
.B(n_558),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_682),
.B(n_671),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_677),
.B(n_388),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_730),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_690),
.B(n_674),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_741),
.B(n_563),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_745),
.B(n_607),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_L g829 ( 
.A1(n_678),
.A2(n_641),
.B1(n_621),
.B2(n_616),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_806),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_741),
.B(n_563),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_767),
.B(n_566),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_767),
.B(n_566),
.Y(n_833)
);

OR2x2_ASAP7_75t_SL g834 ( 
.A(n_729),
.B(n_598),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_773),
.B(n_602),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_806),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_685),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_676),
.B(n_607),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_686),
.Y(n_839)
);

NOR2xp67_ASAP7_75t_L g840 ( 
.A(n_683),
.B(n_649),
.Y(n_840)
);

NOR2xp67_ASAP7_75t_L g841 ( 
.A(n_683),
.B(n_651),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_782),
.B(n_616),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_744),
.B(n_798),
.C(n_776),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_788),
.B(n_616),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_676),
.B(n_598),
.Y(n_845)
);

NOR3xp33_ASAP7_75t_L g846 ( 
.A(n_787),
.B(n_376),
.C(n_398),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_745),
.B(n_616),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_687),
.A2(n_641),
.B1(n_659),
.B2(n_657),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_768),
.B(n_641),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_676),
.B(n_629),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_L g851 ( 
.A(n_800),
.B(n_403),
.C(n_402),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_709),
.B(n_408),
.Y(n_852)
);

NOR3xp33_ASAP7_75t_L g853 ( 
.A(n_774),
.B(n_419),
.C(n_411),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_795),
.Y(n_854)
);

AOI221xp5_ASAP7_75t_L g855 ( 
.A1(n_708),
.A2(n_367),
.B1(n_371),
.B2(n_358),
.C(n_349),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_735),
.B(n_756),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_709),
.B(n_424),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_793),
.B(n_344),
.Y(n_859)
);

INVxp33_ASAP7_75t_L g860 ( 
.A(n_785),
.Y(n_860)
);

BUFx5_ASAP7_75t_L g861 ( 
.A(n_789),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_793),
.B(n_345),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_796),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_717),
.B(n_346),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_732),
.B(n_431),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_694),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_717),
.B(n_352),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_730),
.Y(n_868)
);

NOR2xp67_ASAP7_75t_L g869 ( 
.A(n_688),
.B(n_660),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_715),
.B(n_432),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_681),
.B(n_379),
.Y(n_871)
);

NAND2xp33_ASAP7_75t_L g872 ( 
.A(n_697),
.B(n_393),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_720),
.B(n_385),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_701),
.B(n_394),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_701),
.B(n_791),
.Y(n_875)
);

NAND2xp33_ASAP7_75t_L g876 ( 
.A(n_693),
.B(n_395),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_693),
.A2(n_798),
.B1(n_706),
.B2(n_724),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_799),
.B(n_404),
.Y(n_878)
);

BUFx6f_ASAP7_75t_SL g879 ( 
.A(n_722),
.Y(n_879)
);

AO221x1_ASAP7_75t_L g880 ( 
.A1(n_774),
.A2(n_629),
.B1(n_504),
.B2(n_528),
.C(n_512),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_684),
.B(n_412),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_717),
.B(n_413),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_770),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_792),
.B(n_417),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_726),
.B(n_421),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_705),
.B(n_422),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_729),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_SL g888 ( 
.A(n_725),
.B(n_528),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_705),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_707),
.B(n_389),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_707),
.B(n_426),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_712),
.B(n_429),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_770),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_748),
.B(n_433),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_772),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_L g896 ( 
.A(n_726),
.B(n_436),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_712),
.B(n_439),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_803),
.A2(n_533),
.B1(n_575),
.B2(n_565),
.Y(n_898)
);

BUFx2_ASAP7_75t_R g899 ( 
.A(n_781),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_723),
.B(n_446),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_771),
.B(n_462),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_771),
.B(n_464),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_775),
.B(n_391),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_725),
.B(n_778),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_723),
.B(n_466),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_765),
.B(n_434),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_723),
.B(n_442),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_794),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_724),
.B(n_473),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_724),
.B(n_479),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_SL g911 ( 
.A(n_757),
.B(n_533),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_706),
.A2(n_661),
.B1(n_399),
.B2(n_407),
.Y(n_912)
);

NAND2xp33_ASAP7_75t_L g913 ( 
.A(n_759),
.B(n_484),
.Y(n_913)
);

OAI221xp5_ASAP7_75t_L g914 ( 
.A1(n_731),
.A2(n_416),
.B1(n_423),
.B2(n_410),
.C(n_392),
.Y(n_914)
);

INVx4_ASAP7_75t_SL g915 ( 
.A(n_759),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_786),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_790),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_790),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_L g919 ( 
.A(n_731),
.B(n_451),
.C(n_444),
.Y(n_919)
);

NOR2xp67_ASAP7_75t_L g920 ( 
.A(n_781),
.B(n_18),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_769),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_753),
.Y(n_922)
);

NAND2xp33_ASAP7_75t_L g923 ( 
.A(n_761),
.B(n_499),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_738),
.B(n_400),
.Y(n_924)
);

OR2x6_ASAP7_75t_L g925 ( 
.A(n_686),
.B(n_587),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_739),
.B(n_401),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_739),
.B(n_406),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_769),
.A2(n_438),
.B1(n_440),
.B2(n_430),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_762),
.Y(n_929)
);

INVxp33_ASAP7_75t_L g930 ( 
.A(n_802),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_740),
.B(n_511),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_733),
.B(n_414),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_733),
.B(n_415),
.Y(n_933)
);

NOR3xp33_ASAP7_75t_L g934 ( 
.A(n_762),
.B(n_455),
.C(n_453),
.Y(n_934)
);

OAI21xp33_ASAP7_75t_L g935 ( 
.A1(n_742),
.A2(n_578),
.B(n_574),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_769),
.A2(n_743),
.B1(n_746),
.B2(n_742),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_698),
.B(n_420),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_746),
.B(n_516),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_802),
.B(n_457),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_698),
.B(n_427),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_747),
.B(n_527),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_702),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_754),
.B(n_504),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_755),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_749),
.B(n_461),
.C(n_459),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_749),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_750),
.B(n_531),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_710),
.A2(n_468),
.B1(n_472),
.B2(n_465),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_750),
.B(n_576),
.Y(n_949)
);

NOR2x1p5_ASAP7_75t_L g950 ( 
.A(n_758),
.B(n_476),
.Y(n_950)
);

BUFx6f_ASAP7_75t_SL g951 ( 
.A(n_703),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_752),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_710),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_716),
.B(n_522),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_L g955 ( 
.A(n_716),
.B(n_481),
.C(n_478),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_719),
.B(n_582),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_760),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_727),
.B(n_574),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_760),
.B(n_428),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_763),
.A2(n_450),
.B(n_456),
.C(n_448),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_764),
.B(n_437),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_764),
.B(n_578),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_805),
.A2(n_492),
.B1(n_494),
.B2(n_482),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_777),
.B(n_518),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_801),
.B(n_508),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_779),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_801),
.B(n_513),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_779),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_780),
.B(n_447),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_780),
.B(n_452),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_783),
.B(n_523),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_783),
.B(n_529),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_784),
.B(n_463),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_849),
.A2(n_628),
.B(n_588),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_818),
.A2(n_846),
.B(n_914),
.C(n_810),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_829),
.A2(n_628),
.B(n_588),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_807),
.B(n_536),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_807),
.B(n_538),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_829),
.A2(n_628),
.B(n_588),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_810),
.B(n_539),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_904),
.B(n_811),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_823),
.B(n_540),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_813),
.B(n_575),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_863),
.A2(n_469),
.B1(n_477),
.B2(n_467),
.Y(n_984)
);

BUFx8_ASAP7_75t_SL g985 ( 
.A(n_887),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_823),
.B(n_577),
.Y(n_986)
);

OAI21xp33_ASAP7_75t_L g987 ( 
.A1(n_888),
.A2(n_586),
.B(n_585),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_946),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_852),
.B(n_483),
.Y(n_989)
);

NAND3xp33_ASAP7_75t_L g990 ( 
.A(n_851),
.B(n_647),
.C(n_489),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_853),
.A2(n_493),
.B1(n_495),
.B2(n_490),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_826),
.B(n_828),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_863),
.A2(n_500),
.B1(n_506),
.B2(n_498),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_828),
.B(n_507),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_811),
.B(n_509),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_866),
.B(n_515),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_842),
.A2(n_844),
.B(n_835),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_858),
.B(n_525),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_866),
.A2(n_532),
.B1(n_548),
.B2(n_543),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_809),
.B(n_816),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_846),
.A2(n_559),
.B(n_562),
.C(n_557),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_894),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_837),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_838),
.B(n_567),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_906),
.B(n_572),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_877),
.A2(n_581),
.B1(n_534),
.B2(n_518),
.Y(n_1006)
);

OAI21xp33_ASAP7_75t_L g1007 ( 
.A1(n_857),
.A2(n_534),
.B(n_501),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_838),
.B(n_435),
.Y(n_1008)
);

BUFx4f_ASAP7_75t_L g1009 ( 
.A(n_845),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_877),
.A2(n_475),
.B1(n_517),
.B2(n_510),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_847),
.A2(n_521),
.B1(n_530),
.B2(n_526),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_827),
.B(n_831),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_812),
.A2(n_542),
.B(n_552),
.C(n_549),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_853),
.A2(n_553),
.B(n_570),
.C(n_568),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_939),
.Y(n_1015)
);

BUFx12f_ASAP7_75t_L g1016 ( 
.A(n_834),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_824),
.A2(n_471),
.B1(n_680),
.B2(n_679),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_865),
.B(n_19),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_832),
.B(n_833),
.Y(n_1019)
);

AO21x1_ASAP7_75t_L g1020 ( 
.A1(n_890),
.A2(n_695),
.B(n_692),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_814),
.B(n_20),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_875),
.A2(n_695),
.B(n_692),
.Y(n_1022)
);

AOI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_843),
.A2(n_934),
.B1(n_870),
.B2(n_907),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_873),
.B(n_22),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_851),
.A2(n_714),
.B(n_718),
.C(n_713),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_848),
.A2(n_817),
.B(n_952),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_859),
.B(n_24),
.Y(n_1027)
);

NOR2x1p5_ASAP7_75t_L g1028 ( 
.A(n_881),
.B(n_24),
.Y(n_1028)
);

AND2x2_ASAP7_75t_SL g1029 ( 
.A(n_881),
.B(n_26),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_820),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_821),
.Y(n_1031)
);

AND3x1_ASAP7_75t_L g1032 ( 
.A(n_899),
.B(n_26),
.C(n_27),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_845),
.B(n_28),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_840),
.B(n_29),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_912),
.A2(n_825),
.B1(n_868),
.B2(n_856),
.Y(n_1035)
);

NOR3xp33_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_29),
.C(n_30),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_825),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_873),
.B(n_30),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_960),
.A2(n_35),
.B(n_31),
.C(n_32),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_903),
.B(n_32),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_930),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_903),
.B(n_36),
.Y(n_1042)
);

INVx3_ASAP7_75t_L g1043 ( 
.A(n_808),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_934),
.B(n_37),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_911),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_862),
.B(n_37),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_921),
.A2(n_936),
.B(n_929),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_839),
.B(n_40),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_856),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_936),
.A2(n_797),
.B(n_751),
.Y(n_1050)
);

AO21x1_ASAP7_75t_L g1051 ( 
.A1(n_890),
.A2(n_599),
.B(n_597),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_845),
.B(n_658),
.Y(n_1052)
);

BUFx4f_ASAP7_75t_L g1053 ( 
.A(n_850),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_SL g1054 ( 
.A(n_850),
.B(n_943),
.Y(n_1054)
);

OR2x2_ASAP7_75t_L g1055 ( 
.A(n_898),
.B(n_42),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_854),
.A2(n_46),
.B(n_44),
.C(n_45),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_850),
.B(n_46),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_868),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_830),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_884),
.B(n_905),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_879),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_964),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_889),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_958),
.A2(n_954),
.B(n_908),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_860),
.B(n_47),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_955),
.B(n_48),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_955),
.B(n_49),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_932),
.A2(n_662),
.B(n_669),
.C(n_658),
.Y(n_1068)
);

AO21x1_ASAP7_75t_L g1069 ( 
.A1(n_959),
.A2(n_599),
.B(n_597),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_910),
.B(n_819),
.Y(n_1070)
);

NAND2x2_ASAP7_75t_L g1071 ( 
.A(n_880),
.B(n_51),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_841),
.B(n_950),
.Y(n_1072)
);

O2A1O1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_855),
.A2(n_54),
.B(n_52),
.C(n_53),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_920),
.B(n_658),
.Y(n_1074)
);

BUFx4f_ASAP7_75t_L g1075 ( 
.A(n_925),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_932),
.A2(n_605),
.B(n_599),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_872),
.A2(n_924),
.B(n_927),
.C(n_926),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_933),
.A2(n_605),
.B(n_599),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_963),
.B(n_56),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_R g1080 ( 
.A(n_879),
.B(n_57),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_933),
.A2(n_605),
.B(n_662),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_928),
.A2(n_605),
.B(n_662),
.Y(n_1082)
);

NOR2x1p5_ASAP7_75t_L g1083 ( 
.A(n_919),
.B(n_945),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_948),
.B(n_59),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_883),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_926),
.A2(n_63),
.B(n_60),
.C(n_62),
.Y(n_1086)
);

NOR2xp67_ASAP7_75t_L g1087 ( 
.A(n_869),
.B(n_60),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_937),
.A2(n_669),
.B(n_65),
.C(n_62),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_940),
.A2(n_67),
.B(n_64),
.C(n_66),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_830),
.A2(n_212),
.B(n_208),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_900),
.B(n_67),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_861),
.B(n_68),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_815),
.B(n_69),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_876),
.B(n_73),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_964),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_836),
.A2(n_341),
.B(n_217),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_909),
.B(n_74),
.Y(n_1097)
);

AOI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_938),
.A2(n_75),
.B(n_76),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_964),
.Y(n_1099)
);

AND2x6_ASAP7_75t_SL g1100 ( 
.A(n_925),
.B(n_75),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_901),
.B(n_78),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_927),
.A2(n_81),
.B1(n_78),
.B2(n_79),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_942),
.A2(n_219),
.B(n_213),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_902),
.B(n_79),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_956),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_951),
.Y(n_1106)
);

OAI321xp33_ASAP7_75t_L g1107 ( 
.A1(n_935),
.A2(n_85),
.A3(n_86),
.B1(n_87),
.B2(n_88),
.C(n_89),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_836),
.A2(n_87),
.B1(n_89),
.B2(n_92),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_871),
.B(n_874),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_965),
.A2(n_340),
.B(n_224),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_953),
.A2(n_225),
.B(n_223),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_967),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_886),
.B(n_93),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_971),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_972),
.A2(n_337),
.B(n_230),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_969),
.A2(n_973),
.B(n_970),
.C(n_895),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_931),
.A2(n_94),
.B(n_95),
.C(n_96),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_893),
.Y(n_1118)
);

AO21x1_ASAP7_75t_L g1119 ( 
.A1(n_969),
.A2(n_98),
.B(n_99),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_916),
.A2(n_918),
.B(n_917),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_970),
.A2(n_99),
.B(n_100),
.C(n_101),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_941),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_944),
.Y(n_1123)
);

NOR2x1_ASAP7_75t_L g1124 ( 
.A(n_864),
.B(n_104),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_878),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_822),
.A2(n_336),
.B(n_235),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_973),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_922),
.A2(n_239),
.B(n_234),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_885),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_891),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_947),
.B(n_117),
.Y(n_1131)
);

AND2x2_ASAP7_75t_SL g1132 ( 
.A(n_896),
.B(n_118),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_949),
.B(n_867),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_962),
.A2(n_334),
.B(n_241),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_882),
.B(n_119),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_913),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_923),
.B(n_120),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_892),
.B(n_122),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_897),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_961),
.A2(n_333),
.B(n_243),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_915),
.B(n_123),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_915),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_966),
.A2(n_124),
.B(n_125),
.C(n_126),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_957),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_951),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_SL g1146 ( 
.A(n_968),
.B(n_126),
.Y(n_1146)
);

INVx4_ASAP7_75t_L g1147 ( 
.A(n_944),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_944),
.B(n_127),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_807),
.B(n_127),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_L g1150 ( 
.A(n_839),
.B(n_128),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1145),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1047),
.A2(n_129),
.B(n_130),
.Y(n_1152)
);

BUFx12f_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1020),
.A2(n_131),
.A3(n_132),
.B(n_133),
.Y(n_1154)
);

AND2x2_ASAP7_75t_L g1155 ( 
.A(n_983),
.B(n_132),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1000),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1030),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1031),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1047),
.A2(n_133),
.B(n_134),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1012),
.A2(n_134),
.B(n_135),
.C(n_136),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1130),
.B(n_136),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1037),
.B(n_137),
.Y(n_1162)
);

BUFx10_ASAP7_75t_L g1163 ( 
.A(n_1034),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1059),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1003),
.Y(n_1165)
);

NOR2x1_ASAP7_75t_SL g1166 ( 
.A(n_1035),
.B(n_138),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1049),
.B(n_138),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_981),
.B(n_140),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1001),
.A2(n_140),
.B1(n_143),
.B2(n_144),
.C(n_145),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1019),
.B(n_143),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1015),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_997),
.A2(n_145),
.B(n_146),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_975),
.B(n_147),
.Y(n_1173)
);

INVx8_ASAP7_75t_L g1174 ( 
.A(n_1106),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1075),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_1175)
);

AOI21xp33_ASAP7_75t_L g1176 ( 
.A1(n_1060),
.A2(n_148),
.B(n_149),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_1106),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1023),
.B(n_151),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1062),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_990),
.B(n_1025),
.C(n_1117),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_997),
.A2(n_152),
.B(n_154),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1058),
.B(n_155),
.Y(n_1182)
);

AOI221xp5_ASAP7_75t_L g1183 ( 
.A1(n_995),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.C(n_158),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1027),
.A2(n_157),
.B(n_158),
.C(n_159),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1082),
.A2(n_160),
.B(n_161),
.Y(n_1185)
);

INVx5_ASAP7_75t_L g1186 ( 
.A(n_1100),
.Y(n_1186)
);

AO31x2_ASAP7_75t_L g1187 ( 
.A1(n_1069),
.A2(n_160),
.A3(n_161),
.B(n_162),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1046),
.A2(n_164),
.B(n_165),
.C(n_167),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1052),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_982),
.B(n_167),
.Y(n_1190)
);

NOR2xp33_ASAP7_75t_L g1191 ( 
.A(n_1002),
.B(n_168),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1112),
.A2(n_168),
.B(n_169),
.C(n_170),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_SL g1193 ( 
.A(n_1061),
.B(n_169),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_986),
.B(n_170),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1082),
.A2(n_1064),
.B(n_1026),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_SL g1196 ( 
.A1(n_1029),
.A2(n_1054),
.B1(n_1132),
.B2(n_1045),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1040),
.A2(n_171),
.B(n_173),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_989),
.B(n_174),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_1028),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1042),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_1200)
);

NAND3x1_ASAP7_75t_L g1201 ( 
.A(n_1036),
.B(n_175),
.C(n_177),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1009),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_998),
.B(n_178),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_1139),
.B(n_178),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1055),
.B(n_1004),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1116),
.A2(n_179),
.B(n_181),
.Y(n_1206)
);

AND3x4_ASAP7_75t_L g1207 ( 
.A(n_1009),
.B(n_1053),
.C(n_985),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1063),
.B(n_179),
.Y(n_1208)
);

OR2x6_ASAP7_75t_L g1209 ( 
.A(n_1033),
.B(n_182),
.Y(n_1209)
);

A2O1A1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_1114),
.A2(n_183),
.B(n_249),
.C(n_250),
.Y(n_1210)
);

OA22x2_ASAP7_75t_L g1211 ( 
.A1(n_1057),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_1095),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1144),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1041),
.B(n_1005),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1065),
.Y(n_1215)
);

AND2x2_ASAP7_75t_SL g1216 ( 
.A(n_1032),
.B(n_300),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_987),
.B(n_1122),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1022),
.A2(n_1109),
.B(n_1120),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1081),
.A2(n_1078),
.B(n_1076),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_1099),
.Y(n_1220)
);

AOI21xp33_ASAP7_75t_L g1221 ( 
.A1(n_1039),
.A2(n_1038),
.B(n_1024),
.Y(n_1221)
);

AOI21xp33_ASAP7_75t_L g1222 ( 
.A1(n_1013),
.A2(n_1133),
.B(n_1077),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1119),
.A2(n_1068),
.A3(n_1115),
.B(n_1110),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_991),
.B(n_999),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1034),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1018),
.A2(n_1079),
.B1(n_1084),
.B2(n_984),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1021),
.A2(n_1127),
.B(n_1138),
.C(n_1014),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_996),
.B(n_994),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1073),
.A2(n_1105),
.B(n_1093),
.C(n_1056),
.Y(n_1229)
);

AO21x2_ASAP7_75t_L g1230 ( 
.A1(n_1103),
.A2(n_1111),
.B(n_1128),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1007),
.A2(n_1091),
.B(n_1131),
.C(n_1086),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1088),
.A2(n_1096),
.A3(n_1090),
.B(n_1006),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_977),
.B(n_978),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_993),
.B(n_980),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1146),
.B(n_1072),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1134),
.A2(n_1010),
.A3(n_1148),
.B(n_1121),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1080),
.B(n_1072),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1135),
.B(n_988),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1149),
.B(n_1083),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1113),
.B(n_1011),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1044),
.A2(n_1067),
.B(n_1066),
.Y(n_1241)
);

AND2x2_ASAP7_75t_SL g1242 ( 
.A(n_1141),
.B(n_1129),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1143),
.A2(n_1089),
.A3(n_1108),
.B(n_1126),
.Y(n_1243)
);

CKINVDCx8_ASAP7_75t_R g1244 ( 
.A(n_1048),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1059),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1101),
.B(n_1104),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1136),
.A2(n_1017),
.B1(n_1102),
.B2(n_1094),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1008),
.A2(n_1087),
.B1(n_1137),
.B2(n_1097),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1071),
.A2(n_1124),
.B1(n_1092),
.B2(n_1125),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1142),
.Y(n_1250)
);

NAND2x1_ASAP7_75t_L g1251 ( 
.A(n_1147),
.B(n_1043),
.Y(n_1251)
);

CKINVDCx16_ASAP7_75t_R g1252 ( 
.A(n_1074),
.Y(n_1252)
);

INVxp67_ASAP7_75t_L g1253 ( 
.A(n_1150),
.Y(n_1253)
);

INVx4_ASAP7_75t_L g1254 ( 
.A(n_1123),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1085),
.B(n_1118),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1098),
.B(n_1074),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1140),
.B(n_1107),
.Y(n_1257)
);

AOI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1036),
.A2(n_981),
.B1(n_1029),
.B2(n_745),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_992),
.B(n_981),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1020),
.A2(n_1069),
.A3(n_1051),
.B(n_1050),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_974),
.A2(n_979),
.B(n_976),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_981),
.B(n_725),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1003),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1047),
.A2(n_997),
.B(n_936),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_992),
.B(n_981),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1059),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1037),
.B(n_888),
.Y(n_1267)
);

BUFx4f_ASAP7_75t_L g1268 ( 
.A(n_1016),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_992),
.B(n_981),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1037),
.B(n_888),
.Y(n_1270)
);

AOI21xp33_ASAP7_75t_L g1271 ( 
.A1(n_1070),
.A2(n_904),
.B(n_930),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1047),
.A2(n_997),
.B(n_936),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_974),
.A2(n_979),
.B(n_976),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_974),
.A2(n_979),
.B(n_976),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1047),
.A2(n_997),
.B(n_936),
.Y(n_1275)
);

OA22x2_ASAP7_75t_L g1276 ( 
.A1(n_1033),
.A2(n_803),
.B1(n_850),
.B2(n_845),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_981),
.B(n_725),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1145),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_992),
.B(n_981),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_992),
.B(n_981),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1003),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_983),
.B(n_939),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_992),
.B(n_981),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1000),
.Y(n_1284)
);

OR2x6_ASAP7_75t_L g1285 ( 
.A(n_1016),
.B(n_845),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1030),
.Y(n_1286)
);

OAI22x1_ASAP7_75t_L g1287 ( 
.A1(n_1028),
.A2(n_803),
.B1(n_1055),
.B2(n_785),
.Y(n_1287)
);

NOR3xp33_ASAP7_75t_L g1288 ( 
.A(n_975),
.B(n_904),
.C(n_818),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_992),
.B(n_981),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1130),
.B(n_1139),
.Y(n_1290)
);

BUFx2_ASAP7_75t_L g1291 ( 
.A(n_1003),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_985),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_1037),
.B(n_888),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_992),
.B(n_981),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_985),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_992),
.B(n_981),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_992),
.B(n_981),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_981),
.B(n_725),
.Y(n_1298)
);

INVx5_ASAP7_75t_L g1299 ( 
.A(n_1106),
.Y(n_1299)
);

BUFx4f_ASAP7_75t_L g1300 ( 
.A(n_1016),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1145),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1130),
.B(n_1139),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1059),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1003),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1003),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_1037),
.B(n_888),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_992),
.B(n_981),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1020),
.A2(n_1069),
.A3(n_1051),
.B(n_1050),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1020),
.A2(n_1069),
.A3(n_1051),
.B(n_1050),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1145),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1130),
.B(n_1139),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_992),
.B(n_981),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_992),
.B(n_981),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1037),
.B(n_888),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1047),
.A2(n_997),
.B(n_936),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1145),
.Y(n_1316)
);

AO31x2_ASAP7_75t_L g1317 ( 
.A1(n_1020),
.A2(n_1069),
.A3(n_1051),
.B(n_1050),
.Y(n_1317)
);

OAI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1005),
.A2(n_1019),
.B(n_1012),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1059),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_981),
.B(n_725),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1207),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1318),
.B(n_1156),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1318),
.B(n_1284),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1213),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_1295),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1262),
.B(n_1277),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1288),
.B(n_1224),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_SL g1328 ( 
.A(n_1292),
.B(n_1268),
.Y(n_1328)
);

INVx5_ASAP7_75t_L g1329 ( 
.A(n_1164),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1285),
.B(n_1208),
.Y(n_1330)
);

AO21x1_ASAP7_75t_L g1331 ( 
.A1(n_1152),
.A2(n_1159),
.B(n_1206),
.Y(n_1331)
);

BUFx2_ASAP7_75t_R g1332 ( 
.A(n_1244),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_1161),
.Y(n_1333)
);

NAND2x1p5_ASAP7_75t_L g1334 ( 
.A(n_1302),
.B(n_1311),
.Y(n_1334)
);

BUFx2_ASAP7_75t_R g1335 ( 
.A(n_1267),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1172),
.A2(n_1181),
.B(n_1206),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_1153),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1298),
.B(n_1320),
.Y(n_1338)
);

OA21x2_ASAP7_75t_L g1339 ( 
.A1(n_1195),
.A2(n_1272),
.B(n_1264),
.Y(n_1339)
);

INVx4_ASAP7_75t_SL g1340 ( 
.A(n_1161),
.Y(n_1340)
);

BUFx2_ASAP7_75t_SL g1341 ( 
.A(n_1278),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1264),
.A2(n_1275),
.B(n_1272),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1157),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_SL g1344 ( 
.A1(n_1172),
.A2(n_1181),
.B(n_1166),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1271),
.B(n_1226),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1268),
.Y(n_1346)
);

NOR2xp67_ASAP7_75t_L g1347 ( 
.A(n_1186),
.B(n_1202),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1275),
.A2(n_1315),
.B(n_1219),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1230),
.A2(n_1218),
.B(n_1315),
.Y(n_1349)
);

INVx8_ASAP7_75t_L g1350 ( 
.A(n_1174),
.Y(n_1350)
);

BUFx8_ASAP7_75t_L g1351 ( 
.A(n_1199),
.Y(n_1351)
);

OR2x6_ASAP7_75t_L g1352 ( 
.A(n_1285),
.B(n_1204),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1304),
.Y(n_1353)
);

OR2x6_ASAP7_75t_L g1354 ( 
.A(n_1285),
.B(n_1204),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1240),
.A2(n_1258),
.B1(n_1196),
.B2(n_1225),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1286),
.B(n_1158),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1319),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1180),
.A2(n_1257),
.B(n_1230),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1300),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1152),
.A2(n_1159),
.B(n_1185),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1174),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1174),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1300),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1221),
.A2(n_1248),
.B(n_1227),
.Y(n_1364)
);

NAND3xp33_ASAP7_75t_L g1365 ( 
.A(n_1246),
.B(n_1210),
.C(n_1188),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1252),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1186),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1186),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1205),
.B(n_1214),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1258),
.B(n_1259),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1229),
.A2(n_1239),
.B(n_1241),
.C(n_1234),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1233),
.A2(n_1231),
.B(n_1228),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1245),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1265),
.B(n_1269),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1225),
.A2(n_1297),
.B1(n_1283),
.B2(n_1294),
.Y(n_1375)
);

INVx4_ASAP7_75t_L g1376 ( 
.A(n_1278),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1279),
.B(n_1280),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1289),
.B(n_1296),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1304),
.B(n_1155),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1307),
.B(n_1312),
.Y(n_1380)
);

AO21x2_ASAP7_75t_L g1381 ( 
.A1(n_1256),
.A2(n_1178),
.B(n_1173),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1281),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1291),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1305),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_SL g1385 ( 
.A1(n_1175),
.A2(n_1254),
.B(n_1200),
.Y(n_1385)
);

INVx4_ASAP7_75t_L g1386 ( 
.A(n_1316),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1276),
.A2(n_1242),
.B1(n_1287),
.B2(n_1313),
.Y(n_1387)
);

NAND3xp33_ASAP7_75t_L g1388 ( 
.A(n_1184),
.B(n_1160),
.C(n_1169),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1282),
.B(n_1171),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1220),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1222),
.A2(n_1192),
.B(n_1197),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1211),
.A2(n_1249),
.B(n_1251),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1168),
.A2(n_1209),
.B1(n_1170),
.B2(n_1189),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1249),
.A2(n_1247),
.B(n_1235),
.Y(n_1394)
);

AO21x2_ASAP7_75t_L g1395 ( 
.A1(n_1190),
.A2(n_1194),
.B(n_1197),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1260),
.A2(n_1308),
.B(n_1317),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1198),
.A2(n_1203),
.B(n_1191),
.Y(n_1397)
);

INVx1_ASAP7_75t_SL g1398 ( 
.A(n_1250),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1250),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1260),
.A2(n_1317),
.B(n_1308),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1238),
.B(n_1299),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1209),
.B(n_1165),
.Y(n_1402)
);

INVx1_ASAP7_75t_SL g1403 ( 
.A(n_1220),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1260),
.A2(n_1309),
.B(n_1308),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1215),
.B(n_1217),
.Y(n_1405)
);

AO21x2_ASAP7_75t_L g1406 ( 
.A1(n_1176),
.A2(n_1309),
.B(n_1317),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1299),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1309),
.A2(n_1200),
.B(n_1175),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1316),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1270),
.B(n_1314),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1162),
.A2(n_1167),
.B(n_1182),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1201),
.A2(n_1223),
.B(n_1232),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1223),
.A2(n_1232),
.B(n_1255),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1193),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1154),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1151),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1299),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1183),
.A2(n_1216),
.B(n_1306),
.C(n_1293),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1177),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1177),
.B(n_1237),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1209),
.B(n_1263),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_SL g1422 ( 
.A1(n_1163),
.A2(n_1310),
.B(n_1301),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_SL g1423 ( 
.A(n_1163),
.B(n_1179),
.Y(n_1423)
);

BUFx12f_ASAP7_75t_L g1424 ( 
.A(n_1266),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1187),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1212),
.B(n_1253),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1303),
.A2(n_1243),
.B(n_1236),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1288),
.A2(n_1036),
.B1(n_1318),
.B2(n_1029),
.Y(n_1428)
);

AO21x2_ASAP7_75t_L g1429 ( 
.A1(n_1261),
.A2(n_1274),
.B(n_1273),
.Y(n_1429)
);

BUFx2_ASAP7_75t_SL g1430 ( 
.A(n_1295),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1292),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1226),
.A2(n_1240),
.B1(n_1258),
.B2(n_1318),
.Y(n_1432)
);

AND2x4_ASAP7_75t_L g1433 ( 
.A(n_1290),
.B(n_1302),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1288),
.B(n_990),
.C(n_1246),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_SL g1435 ( 
.A1(n_1172),
.A2(n_1181),
.B(n_1206),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1292),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1290),
.Y(n_1437)
);

AO21x2_ASAP7_75t_L g1438 ( 
.A1(n_1261),
.A2(n_1274),
.B(n_1273),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1304),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1343),
.B(n_1374),
.Y(n_1440)
);

BUFx12f_ASAP7_75t_SL g1441 ( 
.A(n_1321),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1350),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1365),
.A2(n_1388),
.B(n_1434),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1343),
.B(n_1372),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1350),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1340),
.B(n_1333),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_SL g1449 ( 
.A1(n_1333),
.A2(n_1393),
.B1(n_1385),
.B2(n_1354),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1370),
.B(n_1356),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1432),
.B(n_1327),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1424),
.Y(n_1452)
);

OR2x6_ASAP7_75t_L g1453 ( 
.A(n_1352),
.B(n_1354),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1429),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1345),
.A2(n_1338),
.B1(n_1326),
.B2(n_1370),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1345),
.B(n_1369),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1438),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1424),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1322),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1350),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1438),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1326),
.B(n_1338),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_1373),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1418),
.A2(n_1428),
.B(n_1364),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1355),
.A2(n_1387),
.B1(n_1428),
.B2(n_1352),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1387),
.A2(n_1352),
.B1(n_1354),
.B2(n_1321),
.Y(n_1466)
);

AO21x2_ASAP7_75t_L g1467 ( 
.A1(n_1349),
.A2(n_1435),
.B(n_1336),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1353),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1330),
.A2(n_1334),
.B1(n_1366),
.B2(n_1423),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1330),
.A2(n_1375),
.B1(n_1433),
.B2(n_1331),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1390),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1390),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1439),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1324),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1359),
.Y(n_1475)
);

AO21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1323),
.A2(n_1344),
.B(n_1425),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1362),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1389),
.Y(n_1478)
);

INVx4_ASAP7_75t_L g1479 ( 
.A(n_1362),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1394),
.B(n_1379),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1359),
.A2(n_1363),
.B1(n_1399),
.B2(n_1409),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1415),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1394),
.B(n_1371),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1366),
.A2(n_1421),
.B1(n_1402),
.B2(n_1399),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1437),
.B(n_1404),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1409),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1414),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1405),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1426),
.Y(n_1489)
);

CKINVDCx11_ASAP7_75t_R g1490 ( 
.A(n_1363),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1410),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1382),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1410),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1403),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1329),
.B(n_1357),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1411),
.A2(n_1397),
.B1(n_1408),
.B2(n_1401),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1373),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1384),
.Y(n_1498)
);

INVx6_ASAP7_75t_L g1499 ( 
.A(n_1357),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1482),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1499),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1440),
.B(n_1383),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1482),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1451),
.B(n_1342),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1463),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1485),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1485),
.B(n_1413),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1495),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1480),
.B(n_1413),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.Y(n_1510)
);

AND2x4_ASAP7_75t_L g1511 ( 
.A(n_1480),
.B(n_1427),
.Y(n_1511)
);

INVx4_ASAP7_75t_L g1512 ( 
.A(n_1447),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1450),
.B(n_1412),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1450),
.B(n_1404),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1440),
.B(n_1398),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1445),
.B(n_1404),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1445),
.B(n_1342),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1492),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1468),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1451),
.B(n_1408),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1497),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1465),
.A2(n_1411),
.B1(n_1360),
.B2(n_1381),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1483),
.B(n_1342),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1495),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1483),
.B(n_1348),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1471),
.B(n_1339),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1464),
.B(n_1348),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1459),
.B(n_1339),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1455),
.A2(n_1360),
.B1(n_1381),
.B2(n_1395),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1473),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1497),
.Y(n_1531)
);

NOR2x1_ASAP7_75t_L g1532 ( 
.A(n_1469),
.B(n_1419),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1448),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1491),
.B(n_1339),
.Y(n_1534)
);

BUFx3_ASAP7_75t_L g1535 ( 
.A(n_1495),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1447),
.Y(n_1536)
);

OAI211xp5_ASAP7_75t_L g1537 ( 
.A1(n_1466),
.A2(n_1347),
.B(n_1386),
.C(n_1376),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1488),
.B(n_1420),
.Y(n_1538)
);

INVx4_ASAP7_75t_L g1539 ( 
.A(n_1447),
.Y(n_1539)
);

OR2x6_ASAP7_75t_L g1540 ( 
.A(n_1453),
.B(n_1392),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1493),
.B(n_1396),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1472),
.B(n_1396),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1499),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1462),
.A2(n_1395),
.B1(n_1420),
.B2(n_1391),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1467),
.B(n_1400),
.Y(n_1546)
);

OAI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1443),
.A2(n_1335),
.B(n_1392),
.Y(n_1547)
);

INVxp67_ASAP7_75t_R g1548 ( 
.A(n_1481),
.Y(n_1548)
);

BUFx4f_ASAP7_75t_SL g1549 ( 
.A(n_1460),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1456),
.B(n_1358),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1528),
.B(n_1496),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1528),
.B(n_1470),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1514),
.B(n_1454),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1514),
.B(n_1454),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1500),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1457),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1523),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1500),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1506),
.B(n_1525),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1510),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1503),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1521),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1509),
.B(n_1461),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1550),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1526),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1504),
.B(n_1478),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1531),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1527),
.B(n_1509),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1541),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1533),
.B(n_1486),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1508),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1541),
.Y(n_1572)
);

NOR2xp67_ASAP7_75t_L g1573 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1513),
.A2(n_1449),
.B1(n_1453),
.B2(n_1441),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1517),
.B(n_1476),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1517),
.B(n_1476),
.Y(n_1576)
);

INVx2_ASAP7_75t_SL g1577 ( 
.A(n_1512),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1504),
.B(n_1474),
.Y(n_1578)
);

NAND2xp33_ASAP7_75t_SL g1579 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1516),
.B(n_1406),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1536),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1564),
.B(n_1520),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1570),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1559),
.B(n_1519),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1564),
.B(n_1520),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1568),
.B(n_1513),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1555),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1568),
.B(n_1507),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1577),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1559),
.B(n_1530),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1507),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1557),
.B(n_1544),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1558),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1569),
.B(n_1505),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1557),
.B(n_1511),
.Y(n_1596)
);

NAND2x1p5_ASAP7_75t_L g1597 ( 
.A(n_1573),
.B(n_1532),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1563),
.B(n_1511),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1561),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1579),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1569),
.B(n_1516),
.Y(n_1602)
);

NAND2x1p5_ASAP7_75t_L g1603 ( 
.A(n_1573),
.B(n_1532),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1561),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1563),
.B(n_1511),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1566),
.B(n_1518),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1581),
.Y(n_1607)
);

AND2x4_ASAP7_75t_SL g1608 ( 
.A(n_1577),
.B(n_1512),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1566),
.B(n_1542),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1572),
.B(n_1511),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1553),
.B(n_1546),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1594),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1606),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1586),
.B(n_1554),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1594),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1601),
.B(n_1574),
.C(n_1484),
.D(n_1547),
.Y(n_1617)
);

INVx1_ASAP7_75t_SL g1618 ( 
.A(n_1608),
.Y(n_1618)
);

NAND2x1_ASAP7_75t_L g1619 ( 
.A(n_1589),
.B(n_1581),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1587),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1589),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1584),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1582),
.B(n_1572),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1565),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1599),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1600),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1588),
.B(n_1554),
.Y(n_1628)
);

NOR2xp67_ASAP7_75t_SL g1629 ( 
.A(n_1597),
.B(n_1537),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1588),
.B(n_1556),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1604),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1597),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1585),
.B(n_1580),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1585),
.B(n_1580),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1610),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1602),
.B(n_1578),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1602),
.B(n_1578),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1610),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1590),
.B(n_1593),
.Y(n_1639)
);

OAI32xp33_ASAP7_75t_L g1640 ( 
.A1(n_1618),
.A2(n_1603),
.A3(n_1597),
.B1(n_1607),
.B2(n_1583),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1619),
.A2(n_1603),
.B1(n_1548),
.B2(n_1577),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1636),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1636),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1619),
.B(n_1603),
.Y(n_1644)
);

INVx2_ASAP7_75t_SL g1645 ( 
.A(n_1637),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1637),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1632),
.A2(n_1608),
.B1(n_1548),
.B2(n_1539),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1639),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1624),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1617),
.A2(n_1576),
.B(n_1575),
.Y(n_1650)
);

OAI32xp33_ASAP7_75t_L g1651 ( 
.A1(n_1632),
.A2(n_1539),
.A3(n_1571),
.B1(n_1591),
.B2(n_1560),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1614),
.Y(n_1652)
);

OAI31xp33_ASAP7_75t_L g1653 ( 
.A1(n_1632),
.A2(n_1547),
.A3(n_1576),
.B(n_1575),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1629),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1621),
.B(n_1596),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1591),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1629),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1613),
.A2(n_1490),
.B(n_1475),
.C(n_1479),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1612),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1639),
.Y(n_1660)
);

AOI321xp33_ASAP7_75t_L g1661 ( 
.A1(n_1623),
.A2(n_1552),
.A3(n_1551),
.B1(n_1609),
.B2(n_1596),
.C(n_1545),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1622),
.A2(n_1508),
.B(n_1535),
.C(n_1524),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1612),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1633),
.A2(n_1552),
.B1(n_1453),
.B2(n_1538),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_L g1665 ( 
.A1(n_1654),
.A2(n_1633),
.B1(n_1634),
.B2(n_1635),
.C(n_1638),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1650),
.A2(n_1634),
.B(n_1635),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1654),
.A2(n_1567),
.B(n_1615),
.Y(n_1667)
);

OAI31xp33_ASAP7_75t_L g1668 ( 
.A1(n_1657),
.A2(n_1641),
.A3(n_1658),
.B(n_1653),
.Y(n_1668)
);

O2A1O1Ixp5_ASAP7_75t_L g1669 ( 
.A1(n_1658),
.A2(n_1640),
.B(n_1651),
.C(n_1647),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1657),
.A2(n_1638),
.B1(n_1605),
.B2(n_1598),
.Y(n_1670)
);

OAI32xp33_ASAP7_75t_L g1671 ( 
.A1(n_1648),
.A2(n_1630),
.A3(n_1628),
.B1(n_1615),
.B2(n_1539),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1659),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1644),
.A2(n_1549),
.B1(n_1539),
.B2(n_1508),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1663),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1661),
.A2(n_1652),
.B(n_1662),
.C(n_1660),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

AO22x2_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1667),
.B1(n_1674),
.B2(n_1672),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1649),
.Y(n_1678)
);

OAI21xp33_ASAP7_75t_L g1679 ( 
.A1(n_1666),
.A2(n_1664),
.B(n_1645),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1668),
.B(n_1656),
.Y(n_1680)
);

AOI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1671),
.A2(n_1644),
.B(n_1325),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_1643),
.Y(n_1682)
);

O2A1O1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1669),
.A2(n_1644),
.B(n_1328),
.C(n_1487),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1669),
.A2(n_1664),
.B(n_1646),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1673),
.A2(n_1655),
.B(n_1628),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_SL g1686 ( 
.A(n_1665),
.B(n_1368),
.C(n_1367),
.Y(n_1686)
);

NAND4xp25_ASAP7_75t_L g1687 ( 
.A(n_1668),
.B(n_1522),
.C(n_1444),
.D(n_1386),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1668),
.B(n_1655),
.Y(n_1688)
);

AOI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1668),
.A2(n_1494),
.B(n_1422),
.Y(n_1689)
);

AOI22x1_ASAP7_75t_L g1690 ( 
.A1(n_1668),
.A2(n_1430),
.B1(n_1337),
.B2(n_1431),
.Y(n_1690)
);

O2A1O1Ixp33_ASAP7_75t_L g1691 ( 
.A1(n_1675),
.A2(n_1489),
.B(n_1453),
.C(n_1477),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1688),
.B(n_1431),
.Y(n_1692)
);

NAND2x1_ASAP7_75t_L g1693 ( 
.A(n_1677),
.B(n_1630),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1680),
.B(n_1620),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1625),
.Y(n_1695)
);

OAI322xp33_ASAP7_75t_L g1696 ( 
.A1(n_1690),
.A2(n_1562),
.A3(n_1567),
.B1(n_1626),
.B2(n_1631),
.C1(n_1627),
.C2(n_1595),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1682),
.Y(n_1697)
);

NAND4xp25_ASAP7_75t_L g1698 ( 
.A(n_1687),
.B(n_1376),
.C(n_1460),
.D(n_1529),
.Y(n_1698)
);

NAND4xp25_ASAP7_75t_L g1699 ( 
.A(n_1683),
.B(n_1691),
.C(n_1689),
.D(n_1684),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1681),
.B(n_1436),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1679),
.B(n_1436),
.Y(n_1701)
);

NOR3xp33_ASAP7_75t_L g1702 ( 
.A(n_1686),
.B(n_1337),
.C(n_1475),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1685),
.A2(n_1477),
.B(n_1460),
.Y(n_1703)
);

NOR2x1_ASAP7_75t_L g1704 ( 
.A(n_1700),
.B(n_1341),
.Y(n_1704)
);

NOR3xp33_ASAP7_75t_L g1705 ( 
.A(n_1699),
.B(n_1490),
.C(n_1346),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1698),
.A2(n_1346),
.B(n_1368),
.C(n_1367),
.Y(n_1706)
);

NOR3x1_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1677),
.C(n_1351),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1701),
.A2(n_1442),
.B(n_1446),
.C(n_1417),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1695),
.B(n_1598),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1692),
.A2(n_1540),
.B1(n_1502),
.B2(n_1562),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1694),
.B(n_1351),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1703),
.B(n_1605),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1693),
.A2(n_1540),
.B1(n_1535),
.B2(n_1524),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1696),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1714),
.B(n_1702),
.Y(n_1715)
);

NOR3xp33_ASAP7_75t_L g1716 ( 
.A(n_1705),
.B(n_1458),
.C(n_1452),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1711),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1708),
.Y(n_1718)
);

INVxp67_ASAP7_75t_SL g1719 ( 
.A(n_1704),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1709),
.B(n_1616),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1706),
.B(n_1351),
.C(n_1332),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1712),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1707),
.B(n_1611),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1710),
.B(n_1616),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_L g1725 ( 
.A(n_1713),
.B(n_1407),
.C(n_1452),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1714),
.B(n_1611),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1717),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_SL g1728 ( 
.A(n_1723),
.B(n_1442),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1715),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1721),
.B(n_1452),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1718),
.Y(n_1731)
);

NOR2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1719),
.B(n_1416),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1727),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1727),
.Y(n_1734)
);

AND4x1_ASAP7_75t_L g1735 ( 
.A(n_1730),
.B(n_1716),
.C(n_1725),
.D(n_1722),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1731),
.B(n_1726),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1729),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1737),
.Y(n_1738)
);

OA22x2_ASAP7_75t_L g1739 ( 
.A1(n_1736),
.A2(n_1732),
.B1(n_1728),
.B2(n_1724),
.Y(n_1739)
);

AND4x1_ASAP7_75t_L g1740 ( 
.A(n_1739),
.B(n_1734),
.C(n_1733),
.D(n_1721),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1738),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1741),
.A2(n_1738),
.B1(n_1733),
.B2(n_1720),
.Y(n_1742)
);

OAI21xp33_ASAP7_75t_L g1743 ( 
.A1(n_1740),
.A2(n_1735),
.B(n_1458),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1742),
.B(n_1446),
.Y(n_1744)
);

AOI22x1_ASAP7_75t_L g1745 ( 
.A1(n_1743),
.A2(n_1416),
.B1(n_1361),
.B2(n_1458),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1407),
.B(n_1419),
.Y(n_1746)
);

OAI21xp33_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1745),
.B(n_1515),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1747),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1441),
.B1(n_1543),
.B2(n_1501),
.Y(n_1749)
);


endmodule