module real_aes_10461_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_1004;
wire n_580;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_265;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_249;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_1049;
wire n_466;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_1352;
wire n_729;
wire n_394;
wire n_1323;
wire n_1280;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVxp33_ASAP7_75t_L g285 ( .A(n_0), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_0), .A2(n_233), .B1(n_386), .B2(n_391), .Y(n_385) );
OAI222xp33_ASAP7_75t_L g637 ( .A1(n_1), .A2(n_37), .B1(n_140), .B2(n_638), .C1(n_640), .C2(n_642), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_1), .A2(n_140), .B1(n_678), .B2(n_680), .C(n_681), .Y(n_677) );
INVx1_ASAP7_75t_L g1090 ( .A(n_2), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_3), .A2(n_214), .B1(n_392), .B2(n_499), .Y(n_873) );
INVxp33_ASAP7_75t_L g893 ( .A(n_3), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_4), .A2(n_16), .B1(n_322), .B2(n_565), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_4), .A2(n_16), .B1(n_498), .B2(n_606), .Y(n_731) );
INVx1_ASAP7_75t_L g913 ( .A(n_5), .Y(n_913) );
INVxp67_ASAP7_75t_SL g803 ( .A(n_6), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_6), .A2(n_203), .B1(n_391), .B2(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_7), .A2(n_166), .B1(n_486), .B2(n_718), .Y(n_980) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_7), .A2(n_118), .B1(n_287), .B2(n_322), .C(n_1004), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_8), .Y(n_247) );
AND2x2_ASAP7_75t_L g272 ( .A(n_8), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_8), .B(n_187), .Y(n_301) );
INVx1_ASAP7_75t_L g353 ( .A(n_8), .Y(n_353) );
INVx1_ASAP7_75t_L g544 ( .A(n_9), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_9), .A2(n_177), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_10), .A2(n_17), .B1(n_936), .B2(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g962 ( .A(n_10), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g568 ( .A1(n_11), .A2(n_45), .B1(n_564), .B2(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g610 ( .A(n_11), .Y(n_610) );
INVxp67_ASAP7_75t_L g320 ( .A(n_12), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_12), .A2(n_79), .B1(n_391), .B2(n_418), .Y(n_417) );
OA22x2_ASAP7_75t_L g1009 ( .A1(n_13), .A2(n_1010), .B1(n_1071), .B2(n_1072), .Y(n_1009) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_13), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_14), .A2(n_96), .B1(n_392), .B2(n_720), .Y(n_989) );
INVx1_ASAP7_75t_L g998 ( .A(n_14), .Y(n_998) );
OAI332xp33_ASAP7_75t_L g1019 ( .A1(n_15), .A2(n_309), .A3(n_349), .B1(n_1020), .B2(n_1023), .B3(n_1028), .C1(n_1031), .C2(n_1035), .Y(n_1019) );
INVx1_ASAP7_75t_L g1069 ( .A(n_15), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g957 ( .A1(n_17), .A2(n_103), .B1(n_958), .B2(n_959), .C(n_961), .Y(n_957) );
INVx1_ASAP7_75t_L g1189 ( .A(n_18), .Y(n_1189) );
INVx1_ASAP7_75t_L g751 ( .A(n_19), .Y(n_751) );
INVxp67_ASAP7_75t_L g799 ( .A(n_20), .Y(n_799) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_20), .A2(n_141), .B1(n_411), .B2(n_414), .C(n_835), .Y(n_834) );
AO221x2_ASAP7_75t_L g1116 ( .A1(n_21), .A2(n_51), .B1(n_1088), .B2(n_1107), .C(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1135 ( .A(n_22), .Y(n_1135) );
INVx1_ASAP7_75t_L g512 ( .A(n_23), .Y(n_512) );
INVxp33_ASAP7_75t_L g829 ( .A(n_24), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_24), .A2(n_93), .B1(n_841), .B2(n_842), .Y(n_840) );
INVx2_ASAP7_75t_L g366 ( .A(n_25), .Y(n_366) );
OR2x2_ASAP7_75t_L g397 ( .A(n_25), .B(n_364), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_26), .A2(n_99), .B1(n_742), .B2(n_743), .Y(n_741) );
OAI221xp5_ASAP7_75t_L g784 ( .A1(n_26), .A2(n_99), .B1(n_293), .B2(n_785), .C(n_786), .Y(n_784) );
INVx1_ASAP7_75t_L g1118 ( .A(n_27), .Y(n_1118) );
INVx1_ASAP7_75t_L g1311 ( .A(n_28), .Y(n_1311) );
CKINVDCx5p33_ASAP7_75t_R g1022 ( .A(n_29), .Y(n_1022) );
INVx1_ASAP7_75t_L g271 ( .A(n_30), .Y(n_271) );
OR2x2_ASAP7_75t_L g300 ( .A(n_30), .B(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g312 ( .A(n_30), .Y(n_312) );
BUFx2_ASAP7_75t_L g360 ( .A(n_30), .Y(n_360) );
INVxp33_ASAP7_75t_L g828 ( .A(n_31), .Y(n_828) );
AOI21xp33_ASAP7_75t_L g846 ( .A1(n_31), .A2(n_379), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g1187 ( .A(n_32), .Y(n_1187) );
INVx1_ASAP7_75t_L g764 ( .A(n_33), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g969 ( .A1(n_34), .A2(n_134), .B1(n_517), .B2(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_34), .A2(n_125), .B1(n_572), .B2(n_949), .Y(n_1002) );
INVx1_ASAP7_75t_L g812 ( .A(n_35), .Y(n_812) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_36), .A2(n_76), .B1(n_561), .B2(n_691), .Y(n_696) );
INVx1_ASAP7_75t_L g730 ( .A(n_36), .Y(n_730) );
INVx1_ASAP7_75t_L g682 ( .A(n_37), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_38), .A2(n_103), .B1(n_410), .B2(n_414), .C(n_759), .Y(n_934) );
INVx1_ASAP7_75t_L g963 ( .A(n_38), .Y(n_963) );
CKINVDCx16_ASAP7_75t_R g918 ( .A(n_39), .Y(n_918) );
INVx1_ASAP7_75t_L g1183 ( .A(n_40), .Y(n_1183) );
OAI221xp5_ASAP7_75t_SL g869 ( .A1(n_41), .A2(n_209), .B1(n_743), .B2(n_870), .C(n_871), .Y(n_869) );
OAI221xp5_ASAP7_75t_L g898 ( .A1(n_41), .A2(n_209), .B1(n_303), .B2(n_899), .C(n_900), .Y(n_898) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_42), .Y(n_865) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_43), .A2(n_195), .B1(n_561), .B2(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_43), .A2(n_154), .B1(n_717), .B2(n_718), .Y(n_716) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_44), .A2(n_132), .B1(n_879), .B2(n_881), .C(n_884), .Y(n_878) );
INVxp67_ASAP7_75t_SL g908 ( .A(n_44), .Y(n_908) );
INVx1_ASAP7_75t_L g579 ( .A(n_45), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_46), .A2(n_181), .B1(n_627), .B2(n_761), .Y(n_760) );
INVxp67_ASAP7_75t_SL g770 ( .A(n_46), .Y(n_770) );
AOI221xp5_ASAP7_75t_SL g931 ( .A1(n_47), .A2(n_70), .B1(n_379), .B2(n_382), .C(n_623), .Y(n_931) );
INVx1_ASAP7_75t_L g950 ( .A(n_47), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_48), .A2(n_90), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_48), .A2(n_173), .B1(n_391), .B2(n_632), .Y(n_1339) );
INVx1_ASAP7_75t_L g928 ( .A(n_49), .Y(n_928) );
INVx1_ASAP7_75t_L g757 ( .A(n_50), .Y(n_757) );
XNOR2x2_ASAP7_75t_L g683 ( .A(n_51), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g927 ( .A(n_52), .Y(n_927) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_53), .Y(n_1030) );
INVx1_ASAP7_75t_L g877 ( .A(n_54), .Y(n_877) );
INVxp33_ASAP7_75t_L g826 ( .A(n_55), .Y(n_826) );
NAND2xp33_ASAP7_75t_SL g844 ( .A(n_55), .B(n_845), .Y(n_844) );
OAI222xp33_ASAP7_75t_L g644 ( .A1(n_56), .A2(n_122), .B1(n_194), .B2(n_645), .C1(n_646), .C2(n_648), .Y(n_644) );
INVx1_ASAP7_75t_L g654 ( .A(n_56), .Y(n_654) );
INVx1_ASAP7_75t_L g1146 ( .A(n_57), .Y(n_1146) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_58), .A2(n_154), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_58), .A2(n_495), .B(n_720), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g744 ( .A1(n_59), .A2(n_207), .B1(n_745), .B2(n_747), .C(n_749), .Y(n_744) );
INVxp33_ASAP7_75t_L g792 ( .A(n_59), .Y(n_792) );
INVx1_ASAP7_75t_L g737 ( .A(n_60), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_61), .A2(n_185), .B1(n_1013), .B2(n_1014), .Y(n_1012) );
CKINVDCx5p33_ASAP7_75t_R g1067 ( .A(n_61), .Y(n_1067) );
INVxp33_ASAP7_75t_SL g444 ( .A(n_62), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g496 ( .A1(n_62), .A2(n_224), .B1(n_482), .B2(n_497), .C(n_500), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_63), .A2(n_123), .B1(n_391), .B2(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g673 ( .A(n_63), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_64), .A2(n_86), .B1(n_626), .B2(n_627), .Y(n_625) );
INVx1_ASAP7_75t_L g660 ( .A(n_64), .Y(n_660) );
CKINVDCx16_ASAP7_75t_R g1151 ( .A(n_65), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g973 ( .A(n_66), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_67), .A2(n_199), .B1(n_560), .B2(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g593 ( .A(n_67), .Y(n_593) );
INVx1_ASAP7_75t_L g852 ( .A(n_68), .Y(n_852) );
INVxp67_ASAP7_75t_L g314 ( .A(n_69), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_69), .A2(n_160), .B1(n_410), .B2(n_411), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g948 ( .A(n_70), .Y(n_948) );
XOR2x2_ASAP7_75t_L g965 ( .A(n_71), .B(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g553 ( .A(n_72), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_72), .A2(n_94), .B1(n_482), .B2(n_585), .C(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g1096 ( .A(n_73), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g922 ( .A1(n_74), .A2(n_204), .B1(n_923), .B2(n_924), .C(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g955 ( .A(n_74), .Y(n_955) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_75), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_76), .B(n_427), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g1015 ( .A1(n_77), .A2(n_127), .B1(n_357), .B2(n_1016), .Y(n_1015) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_77), .Y(n_1065) );
INVx1_ASAP7_75t_L g708 ( .A(n_78), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_78), .A2(n_114), .B1(n_718), .B2(n_720), .Y(n_724) );
INVxp67_ASAP7_75t_L g326 ( .A(n_79), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g821 ( .A1(n_80), .A2(n_152), .B1(n_293), .B2(n_302), .C(n_786), .Y(n_821) );
INVx1_ASAP7_75t_L g848 ( .A(n_80), .Y(n_848) );
CKINVDCx16_ASAP7_75t_R g1153 ( .A(n_81), .Y(n_1153) );
INVx1_ASAP7_75t_L g889 ( .A(n_82), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_83), .A2(n_124), .B1(n_1101), .B2(n_1104), .Y(n_1113) );
INVx1_ASAP7_75t_L g364 ( .A(n_84), .Y(n_364) );
INVx1_ASAP7_75t_L g384 ( .A(n_84), .Y(n_384) );
INVx1_ASAP7_75t_L g700 ( .A(n_85), .Y(n_700) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_85), .A2(n_486), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g656 ( .A(n_86), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g292 ( .A1(n_87), .A2(n_106), .B1(n_293), .B2(n_302), .C(n_306), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_87), .A2(n_106), .B1(n_399), .B2(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g926 ( .A(n_88), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g951 ( .A1(n_88), .A2(n_204), .B1(n_668), .B2(n_952), .C(n_954), .Y(n_951) );
INVx1_ASAP7_75t_L g1343 ( .A(n_89), .Y(n_1343) );
AOI221xp5_ASAP7_75t_L g1337 ( .A1(n_90), .A2(n_155), .B1(n_414), .B2(n_623), .C(n_1338), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_91), .A2(n_219), .B1(n_1319), .B2(n_1325), .Y(n_1324) );
INVxp67_ASAP7_75t_L g1336 ( .A(n_91), .Y(n_1336) );
INVxp33_ASAP7_75t_SL g1313 ( .A(n_92), .Y(n_1313) );
AOI21xp33_ASAP7_75t_L g1334 ( .A1(n_92), .A2(n_589), .B(n_717), .Y(n_1334) );
INVxp33_ASAP7_75t_L g824 ( .A(n_93), .Y(n_824) );
INVx1_ASAP7_75t_L g548 ( .A(n_94), .Y(n_548) );
INVx1_ASAP7_75t_L g1134 ( .A(n_95), .Y(n_1134) );
OAI211xp5_ASAP7_75t_L g992 ( .A1(n_96), .A2(n_993), .B(n_994), .C(n_996), .Y(n_992) );
INVx1_ASAP7_75t_L g939 ( .A(n_97), .Y(n_939) );
AO221x2_ASAP7_75t_L g1081 ( .A1(n_98), .A2(n_169), .B1(n_1082), .B2(n_1088), .C(n_1089), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_100), .A2(n_144), .B1(n_643), .B2(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g909 ( .A(n_100), .Y(n_909) );
INVx1_ASAP7_75t_L g239 ( .A(n_101), .Y(n_239) );
INVx1_ASAP7_75t_L g815 ( .A(n_102), .Y(n_815) );
INVx1_ASAP7_75t_L g463 ( .A(n_104), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_104), .A2(n_189), .B1(n_482), .B2(n_484), .C(n_487), .Y(n_481) );
XNOR2x1_ASAP7_75t_L g259 ( .A(n_105), .B(n_260), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g986 ( .A(n_107), .Y(n_986) );
INVxp67_ASAP7_75t_SL g1307 ( .A(n_108), .Y(n_1307) );
OAI221xp5_ASAP7_75t_L g1331 ( .A1(n_108), .A2(n_179), .B1(n_404), .B2(n_870), .C(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g335 ( .A(n_109), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_110), .A2(n_161), .B1(n_1088), .B2(n_1107), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_111), .A2(n_129), .B1(n_564), .B2(n_566), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g594 ( .A1(n_111), .A2(n_188), .B1(n_495), .B2(n_595), .C(n_597), .Y(n_594) );
AOI22xp33_ASAP7_75t_SL g1322 ( .A1(n_112), .A2(n_202), .B1(n_1321), .B2(n_1323), .Y(n_1322) );
INVxp33_ASAP7_75t_L g1342 ( .A(n_112), .Y(n_1342) );
INVx1_ASAP7_75t_L g514 ( .A(n_113), .Y(n_514) );
INVx1_ASAP7_75t_L g704 ( .A(n_114), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_115), .A2(n_164), .B1(n_411), .B2(n_495), .C(n_630), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_115), .A2(n_123), .B1(n_668), .B2(n_670), .C(n_672), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g1018 ( .A1(n_116), .A2(n_206), .B1(n_785), .B2(n_786), .C(n_899), .Y(n_1018) );
OAI222xp33_ASAP7_75t_L g1048 ( .A1(n_116), .A2(n_127), .B1(n_206), .B2(n_645), .C1(n_1049), .C2(n_1050), .Y(n_1048) );
INVx1_ASAP7_75t_L g818 ( .A(n_117), .Y(n_818) );
AOI21xp33_ASAP7_75t_L g981 ( .A1(n_118), .A2(n_595), .B(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1119 ( .A(n_119), .Y(n_1119) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_120), .A2(n_131), .B1(n_379), .B2(n_382), .C(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g658 ( .A(n_120), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_121), .A2(n_188), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_121), .A2(n_129), .B1(n_602), .B2(n_605), .Y(n_601) );
INVx1_ASAP7_75t_L g662 ( .A(n_122), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g971 ( .A1(n_125), .A2(n_137), .B1(n_523), .B2(n_628), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_126), .A2(n_197), .B1(n_282), .B2(n_478), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_126), .A2(n_216), .B1(n_517), .B2(n_519), .Y(n_516) );
INVx1_ASAP7_75t_L g346 ( .A(n_128), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_130), .Y(n_687) );
INVx1_ASAP7_75t_L g666 ( .A(n_131), .Y(n_666) );
INVx1_ASAP7_75t_L g906 ( .A(n_132), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g990 ( .A1(n_133), .A2(n_508), .B(n_991), .Y(n_990) );
INVx1_ASAP7_75t_L g997 ( .A(n_133), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g1001 ( .A1(n_134), .A2(n_137), .B1(n_266), .B2(n_693), .Y(n_1001) );
INVxp33_ASAP7_75t_SL g1314 ( .A(n_135), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_135), .A2(n_190), .B1(n_392), .B2(n_493), .Y(n_1333) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_136), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g1123 ( .A1(n_138), .A2(n_148), .B1(n_1101), .B2(n_1104), .Y(n_1123) );
AOI22xp5_ASAP7_75t_L g1353 ( .A1(n_139), .A2(n_1304), .B1(n_1354), .B2(n_1355), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g1354 ( .A(n_139), .Y(n_1354) );
INVxp33_ASAP7_75t_L g808 ( .A(n_141), .Y(n_808) );
INVx1_ASAP7_75t_L g453 ( .A(n_142), .Y(n_453) );
INVx1_ASAP7_75t_L g872 ( .A(n_143), .Y(n_872) );
INVx1_ASAP7_75t_L g905 ( .A(n_144), .Y(n_905) );
INVx1_ASAP7_75t_L g576 ( .A(n_145), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_146), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_147), .A2(n_225), .B1(n_410), .B2(n_414), .C(n_759), .Y(n_758) );
INVxp33_ASAP7_75t_SL g777 ( .A(n_147), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g1124 ( .A1(n_149), .A2(n_193), .B1(n_1082), .B2(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g740 ( .A(n_150), .Y(n_740) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_151), .Y(n_241) );
AND3x2_ASAP7_75t_L g1086 ( .A(n_151), .B(n_239), .C(n_1087), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1093 ( .A(n_151), .B(n_239), .Y(n_1093) );
INVx1_ASAP7_75t_L g849 ( .A(n_152), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g979 ( .A(n_153), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_155), .A2(n_173), .B1(n_569), .B2(n_1321), .Y(n_1320) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_156), .A2(n_200), .B1(n_523), .B2(n_976), .C(n_977), .Y(n_975) );
INVx1_ASAP7_75t_L g995 ( .A(n_156), .Y(n_995) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_157), .Y(n_1029) );
INVx2_ASAP7_75t_L g252 ( .A(n_158), .Y(n_252) );
XOR2xp5_ASAP7_75t_L g734 ( .A(n_159), .B(n_735), .Y(n_734) );
INVxp33_ASAP7_75t_L g333 ( .A(n_160), .Y(n_333) );
XNOR2x2_ASAP7_75t_L g440 ( .A(n_161), .B(n_441), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_162), .Y(n_550) );
INVx1_ASAP7_75t_L g752 ( .A(n_163), .Y(n_752) );
INVx1_ASAP7_75t_L g675 ( .A(n_164), .Y(n_675) );
INVx1_ASAP7_75t_L g929 ( .A(n_165), .Y(n_929) );
INVx1_ASAP7_75t_L g1005 ( .A(n_166), .Y(n_1005) );
CKINVDCx5p33_ASAP7_75t_R g1032 ( .A(n_167), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_168), .A2(n_172), .B1(n_1088), .B2(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g338 ( .A(n_170), .Y(n_338) );
INVx1_ASAP7_75t_L g1087 ( .A(n_171), .Y(n_1087) );
INVx1_ASAP7_75t_L g459 ( .A(n_174), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g1131 ( .A(n_175), .Y(n_1131) );
INVx1_ASAP7_75t_L g446 ( .A(n_176), .Y(n_446) );
INVx1_ASAP7_75t_L g545 ( .A(n_177), .Y(n_545) );
INVx1_ASAP7_75t_L g1185 ( .A(n_178), .Y(n_1185) );
XNOR2x1_ASAP7_75t_L g1303 ( .A(n_178), .B(n_1304), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_178), .A2(n_1350), .B1(n_1352), .B2(n_1356), .Y(n_1349) );
INVxp67_ASAP7_75t_SL g1308 ( .A(n_179), .Y(n_1308) );
AOI22x1_ASAP7_75t_L g793 ( .A1(n_180), .A2(n_794), .B1(n_795), .B2(n_853), .Y(n_793) );
INVx1_ASAP7_75t_L g853 ( .A(n_180), .Y(n_853) );
INVxp33_ASAP7_75t_L g774 ( .A(n_181), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g1021 ( .A(n_182), .Y(n_1021) );
INVx1_ASAP7_75t_L g765 ( .A(n_183), .Y(n_765) );
INVx1_ASAP7_75t_L g709 ( .A(n_184), .Y(n_709) );
OAI211xp5_ASAP7_75t_L g728 ( .A1(n_184), .A2(n_645), .B(n_729), .C(n_732), .Y(n_728) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_185), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_186), .Y(n_1033) );
INVx1_ASAP7_75t_L g254 ( .A(n_187), .Y(n_254) );
INVx2_ASAP7_75t_L g273 ( .A(n_187), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_189), .A2(n_192), .B1(n_465), .B2(n_468), .Y(n_464) );
INVxp33_ASAP7_75t_SL g1310 ( .A(n_190), .Y(n_1310) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_191), .A2(n_215), .B1(n_1101), .B2(n_1104), .Y(n_1100) );
INVx1_ASAP7_75t_L g491 ( .A(n_192), .Y(n_491) );
INVx1_ASAP7_75t_L g653 ( .A(n_194), .Y(n_653) );
INVx1_ASAP7_75t_L g714 ( .A(n_195), .Y(n_714) );
INVxp33_ASAP7_75t_L g280 ( .A(n_196), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_196), .A2(n_201), .B1(n_376), .B2(n_379), .C(n_382), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g521 ( .A1(n_197), .A2(n_220), .B1(n_522), .B2(n_523), .Y(n_521) );
XOR2x1_ASAP7_75t_L g540 ( .A(n_198), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g609 ( .A(n_199), .Y(n_609) );
INVx1_ASAP7_75t_L g1008 ( .A(n_200), .Y(n_1008) );
INVxp33_ASAP7_75t_L g274 ( .A(n_201), .Y(n_274) );
INVxp67_ASAP7_75t_L g1330 ( .A(n_202), .Y(n_1330) );
INVxp33_ASAP7_75t_L g805 ( .A(n_203), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_205), .A2(n_217), .B1(n_585), .B2(n_745), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g944 ( .A1(n_205), .A2(n_217), .B1(n_945), .B2(n_946), .C(n_947), .Y(n_944) );
INVxp33_ASAP7_75t_L g789 ( .A(n_207), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_208), .Y(n_1026) );
INVx1_ASAP7_75t_L g1147 ( .A(n_210), .Y(n_1147) );
INVx1_ASAP7_75t_L g342 ( .A(n_211), .Y(n_342) );
INVx1_ASAP7_75t_L g1085 ( .A(n_212), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_212), .B(n_1095), .Y(n_1098) );
AOI21xp33_ASAP7_75t_L g874 ( .A1(n_213), .A2(n_382), .B(n_875), .Y(n_874) );
INVxp33_ASAP7_75t_L g896 ( .A(n_213), .Y(n_896) );
INVxp33_ASAP7_75t_L g897 ( .A(n_214), .Y(n_897) );
INVxp67_ASAP7_75t_SL g476 ( .A(n_216), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_218), .Y(n_372) );
INVxp33_ASAP7_75t_L g1341 ( .A(n_219), .Y(n_1341) );
INVxp67_ASAP7_75t_SL g474 ( .A(n_220), .Y(n_474) );
INVx1_ASAP7_75t_L g820 ( .A(n_221), .Y(n_820) );
INVx2_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
XNOR2x1_ASAP7_75t_L g618 ( .A(n_223), .B(n_619), .Y(n_618) );
INVxp33_ASAP7_75t_SL g448 ( .A(n_224), .Y(n_448) );
INVxp67_ASAP7_75t_L g769 ( .A(n_225), .Y(n_769) );
INVx1_ASAP7_75t_L g888 ( .A(n_226), .Y(n_888) );
INVx1_ASAP7_75t_L g450 ( .A(n_227), .Y(n_450) );
BUFx3_ASAP7_75t_L g369 ( .A(n_228), .Y(n_369) );
INVx1_ASAP7_75t_L g394 ( .A(n_228), .Y(n_394) );
BUFx3_ASAP7_75t_L g371 ( .A(n_229), .Y(n_371) );
INVx1_ASAP7_75t_L g390 ( .A(n_229), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_230), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g868 ( .A(n_231), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_232), .Y(n_705) );
INVxp33_ASAP7_75t_L g264 ( .A(n_233), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_255), .B(n_1074), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_237), .B(n_242), .Y(n_236) );
AND2x4_ASAP7_75t_L g1348 ( .A(n_237), .B(n_243), .Y(n_1348) );
NOR2xp33_ASAP7_75t_SL g237 ( .A(n_238), .B(n_240), .Y(n_237) );
INVx1_ASAP7_75t_SL g1351 ( .A(n_238), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_238), .B(n_240), .Y(n_1361) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_240), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVxp67_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g558 ( .A(n_246), .B(n_254), .Y(n_558) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g310 ( .A(n_247), .B(n_311), .Y(n_310) );
OR2x6_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
INVx2_ASAP7_75t_SL g325 ( .A(n_249), .Y(n_325) );
INVx2_ASAP7_75t_SL g341 ( .A(n_249), .Y(n_341) );
OR2x2_ASAP7_75t_L g357 ( .A(n_249), .B(n_300), .Y(n_357) );
BUFx2_ASAP7_75t_L g674 ( .A(n_249), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_249), .A2(n_329), .B1(n_636), .B2(n_682), .Y(n_681) );
BUFx6f_ASAP7_75t_L g776 ( .A(n_249), .Y(n_776) );
INVx1_ASAP7_75t_L g904 ( .A(n_249), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_249), .A2(n_329), .B1(n_979), .B2(n_1005), .Y(n_1004) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
AND2x4_ASAP7_75t_L g268 ( .A(n_251), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g278 ( .A(n_251), .Y(n_278) );
AND2x2_ASAP7_75t_L g284 ( .A(n_251), .B(n_252), .Y(n_284) );
INVx2_ASAP7_75t_L g289 ( .A(n_251), .Y(n_289) );
INVx1_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
INVx2_ASAP7_75t_L g269 ( .A(n_252), .Y(n_269) );
INVx1_ASAP7_75t_L g291 ( .A(n_252), .Y(n_291) );
INVx1_ASAP7_75t_L g298 ( .A(n_252), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_252), .B(n_289), .Y(n_319) );
INVx1_ASAP7_75t_L g331 ( .A(n_252), .Y(n_331) );
INVx2_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
XNOR2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_857), .Y(n_255) );
XOR2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_613), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_437), .B1(n_438), .B2(n_612), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx2_ASAP7_75t_SL g612 ( .A(n_259), .Y(n_612) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_354), .Y(n_260) );
NOR3xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_292), .C(n_308), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_279), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B1(n_274), .B2(n_275), .Y(n_263) );
BUFx2_ASAP7_75t_L g445 ( .A(n_265), .Y(n_445) );
BUFx2_ASAP7_75t_L g549 ( .A(n_265), .Y(n_549) );
BUFx2_ASAP7_75t_L g661 ( .A(n_265), .Y(n_661) );
BUFx2_ASAP7_75t_L g790 ( .A(n_265), .Y(n_790) );
BUFx2_ASAP7_75t_L g825 ( .A(n_265), .Y(n_825) );
BUFx2_ASAP7_75t_L g894 ( .A(n_265), .Y(n_894) );
AND2x4_ASAP7_75t_L g265 ( .A(n_266), .B(n_270), .Y(n_265) );
BUFx3_ASAP7_75t_L g772 ( .A(n_266), .Y(n_772) );
INVx1_ASAP7_75t_L g782 ( .A(n_266), .Y(n_782) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g337 ( .A(n_267), .Y(n_337) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_267), .Y(n_462) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_268), .Y(n_322) );
AND2x4_ASAP7_75t_L g277 ( .A(n_269), .B(n_278), .Y(n_277) );
AND2x6_ASAP7_75t_L g275 ( .A(n_270), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g281 ( .A(n_270), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g286 ( .A(n_270), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g449 ( .A(n_270), .B(n_287), .Y(n_449) );
AND2x2_ASAP7_75t_L g554 ( .A(n_270), .B(n_287), .Y(n_554) );
AND2x2_ASAP7_75t_L g657 ( .A(n_270), .B(n_287), .Y(n_657) );
AND2x2_ASAP7_75t_L g664 ( .A(n_270), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g703 ( .A(n_270), .B(n_287), .Y(n_703) );
AND2x2_ASAP7_75t_L g707 ( .A(n_270), .B(n_337), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_270), .A2(n_573), .B1(n_944), .B2(n_951), .Y(n_943) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_270), .B(n_572), .Y(n_1006) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g350 ( .A(n_271), .Y(n_350) );
INVx1_ASAP7_75t_L g311 ( .A(n_273), .Y(n_311) );
INVx1_ASAP7_75t_L g352 ( .A(n_273), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_275), .A2(n_444), .B1(n_445), .B2(n_446), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_275), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_275), .A2(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_275), .A2(n_703), .B1(n_704), .B2(n_705), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_275), .A2(n_751), .B1(n_789), .B2(n_790), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_275), .A2(n_824), .B1(n_825), .B2(n_826), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_275), .A2(n_872), .B1(n_893), .B2(n_894), .Y(n_892) );
INVx1_ASAP7_75t_SL g1014 ( .A(n_275), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_275), .A2(n_825), .B1(n_1310), .B2(n_1311), .Y(n_1309) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_276), .B(n_299), .Y(n_307) );
BUFx2_ASAP7_75t_L g1319 ( .A(n_276), .Y(n_1319) );
BUFx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_277), .Y(n_470) );
BUFx3_ASAP7_75t_L g479 ( .A(n_277), .Y(n_479) );
BUFx2_ASAP7_75t_L g538 ( .A(n_277), .Y(n_538) );
INVx1_ASAP7_75t_L g562 ( .A(n_277), .Y(n_562) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_277), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B1(n_285), .B2(n_286), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_281), .A2(n_453), .B(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_281), .A2(n_552), .B1(n_553), .B2(n_554), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_281), .B(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_281), .A2(n_657), .B1(n_752), .B2(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_281), .A2(n_657), .B1(n_828), .B2(n_829), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_281), .A2(n_554), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g1312 ( .A1(n_281), .A2(n_554), .B1(n_1313), .B2(n_1314), .Y(n_1312) );
INVx2_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_SL g665 ( .A(n_283), .Y(n_665) );
INVx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_284), .Y(n_467) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_288), .Y(n_565) );
INVx1_ASAP7_75t_L g669 ( .A(n_288), .Y(n_669) );
INVx1_ASAP7_75t_L g679 ( .A(n_288), .Y(n_679) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_288), .Y(n_693) );
BUFx2_ASAP7_75t_L g1321 ( .A(n_288), .Y(n_1321) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g305 ( .A(n_289), .Y(n_305) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g899 ( .A(n_294), .Y(n_899) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2x1_ASAP7_75t_SL g295 ( .A(n_296), .B(n_299), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_298), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g303 ( .A(n_299), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g530 ( .A(n_299), .B(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g535 ( .A(n_299), .B(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g537 ( .A(n_299), .B(n_538), .Y(n_537) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx4f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx4f_ASAP7_75t_L g785 ( .A(n_303), .Y(n_785) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g786 ( .A(n_307), .Y(n_786) );
BUFx2_ASAP7_75t_L g900 ( .A(n_307), .Y(n_900) );
OAI33xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_313), .A3(n_323), .B1(n_334), .B2(n_339), .B3(n_347), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_309), .A2(n_347), .B1(n_455), .B2(n_471), .Y(n_454) );
OAI33xp33_ASAP7_75t_L g767 ( .A1(n_309), .A2(n_347), .A3(n_768), .B1(n_773), .B2(n_780), .B3(n_783), .Y(n_767) );
OAI33xp33_ASAP7_75t_L g797 ( .A1(n_309), .A2(n_347), .A3(n_798), .B1(n_804), .B2(n_809), .B3(n_816), .Y(n_797) );
OAI33xp33_ASAP7_75t_L g901 ( .A1(n_309), .A2(n_347), .A3(n_902), .B1(n_907), .B2(n_910), .B3(n_912), .Y(n_901) );
OR2x6_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
BUFx2_ASAP7_75t_L g436 ( .A(n_312), .Y(n_436) );
INVx2_ASAP7_75t_L g526 ( .A(n_312), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_320), .B2(n_321), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_315), .A2(n_335), .B1(n_336), .B2(n_338), .Y(n_334) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_315), .A2(n_769), .B1(n_770), .B2(n_771), .Y(n_768) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g781 ( .A(n_316), .Y(n_781) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g473 ( .A(n_318), .Y(n_473) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g458 ( .A(n_319), .Y(n_458) );
INVx1_ASAP7_75t_L g802 ( .A(n_319), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_321), .A2(n_817), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
INVx4_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_SL g475 ( .A(n_322), .Y(n_475) );
INVx2_ASAP7_75t_SL g567 ( .A(n_322), .Y(n_567) );
BUFx3_ASAP7_75t_L g569 ( .A(n_322), .Y(n_569) );
INVx2_ASAP7_75t_SL g946 ( .A(n_322), .Y(n_946) );
INVx2_ASAP7_75t_SL g960 ( .A(n_322), .Y(n_960) );
OAI22xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_326), .B1(n_327), .B2(n_333), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_327), .A2(n_805), .B1(n_806), .B2(n_808), .Y(n_804) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g1034 ( .A(n_328), .Y(n_1034) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_329), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
BUFx3_ASAP7_75t_L g1027 ( .A(n_329), .Y(n_1027) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g345 ( .A(n_331), .B(n_332), .Y(n_345) );
INVx1_ASAP7_75t_L g532 ( .A(n_332), .Y(n_532) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_335), .A2(n_375), .B1(n_385), .B2(n_395), .C(n_398), .Y(n_374) );
INVx2_ASAP7_75t_L g680 ( .A(n_336), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_336), .A2(n_799), .B1(n_800), .B2(n_803), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_336), .A2(n_456), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g671 ( .A(n_337), .Y(n_671) );
INVx1_ASAP7_75t_L g953 ( .A(n_337), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_338), .A2(n_342), .B1(n_426), .B2(n_431), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_343), .B2(n_346), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_340), .A2(n_343), .B1(n_757), .B2(n_764), .Y(n_783) );
INVx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_343), .A2(n_806), .B1(n_877), .B2(n_888), .Y(n_912) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g779 ( .A(n_344), .Y(n_779) );
OAI22xp33_ASAP7_75t_L g954 ( .A1(n_344), .A2(n_776), .B1(n_927), .B2(n_955), .Y(n_954) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_344), .A2(n_776), .B1(n_962), .B2(n_963), .Y(n_961) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g814 ( .A(n_345), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_346), .A2(n_409), .B1(n_417), .B2(n_420), .C(n_422), .Y(n_408) );
CKINVDCx8_ASAP7_75t_R g347 ( .A(n_348), .Y(n_347) );
INVx5_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx6_ASAP7_75t_L g573 ( .A(n_349), .Y(n_573) );
OR2x6_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx2_ASAP7_75t_L g698 ( .A(n_351), .Y(n_698) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AOI21xp33_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_372), .B(n_373), .Y(n_354) );
AOI21xp33_ASAP7_75t_L g736 ( .A1(n_355), .A2(n_737), .B(n_738), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g830 ( .A1(n_355), .A2(n_831), .B1(n_832), .B2(n_852), .Y(n_830) );
AOI21xp33_ASAP7_75t_SL g864 ( .A1(n_355), .A2(n_865), .B(n_866), .Y(n_864) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_355), .A2(n_831), .B1(n_1328), .B2(n_1343), .Y(n_1327) );
INVx5_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g575 ( .A(n_356), .Y(n_575) );
AND2x4_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx2_ASAP7_75t_L g451 ( .A(n_357), .Y(n_451) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx2_ASAP7_75t_L g645 ( .A(n_361), .Y(n_645) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_367), .Y(n_361) );
AND2x4_ASAP7_75t_L g400 ( .A(n_362), .B(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g405 ( .A(n_362), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
BUFx2_ASAP7_75t_L g510 ( .A(n_362), .Y(n_510) );
AND2x2_ASAP7_75t_L g513 ( .A(n_362), .B(n_406), .Y(n_513) );
AND2x2_ASAP7_75t_L g583 ( .A(n_362), .B(n_406), .Y(n_583) );
AND2x4_ASAP7_75t_L g647 ( .A(n_362), .B(n_401), .Y(n_647) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x4_ASAP7_75t_L g383 ( .A(n_365), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g416 ( .A(n_366), .B(n_384), .Y(n_416) );
INVx6_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
BUFx2_ASAP7_75t_L g508 ( .A(n_367), .Y(n_508) );
INVx2_ASAP7_75t_L g604 ( .A(n_367), .Y(n_604) );
AND2x4_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g407 ( .A(n_368), .Y(n_407) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g378 ( .A(n_369), .B(n_371), .Y(n_378) );
AND2x4_ASAP7_75t_L g389 ( .A(n_369), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g403 ( .A(n_370), .Y(n_403) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g393 ( .A(n_371), .B(n_394), .Y(n_393) );
AOI31xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_408), .A3(n_425), .B(n_434), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g729 ( .A1(n_376), .A2(n_396), .B(n_730), .C(n_731), .Y(n_729) );
BUFx4f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g421 ( .A(n_377), .B(n_396), .Y(n_421) );
INVx2_ASAP7_75t_SL g624 ( .A(n_377), .Y(n_624) );
AND2x4_ASAP7_75t_L g634 ( .A(n_377), .B(n_510), .Y(n_634) );
BUFx3_ASAP7_75t_L g759 ( .A(n_377), .Y(n_759) );
BUFx6f_ASAP7_75t_L g1046 ( .A(n_377), .Y(n_1046) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g762 ( .A(n_380), .Y(n_762) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
INVx1_ASAP7_75t_L g486 ( .A(n_381), .Y(n_486) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_381), .Y(n_633) );
INVx2_ASAP7_75t_SL g717 ( .A(n_381), .Y(n_717) );
INVx2_ASAP7_75t_L g875 ( .A(n_381), .Y(n_875) );
INVx1_ASAP7_75t_L g936 ( .A(n_381), .Y(n_936) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_383), .Y(n_505) );
INVx2_ASAP7_75t_L g589 ( .A(n_383), .Y(n_589) );
INVx2_ASAP7_75t_SL g726 ( .A(n_383), .Y(n_726) );
INVx1_ASAP7_75t_L g991 ( .A(n_383), .Y(n_991) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g395 ( .A(n_388), .B(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g585 ( .A(n_388), .Y(n_585) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g410 ( .A(n_389), .Y(n_410) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_389), .Y(n_493) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_389), .Y(n_499) );
INVx2_ASAP7_75t_SL g596 ( .A(n_389), .Y(n_596) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_389), .Y(n_630) );
BUFx2_ASAP7_75t_L g641 ( .A(n_389), .Y(n_641) );
BUFx3_ASAP7_75t_L g720 ( .A(n_389), .Y(n_720) );
BUFx6f_ASAP7_75t_L g835 ( .A(n_389), .Y(n_835) );
INVx1_ASAP7_75t_L g430 ( .A(n_390), .Y(n_430) );
INVx1_ASAP7_75t_L g1056 ( .A(n_391), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g433 ( .A(n_393), .Y(n_433) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_393), .Y(n_483) );
INVx1_ASAP7_75t_L g746 ( .A(n_393), .Y(n_746) );
INVx1_ASAP7_75t_L g1041 ( .A(n_393), .Y(n_1041) );
INVx1_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_395), .A2(n_579), .B(n_580), .C(n_584), .Y(n_578) );
AOI211xp5_ASAP7_75t_L g739 ( .A1(n_395), .A2(n_740), .B(n_741), .C(n_744), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_395), .A2(n_426), .B1(n_812), .B2(n_818), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_395), .A2(n_868), .B(n_869), .Y(n_867) );
AOI21xp33_ASAP7_75t_L g1329 ( .A1(n_395), .A2(n_1330), .B(n_1331), .Y(n_1329) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_396), .A2(n_516), .B(n_521), .Y(n_515) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_396), .A2(n_426), .B1(n_636), .B2(n_637), .C(n_644), .Y(n_635) );
AOI222xp33_ASAP7_75t_L g921 ( .A1(n_396), .A2(n_400), .B1(n_513), .B2(n_922), .C1(n_928), .C2(n_929), .Y(n_921) );
OAI21xp5_ASAP7_75t_L g968 ( .A1(n_396), .A2(n_969), .B(n_971), .Y(n_968) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g427 ( .A(n_397), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g432 ( .A(n_397), .B(n_433), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_SL g1037 ( .A1(n_397), .A2(n_1038), .B(n_1042), .C(n_1047), .Y(n_1037) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_400), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_511) );
INVx1_ASAP7_75t_L g581 ( .A(n_400), .Y(n_581) );
INVx1_ASAP7_75t_L g742 ( .A(n_400), .Y(n_742) );
AOI322xp5_ASAP7_75t_L g839 ( .A1(n_400), .A2(n_583), .A3(n_840), .B1(n_844), .B2(n_846), .C1(n_848), .C2(n_849), .Y(n_839) );
INVx2_ASAP7_75t_SL g1049 ( .A(n_400), .Y(n_1049) );
INVxp67_ASAP7_75t_L g976 ( .A(n_401), .Y(n_976) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g648 ( .A(n_405), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_405), .A2(n_647), .B1(n_687), .B2(n_688), .Y(n_732) );
INVx1_ASAP7_75t_L g977 ( .A(n_406), .Y(n_977) );
INVx2_ASAP7_75t_L g1051 ( .A(n_406), .Y(n_1051) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_411), .A2(n_450), .B(n_508), .C(n_509), .Y(n_507) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g422 ( .A(n_412), .B(n_423), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g925 ( .A1(n_412), .A2(n_835), .B1(n_926), .B2(n_927), .Y(n_925) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g600 ( .A(n_413), .Y(n_600) );
INVx1_ASAP7_75t_L g883 ( .A(n_413), .Y(n_883) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_415), .A2(n_1021), .B1(n_1026), .B2(n_1058), .C(n_1060), .Y(n_1057) );
BUFx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g495 ( .A(n_416), .Y(n_495) );
INVx2_ASAP7_75t_L g984 ( .A(n_416), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_418), .A2(n_1030), .B1(n_1032), .B2(n_1039), .Y(n_1038) );
INVx4_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g974 ( .A(n_419), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_420), .A2(n_422), .B1(n_877), .B2(n_878), .C(n_885), .Y(n_876) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g592 ( .A(n_421), .Y(n_592) );
INVx1_ASAP7_75t_L g756 ( .A(n_421), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_422), .A2(n_591), .B1(n_593), .B2(n_594), .C(n_601), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g754 ( .A1(n_422), .A2(n_755), .B1(n_757), .B2(n_758), .C(n_760), .Y(n_754) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_422), .A2(n_755), .B1(n_815), .B2(n_834), .C(n_836), .Y(n_833) );
AOI21xp33_ASAP7_75t_L g930 ( .A1(n_422), .A2(n_931), .B(n_932), .Y(n_930) );
INVx1_ASAP7_75t_L g1047 ( .A(n_422), .Y(n_1047) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_424), .B(n_1051), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_426), .A2(n_431), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_426), .A2(n_431), .B1(n_764), .B2(n_765), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_426), .A2(n_431), .B1(n_888), .B2(n_889), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_426), .A2(n_431), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
INVx6_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g504 ( .A(n_428), .Y(n_504) );
INVx2_ASAP7_75t_L g518 ( .A(n_428), .Y(n_518) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
AND2x2_ASAP7_75t_L g490 ( .A(n_429), .B(n_430), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_431), .B(n_820), .Y(n_851) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g520 ( .A(n_433), .Y(n_520) );
INVx2_ASAP7_75t_L g607 ( .A(n_433), .Y(n_607) );
AOI31xp33_ASAP7_75t_L g738 ( .A1(n_434), .A2(n_739), .A3(n_754), .B(n_763), .Y(n_738) );
BUFx8_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g831 ( .A(n_435), .Y(n_831) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g650 ( .A(n_436), .Y(n_650) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AO22x2_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_539), .B1(n_540), .B2(n_611), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g611 ( .A(n_440), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_442), .B(n_452), .C(n_480), .D(n_527), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_447), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g500 ( .A1(n_446), .A2(n_453), .B1(n_501), .B2(n_503), .C(n_505), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .B1(n_450), .B2(n_451), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_451), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_451), .A2(n_707), .B1(n_708), .B2(n_709), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g956 ( .A1(n_451), .A2(n_676), .B1(n_939), .B2(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_451), .A2(n_530), .B1(n_973), .B2(n_995), .Y(n_994) );
OAI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_459), .B1(n_460), .B2(n_463), .C(n_464), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_459), .A2(n_488), .B1(n_491), .B2(n_492), .C(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g694 ( .A(n_462), .Y(n_694) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g691 ( .A(n_466), .Y(n_691) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g560 ( .A(n_467), .Y(n_560) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_467), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g947 ( .A1(n_468), .A2(n_948), .B1(n_949), .B2(n_950), .Y(n_947) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B1(n_475), .B2(n_476), .C(n_477), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g817 ( .A(n_473), .Y(n_817) );
INVx2_ASAP7_75t_L g945 ( .A(n_473), .Y(n_945) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OAI31xp33_ASAP7_75t_SL g480 ( .A1(n_481), .A2(n_496), .A3(n_506), .B(n_524), .Y(n_480) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g628 ( .A(n_483), .Y(n_628) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_483), .Y(n_643) );
INVx1_ASAP7_75t_L g843 ( .A(n_483), .Y(n_843) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx4f_ASAP7_75t_L g502 ( .A(n_490), .Y(n_502) );
INVx1_ASAP7_75t_L g639 ( .A(n_490), .Y(n_639) );
INVx2_ASAP7_75t_L g723 ( .A(n_490), .Y(n_723) );
INVx1_ASAP7_75t_L g750 ( .A(n_490), .Y(n_750) );
INVx1_ASAP7_75t_L g1059 ( .A(n_490), .Y(n_1059) );
INVx2_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g748 ( .A(n_493), .Y(n_748) );
BUFx3_ASAP7_75t_L g1061 ( .A(n_493), .Y(n_1061) );
INVx1_ASAP7_75t_L g884 ( .A(n_494), .Y(n_884) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g522 ( .A(n_499), .Y(n_522) );
BUFx3_ASAP7_75t_L g626 ( .A(n_499), .Y(n_626) );
OAI211xp5_ASAP7_75t_L g871 ( .A1(n_501), .A2(n_872), .B(n_873), .C(n_874), .Y(n_871) );
OAI211xp5_ASAP7_75t_L g1332 ( .A1(n_501), .A2(n_1311), .B(n_1333), .C(n_1334), .Y(n_1332) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g523 ( .A(n_502), .Y(n_523) );
INVx1_ASAP7_75t_L g587 ( .A(n_502), .Y(n_587) );
INVx1_ASAP7_75t_L g715 ( .A(n_502), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_503), .A2(n_550), .B1(n_552), .B2(n_587), .C(n_588), .Y(n_586) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_503), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_749) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .C(n_515), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g972 ( .A1(n_509), .A2(n_973), .B(n_974), .C(n_975), .Y(n_972) );
BUFx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_512), .A2(n_514), .B1(n_528), .B2(n_533), .C(n_537), .Y(n_527) );
INVx3_ASAP7_75t_L g743 ( .A(n_513), .Y(n_743) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g923 ( .A(n_518), .Y(n_923) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_518), .Y(n_1055) );
INVx2_ASAP7_75t_L g1068 ( .A(n_518), .Y(n_1068) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g1338 ( .A(n_522), .Y(n_1338) );
OAI31xp33_ASAP7_75t_L g1036 ( .A1(n_524), .A2(n_1037), .A3(n_1048), .B(n_1052), .Y(n_1036) );
CKINVDCx8_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
AOI31xp33_ASAP7_75t_L g577 ( .A1(n_525), .A2(n_578), .A3(n_590), .B(n_608), .Y(n_577) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g557 ( .A(n_526), .B(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g676 ( .A(n_526), .B(n_558), .Y(n_676) );
AND2x2_ASAP7_75t_L g697 ( .A(n_526), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g941 ( .A(n_526), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_528), .A2(n_535), .B1(n_544), .B2(n_545), .C(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_530), .A2(n_535), .B1(n_537), .B2(n_653), .C(n_654), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_530), .A2(n_535), .B1(n_537), .B2(n_687), .C(n_688), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g964 ( .A1(n_530), .A2(n_535), .B1(n_537), .B2(n_928), .C(n_929), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g1306 ( .A1(n_530), .A2(n_535), .B1(n_537), .B2(n_1307), .C(n_1308), .Y(n_1306) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g1007 ( .A1(n_535), .A2(n_537), .B(n_1008), .Y(n_1007) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_537), .Y(n_546) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_574), .Y(n_541) );
AND4x1_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .C(n_551), .D(n_555), .Y(n_542) );
AOI33xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .A3(n_563), .B1(n_568), .B2(n_570), .B3(n_573), .Y(n_555) );
BUFx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g819 ( .A(n_569), .Y(n_819) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI222xp33_ASAP7_75t_L g663 ( .A1(n_573), .A2(n_664), .B1(n_666), .B2(n_667), .C1(n_676), .C2(n_677), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g1000 ( .A1(n_573), .A2(n_676), .A3(n_986), .B1(n_1001), .B2(n_1002), .C1(n_1003), .C2(n_1006), .Y(n_1000) );
AOI33xp33_ASAP7_75t_L g1315 ( .A1(n_573), .A2(n_1316), .A3(n_1317), .B1(n_1320), .B2(n_1322), .B3(n_1324), .Y(n_1315) );
AOI21xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B(n_577), .Y(n_574) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVxp67_ASAP7_75t_L g1064 ( .A(n_585), .Y(n_1064) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx2_ASAP7_75t_L g847 ( .A(n_589), .Y(n_847) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g841 ( .A(n_596), .Y(n_841) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx2_ASAP7_75t_L g718 ( .A(n_607), .Y(n_718) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_733), .B1(n_854), .B2(n_855), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g856 ( .A(n_616), .Y(n_856) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
XNOR2x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_683), .Y(n_617) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_620), .B(n_651), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_635), .B(n_649), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B1(n_629), .B2(n_631), .C(n_634), .Y(n_621) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g845 ( .A(n_624), .Y(n_845) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_628), .A2(n_1063), .B1(n_1064), .B2(n_1065), .Y(n_1062) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g727 ( .A(n_634), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_634), .A2(n_755), .B1(n_1336), .B2(n_1337), .C(n_1339), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g938 ( .A(n_645), .Y(n_938) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g870 ( .A(n_647), .Y(n_870) );
AOI31xp33_ASAP7_75t_L g866 ( .A1(n_649), .A2(n_867), .A3(n_876), .B(n_887), .Y(n_866) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI31xp33_ASAP7_75t_L g710 ( .A1(n_650), .A2(n_711), .A3(n_712), .B(n_728), .Y(n_710) );
NAND4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .C(n_659), .D(n_663), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_664), .A2(n_707), .B1(n_997), .B2(n_998), .Y(n_996) );
INVx1_ASAP7_75t_L g1035 ( .A(n_664), .Y(n_1035) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_671), .Y(n_911) );
AOI33xp33_ASAP7_75t_L g689 ( .A1(n_676), .A2(n_690), .A3(n_692), .B1(n_695), .B2(n_696), .B3(n_697), .Y(n_689) );
BUFx2_ASAP7_75t_L g1316 ( .A(n_676), .Y(n_1316) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g958 ( .A(n_679), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_701), .C(n_710), .Y(n_684) );
AND3x1_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .C(n_699), .Y(n_685) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g993 ( .A(n_703), .Y(n_993) );
INVx1_ASAP7_75t_L g1013 ( .A(n_703), .Y(n_1013) );
OAI211xp5_ASAP7_75t_L g721 ( .A1(n_705), .A2(n_722), .B(n_724), .C(n_725), .Y(n_721) );
INVx2_ASAP7_75t_L g1016 ( .A(n_707), .Y(n_1016) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_721), .C(n_727), .Y(n_712) );
OAI211xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B(n_716), .C(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g838 ( .A(n_717), .Y(n_838) );
INVx1_ASAP7_75t_L g924 ( .A(n_718), .Y(n_924) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_720), .Y(n_1044) );
OAI211xp5_ASAP7_75t_L g978 ( .A1(n_722), .A2(n_979), .B(n_980), .C(n_981), .Y(n_978) );
BUFx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g988 ( .A(n_723), .Y(n_988) );
INVx1_ASAP7_75t_L g753 ( .A(n_726), .Y(n_753) );
INVx1_ASAP7_75t_L g854 ( .A(n_733), .Y(n_854) );
XOR2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_793), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_766), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_740), .A2(n_765), .B1(n_781), .B2(n_782), .Y(n_780) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g937 ( .A(n_746), .Y(n_937) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NOR3xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_784), .C(n_787), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_773) );
BUFx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g807 ( .A(n_776), .Y(n_807) );
INVx1_ASAP7_75t_L g811 ( .A(n_776), .Y(n_811) );
OAI22xp5_ASAP7_75t_SL g1031 ( .A1(n_776), .A2(n_1032), .B1(n_1033), .B2(n_1034), .Y(n_1031) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_791), .Y(n_787) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_830), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_821), .C(n_822), .Y(n_796) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_801), .A2(n_819), .B1(n_908), .B2(n_909), .Y(n_907) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B1(n_813), .B2(n_815), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_813), .A2(n_903), .B1(n_905), .B2(n_906), .Y(n_902) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_817), .A2(n_868), .B1(n_889), .B2(n_911), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_827), .Y(n_822) );
NAND4xp25_ASAP7_75t_L g832 ( .A(n_833), .B(n_839), .C(n_850), .D(n_851), .Y(n_832) );
INVx1_ASAP7_75t_L g880 ( .A(n_835), .Y(n_880) );
INVx1_ASAP7_75t_L g970 ( .A(n_835), .Y(n_970) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
XNOR2x1_ASAP7_75t_L g860 ( .A(n_861), .B(n_914), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
XNOR2x1_ASAP7_75t_L g862 ( .A(n_863), .B(n_913), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_890), .Y(n_863) );
BUFx3_ASAP7_75t_L g886 ( .A(n_875), .Y(n_886) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
HB1xp67_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR3xp33_ASAP7_75t_SL g890 ( .A(n_891), .B(n_898), .C(n_901), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_892), .B(n_895), .Y(n_891) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g1025 ( .A(n_904), .Y(n_1025) );
OAI22x1_ASAP7_75t_L g914 ( .A1(n_915), .A2(n_916), .B1(n_1009), .B2(n_1073), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
XNOR2x1_ASAP7_75t_L g916 ( .A(n_917), .B(n_965), .Y(n_916) );
XNOR2x1_ASAP7_75t_L g917 ( .A(n_918), .B(n_919), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_918), .A2(n_1130), .B1(n_1131), .B2(n_1132), .Y(n_1129) );
OR2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_942), .Y(n_919) );
AOI31xp33_ASAP7_75t_SL g920 ( .A1(n_921), .A2(n_930), .A3(n_933), .B(n_940), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_935), .B1(n_938), .B2(n_939), .Y(n_933) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
AOI211xp5_ASAP7_75t_L g966 ( .A1(n_941), .A2(n_967), .B(n_992), .C(n_999), .Y(n_966) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_956), .C(n_964), .Y(n_942) );
HB1xp67_ASAP7_75t_L g1318 ( .A(n_949), .Y(n_1318) );
INVx1_ASAP7_75t_L g1326 ( .A(n_949), .Y(n_1326) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g1323 ( .A(n_953), .Y(n_1323) );
INVxp67_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND4xp25_ASAP7_75t_L g967 ( .A(n_968), .B(n_972), .C(n_978), .D(n_985), .Y(n_967) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OAI211xp5_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_987), .B(n_989), .C(n_990), .Y(n_985) );
INVx2_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1070 ( .A(n_991), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1007), .Y(n_999) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1009), .Y(n_1073) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1010), .Y(n_1071) );
NAND3xp33_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1017), .C(n_1036), .Y(n_1010) );
NOR2xp33_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1015), .Y(n_1011) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_1022), .A2(n_1024), .B1(n_1054), .B2(n_1056), .Y(n_1053) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1025), .B1(n_1026), .B2(n_1027), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_1029), .A2(n_1033), .B1(n_1043), .B2(n_1045), .Y(n_1042) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
BUFx2_ASAP7_75t_SL g1045 ( .A(n_1046), .Y(n_1045) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_1053), .A2(n_1057), .B1(n_1062), .B2(n_1066), .Y(n_1052) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
OAI221xp5_ASAP7_75t_L g1066 ( .A1(n_1058), .A2(n_1067), .B1(n_1068), .B2(n_1069), .C(n_1070), .Y(n_1066) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1074 ( .A1(n_1075), .A2(n_1300), .B1(n_1302), .B2(n_1344), .C(n_1349), .Y(n_1074) );
NOR2x1_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1237), .Y(n_1075) );
NAND3xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1174), .C(n_1198), .Y(n_1076) );
AOI211xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1108), .B(n_1136), .C(n_1166), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1078), .B(n_1157), .Y(n_1240) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_1079), .A2(n_1099), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1099), .Y(n_1079) );
INVx2_ASAP7_75t_SL g1162 ( .A(n_1080), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1080), .B(n_1122), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1080), .B(n_1099), .Y(n_1246) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_1081), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1141 ( .A(n_1081), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1081), .B(n_1099), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1081), .B(n_1099), .Y(n_1219) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1082), .Y(n_1152) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1082), .Y(n_1184) );
AND2x4_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1086), .Y(n_1082) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1083), .B(n_1086), .Y(n_1107) );
HB1xp67_ASAP7_75t_L g1358 ( .A(n_1083), .Y(n_1358) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
AND2x4_ASAP7_75t_L g1088 ( .A(n_1084), .B(n_1086), .Y(n_1088) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_1085), .B(n_1095), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1087), .Y(n_1095) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1088), .Y(n_1126) );
INVx1_ASAP7_75t_SL g1132 ( .A(n_1088), .Y(n_1132) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1091), .B1(n_1096), .B2(n_1097), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_1091), .A2(n_1097), .B1(n_1134), .B2(n_1135), .Y(n_1133) );
OAI22xp33_ASAP7_75t_L g1145 ( .A1(n_1091), .A2(n_1146), .B1(n_1147), .B2(n_1148), .Y(n_1145) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_1091), .Y(n_1188) );
BUFx6f_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_1092), .A2(n_1097), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .Y(n_1092) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1093), .B(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1093), .Y(n_1103) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1094), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g1360 ( .A(n_1095), .Y(n_1360) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1097), .Y(n_1149) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1098), .Y(n_1105) );
INVx2_ASAP7_75t_L g1154 ( .A(n_1099), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1099), .B(n_1143), .Y(n_1169) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1099), .B(n_1143), .Y(n_1195) );
OAI21xp33_ASAP7_75t_L g1199 ( .A1(n_1099), .A2(n_1200), .B(n_1202), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1099), .B(n_1144), .Y(n_1230) );
AND2x4_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1106), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1103), .Y(n_1101) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_1103), .B(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1107), .Y(n_1130) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1120), .Y(n_1109) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1110), .B(n_1221), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1231 ( .A(n_1110), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1111), .B(n_1127), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1111), .B(n_1128), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1115), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1112), .B(n_1116), .Y(n_1139) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1112), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1112), .B(n_1128), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1259 ( .A(n_1112), .B(n_1116), .Y(n_1259) );
NOR2xp33_ASAP7_75t_SL g1289 ( .A(n_1112), .B(n_1290), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1114), .Y(n_1112) );
OR2x2_ASAP7_75t_L g1159 ( .A(n_1115), .B(n_1127), .Y(n_1159) );
NOR3xp33_ASAP7_75t_L g1179 ( .A(n_1115), .B(n_1157), .C(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1115), .B(n_1127), .Y(n_1210) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1116), .B(n_1127), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1116), .B(n_1172), .Y(n_1171) );
OAI322xp33_ASAP7_75t_L g1243 ( .A1(n_1116), .A2(n_1244), .A3(n_1247), .B1(n_1248), .B2(n_1250), .C1(n_1252), .C2(n_1254), .Y(n_1243) );
NOR2xp33_ASAP7_75t_L g1253 ( .A(n_1116), .B(n_1127), .Y(n_1253) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1127), .Y(n_1121) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1122), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1122), .B(n_1127), .Y(n_1173) );
INVx4_ASAP7_75t_L g1178 ( .A(n_1122), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1122), .B(n_1209), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1122), .B(n_1246), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1122), .B(n_1249), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1122), .B(n_1144), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1122), .B(n_1162), .Y(n_1290) );
AND2x6_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1124), .Y(n_1122) );
INVx2_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1182 ( .A1(n_1126), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1182) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1126), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1127), .B(n_1139), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1127), .B(n_1177), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1127), .B(n_1171), .Y(n_1233) );
CKINVDCx6p67_ASAP7_75t_R g1127 ( .A(n_1128), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_1128), .B(n_1177), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1128), .B(n_1171), .Y(n_1213) );
AOI32xp33_ASAP7_75t_L g1215 ( .A1(n_1128), .A2(n_1194), .A3(n_1216), .B1(n_1220), .B2(n_1222), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1128), .B(n_1139), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1128), .B(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1128), .B(n_1288), .Y(n_1287) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1128), .B(n_1294), .Y(n_1293) );
OR2x6_ASAP7_75t_SL g1128 ( .A(n_1129), .B(n_1133), .Y(n_1128) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_1132), .A2(n_1151), .B1(n_1152), .B2(n_1153), .Y(n_1150) );
OAI221xp5_ASAP7_75t_L g1136 ( .A1(n_1137), .A2(n_1140), .B1(n_1155), .B2(n_1160), .C(n_1163), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1139), .B(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1139), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1141), .Y(n_1272) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1141), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1142), .B(n_1164), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1154), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1143), .B(n_1162), .Y(n_1161) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1143), .Y(n_1207) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1143), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1143), .B(n_1191), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1143), .B(n_1181), .Y(n_1247) );
INVx3_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1144), .B(n_1219), .Y(n_1257) );
OR2x2_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1150), .Y(n_1144) );
HB1xp67_ASAP7_75t_L g1190 ( .A(n_1148), .Y(n_1190) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NOR2x1_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1159), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1157), .B(n_1213), .Y(n_1212) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1157), .B(n_1265), .Y(n_1264) );
NOR2x1_ASAP7_75t_R g1280 ( .A(n_1157), .B(n_1221), .Y(n_1280) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1158), .B(n_1165), .Y(n_1164) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1158), .B(n_1209), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1158), .B(n_1225), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1158), .B(n_1213), .Y(n_1298) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1159), .Y(n_1227) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
AOI322xp5_ASAP7_75t_L g1226 ( .A1(n_1161), .A2(n_1207), .A3(n_1227), .B1(n_1228), .B2(n_1230), .C1(n_1231), .C2(n_1233), .Y(n_1226) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1162), .Y(n_1168) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1162), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1162), .B(n_1230), .Y(n_1251) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1162), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1170), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1169), .Y(n_1167) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1169), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1173), .Y(n_1170) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1171), .Y(n_1221) );
AOI211xp5_ASAP7_75t_L g1275 ( .A1(n_1172), .A2(n_1276), .B(n_1277), .C(n_1280), .Y(n_1275) );
O2A1O1Ixp33_ASAP7_75t_L g1174 ( .A1(n_1175), .A2(n_1179), .B(n_1191), .C(n_1192), .Y(n_1174) );
INVxp67_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1178), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1178), .Y(n_1204) );
NOR2xp33_ASAP7_75t_L g1294 ( .A(n_1178), .B(n_1259), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1178), .B(n_1218), .Y(n_1296) );
OAI31xp33_ASAP7_75t_L g1198 ( .A1(n_1180), .A2(n_1199), .A3(n_1211), .B(n_1214), .Y(n_1198) );
OAI221xp5_ASAP7_75t_L g1285 ( .A1(n_1180), .A2(n_1219), .B1(n_1286), .B2(n_1291), .C(n_1295), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_1181), .Y(n_1180) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_1181), .A2(n_1261), .B1(n_1270), .B2(n_1271), .Y(n_1260) );
OR2x6_ASAP7_75t_SL g1181 ( .A(n_1182), .B(n_1186), .Y(n_1181) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_1187), .A2(n_1188), .B1(n_1189), .B2(n_1190), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1191), .B(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1196), .Y(n_1193) );
AOI322xp5_ASAP7_75t_L g1286 ( .A1(n_1194), .A2(n_1207), .A3(n_1210), .B1(n_1245), .B2(n_1246), .C1(n_1287), .C2(n_1289), .Y(n_1286) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1196), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1197), .Y(n_1223) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
OAI21xp5_ASAP7_75t_SL g1202 ( .A1(n_1203), .A2(n_1205), .B(n_1210), .Y(n_1202) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1204), .B(n_1225), .Y(n_1224) );
NOR2xp33_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_SL g1206 ( .A(n_1207), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1207), .B(n_1212), .Y(n_1211) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1207), .B(n_1233), .Y(n_1269) );
AOI21xp5_ASAP7_75t_L g1268 ( .A1(n_1208), .A2(n_1221), .B(n_1262), .Y(n_1268) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1208), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1210), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1213), .Y(n_1242) );
NAND3xp33_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1226), .C(n_1234), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1218), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1218), .B(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1241 ( .A(n_1223), .B(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1225), .Y(n_1262) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
A2O1A1Ixp33_ASAP7_75t_L g1282 ( .A1(n_1229), .A2(n_1242), .B(n_1258), .C(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1230), .Y(n_1265) );
AOI211xp5_ASAP7_75t_SL g1281 ( .A1(n_1230), .A2(n_1282), .B(n_1285), .C(n_1297), .Y(n_1281) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1232), .Y(n_1284) );
NOR2xp33_ASAP7_75t_L g1252 ( .A(n_1233), .B(n_1253), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1233), .B(n_1267), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1233), .B(n_1284), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1236), .Y(n_1234) );
AOI211xp5_ASAP7_75t_L g1263 ( .A1(n_1235), .A2(n_1264), .B(n_1266), .C(n_1268), .Y(n_1263) );
NAND3xp33_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1260), .C(n_1281), .Y(n_1237) );
AOI211xp5_ASAP7_75t_SL g1238 ( .A1(n_1239), .A2(n_1241), .B(n_1243), .C(n_1256), .Y(n_1238) );
INVxp67_ASAP7_75t_SL g1239 ( .A(n_1240), .Y(n_1239) );
OAI211xp5_ASAP7_75t_L g1271 ( .A1(n_1242), .A2(n_1272), .B(n_1273), .C(n_1275), .Y(n_1271) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1247), .Y(n_1270) );
OAI211xp5_ASAP7_75t_L g1261 ( .A1(n_1250), .A2(n_1262), .B(n_1263), .C(n_1269), .Y(n_1261) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
NOR2xp33_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1258), .Y(n_1256) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1259), .Y(n_1288) );
AOI21xp5_ASAP7_75t_L g1297 ( .A1(n_1291), .A2(n_1298), .B(n_1299), .Y(n_1297) );
INVxp67_ASAP7_75t_SL g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1304), .Y(n_1355) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1327), .Y(n_1304) );
AND4x1_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1309), .C(n_1312), .D(n_1315), .Y(n_1305) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1335), .C(n_1340), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g1344 ( .A(n_1345), .Y(n_1344) );
BUFx2_ASAP7_75t_L g1345 ( .A(n_1346), .Y(n_1345) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1347), .Y(n_1346) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
A2O1A1Ixp33_ASAP7_75t_L g1356 ( .A1(n_1351), .A2(n_1357), .B(n_1359), .C(n_1361), .Y(n_1356) );
INVxp33_ASAP7_75t_SL g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
endmodule